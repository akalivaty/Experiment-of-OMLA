

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U557 ( .A1(n529), .A2(n528), .ZN(n535) );
  XOR2_X1 U558 ( .A(KEYINPUT97), .B(n748), .Z(n524) );
  INV_X1 U559 ( .A(KEYINPUT94), .ZN(n684) );
  XNOR2_X1 U560 ( .A(n685), .B(n684), .ZN(n738) );
  NOR2_X1 U561 ( .A1(G651), .A2(n564), .ZN(n639) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n641) );
  NOR2_X1 U563 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n525), .Z(n881) );
  NAND2_X1 U565 ( .A1(G137), .A2(n881), .ZN(n526) );
  XNOR2_X1 U566 ( .A(KEYINPUT65), .B(n526), .ZN(n529) );
  INV_X1 U567 ( .A(G2105), .ZN(n530) );
  NOR2_X2 U568 ( .A1(G2104), .A2(n530), .ZN(n876) );
  NAND2_X1 U569 ( .A1(G125), .A2(n876), .ZN(n527) );
  XOR2_X1 U570 ( .A(KEYINPUT64), .B(n527), .Z(n528) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n877) );
  NAND2_X1 U572 ( .A1(n877), .A2(G113), .ZN(n533) );
  AND2_X1 U573 ( .A1(n530), .A2(G2104), .ZN(n880) );
  NAND2_X1 U574 ( .A1(G101), .A2(n880), .ZN(n531) );
  XOR2_X1 U575 ( .A(KEYINPUT23), .B(n531), .Z(n532) );
  NAND2_X1 U576 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U577 ( .A1(n535), .A2(n534), .ZN(G160) );
  NAND2_X1 U578 ( .A1(G91), .A2(n641), .ZN(n536) );
  XNOR2_X1 U579 ( .A(n536), .B(KEYINPUT68), .ZN(n545) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n564) );
  INV_X1 U581 ( .A(G651), .ZN(n537) );
  NOR2_X1 U582 ( .A1(n564), .A2(n537), .ZN(n640) );
  NAND2_X1 U583 ( .A1(G78), .A2(n640), .ZN(n540) );
  NOR2_X1 U584 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U585 ( .A(KEYINPUT1), .B(n538), .Z(n644) );
  NAND2_X1 U586 ( .A1(G65), .A2(n644), .ZN(n539) );
  NAND2_X1 U587 ( .A1(n540), .A2(n539), .ZN(n543) );
  NAND2_X1 U588 ( .A1(G53), .A2(n639), .ZN(n541) );
  XNOR2_X1 U589 ( .A(KEYINPUT69), .B(n541), .ZN(n542) );
  NOR2_X1 U590 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U591 ( .A1(n545), .A2(n544), .ZN(G299) );
  NAND2_X1 U592 ( .A1(G60), .A2(n644), .ZN(n547) );
  NAND2_X1 U593 ( .A1(G85), .A2(n641), .ZN(n546) );
  NAND2_X1 U594 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U595 ( .A1(G72), .A2(n640), .ZN(n549) );
  NAND2_X1 U596 ( .A1(G47), .A2(n639), .ZN(n548) );
  NAND2_X1 U597 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U598 ( .A1(n551), .A2(n550), .ZN(G290) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U600 ( .A(G57), .ZN(G237) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  NAND2_X1 U603 ( .A1(G64), .A2(n644), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G52), .A2(n639), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n559) );
  NAND2_X1 U606 ( .A1(n641), .A2(G90), .ZN(n554) );
  XNOR2_X1 U607 ( .A(n554), .B(KEYINPUT66), .ZN(n556) );
  NAND2_X1 U608 ( .A1(G77), .A2(n640), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n557), .Z(n558) );
  NOR2_X1 U611 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U612 ( .A(KEYINPUT67), .B(n560), .Z(G171) );
  NAND2_X1 U613 ( .A1(G49), .A2(n639), .ZN(n562) );
  NAND2_X1 U614 ( .A1(G74), .A2(G651), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U616 ( .A1(n644), .A2(n563), .ZN(n566) );
  NAND2_X1 U617 ( .A1(n564), .A2(G87), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(G288) );
  NAND2_X1 U619 ( .A1(G63), .A2(n644), .ZN(n568) );
  NAND2_X1 U620 ( .A1(G51), .A2(n639), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(n569), .ZN(n576) );
  NAND2_X1 U623 ( .A1(G89), .A2(n641), .ZN(n570) );
  XOR2_X1 U624 ( .A(KEYINPUT75), .B(n570), .Z(n571) );
  XNOR2_X1 U625 ( .A(n571), .B(KEYINPUT4), .ZN(n573) );
  NAND2_X1 U626 ( .A1(G76), .A2(n640), .ZN(n572) );
  NAND2_X1 U627 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U628 ( .A(n574), .B(KEYINPUT5), .Z(n575) );
  NOR2_X1 U629 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U630 ( .A(KEYINPUT76), .B(n577), .Z(n578) );
  XNOR2_X1 U631 ( .A(KEYINPUT7), .B(n578), .ZN(G168) );
  XOR2_X1 U632 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U634 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U635 ( .A(KEYINPUT71), .B(KEYINPUT11), .Z(n581) );
  INV_X1 U636 ( .A(G223), .ZN(n826) );
  NAND2_X1 U637 ( .A1(G567), .A2(n826), .ZN(n580) );
  XNOR2_X1 U638 ( .A(n581), .B(n580), .ZN(n582) );
  XOR2_X1 U639 ( .A(KEYINPUT70), .B(n582), .Z(G234) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n584) );
  NAND2_X1 U641 ( .A1(G56), .A2(n644), .ZN(n583) );
  XNOR2_X1 U642 ( .A(n584), .B(n583), .ZN(n591) );
  XNOR2_X1 U643 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n589) );
  NAND2_X1 U644 ( .A1(n641), .A2(G81), .ZN(n585) );
  XNOR2_X1 U645 ( .A(n585), .B(KEYINPUT12), .ZN(n587) );
  NAND2_X1 U646 ( .A1(G68), .A2(n640), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U648 ( .A(n589), .B(n588), .ZN(n590) );
  NOR2_X1 U649 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U650 ( .A1(n639), .A2(G43), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n593), .A2(n592), .ZN(n922) );
  INV_X1 U652 ( .A(G860), .ZN(n607) );
  OR2_X1 U653 ( .A1(n922), .A2(n607), .ZN(G153) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(G79), .A2(n640), .ZN(n595) );
  NAND2_X1 U656 ( .A1(G54), .A2(n639), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U658 ( .A1(G66), .A2(n644), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G92), .A2(n641), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U661 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U662 ( .A(n600), .B(KEYINPUT15), .ZN(n925) );
  INV_X1 U663 ( .A(G868), .ZN(n660) );
  NAND2_X1 U664 ( .A1(n925), .A2(n660), .ZN(n601) );
  XNOR2_X1 U665 ( .A(n601), .B(KEYINPUT74), .ZN(n603) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n602) );
  NAND2_X1 U667 ( .A1(n603), .A2(n602), .ZN(G284) );
  NOR2_X1 U668 ( .A1(G286), .A2(n660), .ZN(n604) );
  XOR2_X1 U669 ( .A(KEYINPUT77), .B(n604), .Z(n606) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U671 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n607), .A2(G559), .ZN(n608) );
  INV_X1 U673 ( .A(n925), .ZN(n656) );
  NAND2_X1 U674 ( .A1(n608), .A2(n656), .ZN(n609) );
  XNOR2_X1 U675 ( .A(n609), .B(KEYINPUT16), .ZN(n610) );
  XNOR2_X1 U676 ( .A(KEYINPUT78), .B(n610), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n922), .ZN(n613) );
  NAND2_X1 U678 ( .A1(G868), .A2(n656), .ZN(n611) );
  NOR2_X1 U679 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U680 ( .A1(n613), .A2(n612), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G123), .A2(n876), .ZN(n614) );
  XOR2_X1 U682 ( .A(KEYINPUT18), .B(n614), .Z(n615) );
  XNOR2_X1 U683 ( .A(n615), .B(KEYINPUT79), .ZN(n617) );
  NAND2_X1 U684 ( .A1(G111), .A2(n877), .ZN(n616) );
  NAND2_X1 U685 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U686 ( .A1(G99), .A2(n880), .ZN(n619) );
  NAND2_X1 U687 ( .A1(G135), .A2(n881), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U689 ( .A1(n621), .A2(n620), .ZN(n974) );
  XNOR2_X1 U690 ( .A(n974), .B(G2096), .ZN(n623) );
  INV_X1 U691 ( .A(G2100), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G62), .A2(n644), .ZN(n625) );
  NAND2_X1 U694 ( .A1(G50), .A2(n639), .ZN(n624) );
  NAND2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U696 ( .A(KEYINPUT84), .B(n626), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G75), .A2(n640), .ZN(n628) );
  NAND2_X1 U698 ( .A1(G88), .A2(n641), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U700 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U701 ( .A1(G61), .A2(n644), .ZN(n632) );
  NAND2_X1 U702 ( .A1(G48), .A2(n639), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n636) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n634) );
  NAND2_X1 U705 ( .A1(n640), .A2(G73), .ZN(n633) );
  XOR2_X1 U706 ( .A(n634), .B(n633), .Z(n635) );
  NOR2_X1 U707 ( .A1(n636), .A2(n635), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n641), .A2(G86), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G55), .A2(n639), .ZN(n649) );
  NAND2_X1 U711 ( .A1(G80), .A2(n640), .ZN(n643) );
  NAND2_X1 U712 ( .A1(G93), .A2(n641), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U714 ( .A1(G67), .A2(n644), .ZN(n645) );
  XNOR2_X1 U715 ( .A(KEYINPUT81), .B(n645), .ZN(n646) );
  NOR2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT82), .ZN(n918) );
  XNOR2_X1 U719 ( .A(n918), .B(KEYINPUT19), .ZN(n652) );
  INV_X1 U720 ( .A(G299), .ZN(n930) );
  XNOR2_X1 U721 ( .A(G288), .B(n930), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n652), .B(n651), .ZN(n653) );
  XOR2_X1 U723 ( .A(n653), .B(G305), .Z(n654) );
  XNOR2_X1 U724 ( .A(G290), .B(n654), .ZN(n655) );
  XNOR2_X1 U725 ( .A(G166), .B(n655), .ZN(n894) );
  NAND2_X1 U726 ( .A1(G559), .A2(n656), .ZN(n657) );
  XNOR2_X1 U727 ( .A(n657), .B(n922), .ZN(n915) );
  XNOR2_X1 U728 ( .A(n894), .B(n915), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n658), .A2(G868), .ZN(n659) );
  XOR2_X1 U730 ( .A(KEYINPUT85), .B(n659), .Z(n662) );
  NAND2_X1 U731 ( .A1(n918), .A2(n660), .ZN(n661) );
  NAND2_X1 U732 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U735 ( .A1(n664), .A2(G2090), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n665), .B(KEYINPUT21), .ZN(n666) );
  XNOR2_X1 U737 ( .A(KEYINPUT86), .B(n666), .ZN(n667) );
  NAND2_X1 U738 ( .A1(G2072), .A2(n667), .ZN(G158) );
  XNOR2_X1 U739 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U740 ( .A1(G220), .A2(G219), .ZN(n668) );
  XOR2_X1 U741 ( .A(KEYINPUT22), .B(n668), .Z(n669) );
  NOR2_X1 U742 ( .A1(G218), .A2(n669), .ZN(n670) );
  NAND2_X1 U743 ( .A1(G96), .A2(n670), .ZN(n919) );
  NAND2_X1 U744 ( .A1(n919), .A2(G2106), .ZN(n674) );
  NAND2_X1 U745 ( .A1(G69), .A2(G120), .ZN(n671) );
  NOR2_X1 U746 ( .A1(G237), .A2(n671), .ZN(n672) );
  NAND2_X1 U747 ( .A1(G108), .A2(n672), .ZN(n920) );
  NAND2_X1 U748 ( .A1(n920), .A2(G567), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n674), .A2(n673), .ZN(n830) );
  NAND2_X1 U750 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U751 ( .A1(n830), .A2(n675), .ZN(n676) );
  XOR2_X1 U752 ( .A(KEYINPUT87), .B(n676), .Z(n829) );
  NAND2_X1 U753 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U754 ( .A1(G102), .A2(n880), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G138), .A2(n881), .ZN(n677) );
  NAND2_X1 U756 ( .A1(n678), .A2(n677), .ZN(n682) );
  NAND2_X1 U757 ( .A1(G126), .A2(n876), .ZN(n680) );
  NAND2_X1 U758 ( .A1(G114), .A2(n877), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U760 ( .A1(n682), .A2(n681), .ZN(G164) );
  INV_X1 U761 ( .A(G166), .ZN(G303) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n772) );
  INV_X1 U763 ( .A(n772), .ZN(n683) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n771) );
  NAND2_X2 U765 ( .A1(n683), .A2(n771), .ZN(n720) );
  NOR2_X1 U766 ( .A1(G2084), .A2(n720), .ZN(n736) );
  NAND2_X2 U767 ( .A1(G8), .A2(n720), .ZN(n800) );
  NOR2_X1 U768 ( .A1(G1966), .A2(n800), .ZN(n685) );
  NAND2_X1 U769 ( .A1(n738), .A2(G8), .ZN(n686) );
  NOR2_X1 U770 ( .A1(n736), .A2(n686), .ZN(n687) );
  XOR2_X1 U771 ( .A(KEYINPUT30), .B(n687), .Z(n688) );
  NOR2_X1 U772 ( .A1(G168), .A2(n688), .ZN(n693) );
  XOR2_X1 U773 ( .A(KEYINPUT25), .B(G2078), .Z(n1011) );
  NOR2_X1 U774 ( .A1(n1011), .A2(n720), .ZN(n689) );
  XNOR2_X1 U775 ( .A(n689), .B(KEYINPUT95), .ZN(n691) );
  INV_X1 U776 ( .A(G1961), .ZN(n957) );
  NAND2_X1 U777 ( .A1(n957), .A2(n720), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n691), .A2(n690), .ZN(n695) );
  NOR2_X1 U779 ( .A1(G171), .A2(n695), .ZN(n692) );
  NOR2_X2 U780 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U781 ( .A(KEYINPUT31), .B(n694), .Z(n734) );
  NAND2_X1 U782 ( .A1(n695), .A2(G171), .ZN(n719) );
  INV_X1 U783 ( .A(n720), .ZN(n705) );
  NAND2_X1 U784 ( .A1(n705), .A2(G2072), .ZN(n696) );
  XNOR2_X1 U785 ( .A(n696), .B(KEYINPUT27), .ZN(n698) );
  INV_X1 U786 ( .A(G1956), .ZN(n948) );
  NOR2_X1 U787 ( .A1(n948), .A2(n705), .ZN(n697) );
  NOR2_X1 U788 ( .A1(n698), .A2(n697), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n930), .A2(n700), .ZN(n699) );
  XOR2_X1 U790 ( .A(n699), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U791 ( .A1(n930), .A2(n700), .ZN(n714) );
  INV_X1 U792 ( .A(G1996), .ZN(n1003) );
  NOR2_X1 U793 ( .A1(n720), .A2(n1003), .ZN(n701) );
  XOR2_X1 U794 ( .A(n701), .B(KEYINPUT26), .Z(n703) );
  NAND2_X1 U795 ( .A1(n720), .A2(G1341), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U797 ( .A1(n922), .A2(n704), .ZN(n709) );
  NAND2_X1 U798 ( .A1(G1348), .A2(n720), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n705), .A2(G2067), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n710) );
  NOR2_X1 U801 ( .A1(n925), .A2(n710), .ZN(n708) );
  OR2_X1 U802 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U803 ( .A1(n925), .A2(n710), .ZN(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U807 ( .A(KEYINPUT29), .B(n717), .Z(n718) );
  NAND2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n735) );
  INV_X1 U809 ( .A(G8), .ZN(n725) );
  NOR2_X1 U810 ( .A1(G1971), .A2(n800), .ZN(n722) );
  NOR2_X1 U811 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U813 ( .A1(n723), .A2(G303), .ZN(n724) );
  OR2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n727) );
  AND2_X1 U815 ( .A1(n735), .A2(n727), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n734), .A2(n726), .ZN(n731) );
  INV_X1 U817 ( .A(n727), .ZN(n729) );
  AND2_X1 U818 ( .A1(G286), .A2(G8), .ZN(n728) );
  OR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U821 ( .A(n732), .B(KEYINPUT32), .ZN(n796) );
  AND2_X1 U822 ( .A1(G1976), .A2(G288), .ZN(n927) );
  OR2_X1 U823 ( .A1(n800), .A2(n927), .ZN(n744) );
  INV_X1 U824 ( .A(n744), .ZN(n733) );
  AND2_X1 U825 ( .A1(n796), .A2(n733), .ZN(n742) );
  NAND2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n740) );
  NAND2_X1 U827 ( .A1(G8), .A2(n736), .ZN(n737) );
  AND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U830 ( .A(n741), .B(KEYINPUT96), .ZN(n797) );
  NAND2_X1 U831 ( .A1(n742), .A2(n797), .ZN(n746) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n743) );
  NOR2_X1 U834 ( .A1(n749), .A2(n743), .ZN(n942) );
  OR2_X1 U835 ( .A1(n744), .A2(n942), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U837 ( .A1(KEYINPUT33), .A2(n747), .ZN(n748) );
  NAND2_X1 U838 ( .A1(KEYINPUT33), .A2(n749), .ZN(n750) );
  NOR2_X1 U839 ( .A1(n800), .A2(n750), .ZN(n751) );
  NOR2_X1 U840 ( .A1(n524), .A2(n751), .ZN(n790) );
  XOR2_X1 U841 ( .A(KEYINPUT98), .B(G1981), .Z(n752) );
  XNOR2_X1 U842 ( .A(G305), .B(n752), .ZN(n937) );
  NAND2_X1 U843 ( .A1(G95), .A2(n880), .ZN(n753) );
  XNOR2_X1 U844 ( .A(n753), .B(KEYINPUT92), .ZN(n756) );
  NAND2_X1 U845 ( .A1(G119), .A2(n876), .ZN(n754) );
  XOR2_X1 U846 ( .A(KEYINPUT91), .B(n754), .Z(n755) );
  NAND2_X1 U847 ( .A1(n756), .A2(n755), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G131), .A2(n881), .ZN(n758) );
  NAND2_X1 U849 ( .A1(G107), .A2(n877), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U851 ( .A1(n760), .A2(n759), .ZN(n865) );
  INV_X1 U852 ( .A(G1991), .ZN(n1008) );
  NOR2_X1 U853 ( .A1(n865), .A2(n1008), .ZN(n770) );
  NAND2_X1 U854 ( .A1(G129), .A2(n876), .ZN(n762) );
  NAND2_X1 U855 ( .A1(G141), .A2(n881), .ZN(n761) );
  NAND2_X1 U856 ( .A1(n762), .A2(n761), .ZN(n766) );
  NAND2_X1 U857 ( .A1(G105), .A2(n880), .ZN(n763) );
  XNOR2_X1 U858 ( .A(n763), .B(KEYINPUT38), .ZN(n764) );
  XNOR2_X1 U859 ( .A(n764), .B(KEYINPUT93), .ZN(n765) );
  NOR2_X1 U860 ( .A1(n766), .A2(n765), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n877), .A2(G117), .ZN(n767) );
  NAND2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n866) );
  AND2_X1 U863 ( .A1(n866), .A2(G1996), .ZN(n769) );
  NOR2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n981) );
  NOR2_X1 U865 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U866 ( .A(n773), .B(KEYINPUT88), .Z(n785) );
  NOR2_X1 U867 ( .A1(n981), .A2(n785), .ZN(n812) );
  INV_X1 U868 ( .A(n812), .ZN(n786) );
  XNOR2_X1 U869 ( .A(G2067), .B(KEYINPUT37), .ZN(n817) );
  NAND2_X1 U870 ( .A1(n881), .A2(G140), .ZN(n774) );
  XOR2_X1 U871 ( .A(KEYINPUT89), .B(n774), .Z(n776) );
  NAND2_X1 U872 ( .A1(n880), .A2(G104), .ZN(n775) );
  NAND2_X1 U873 ( .A1(n776), .A2(n775), .ZN(n778) );
  XNOR2_X1 U874 ( .A(KEYINPUT90), .B(KEYINPUT34), .ZN(n777) );
  XNOR2_X1 U875 ( .A(n778), .B(n777), .ZN(n783) );
  NAND2_X1 U876 ( .A1(G128), .A2(n876), .ZN(n780) );
  NAND2_X1 U877 ( .A1(G116), .A2(n877), .ZN(n779) );
  NAND2_X1 U878 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U879 ( .A(KEYINPUT35), .B(n781), .Z(n782) );
  NOR2_X1 U880 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U881 ( .A(KEYINPUT36), .B(n784), .ZN(n891) );
  NOR2_X1 U882 ( .A1(n817), .A2(n891), .ZN(n996) );
  INV_X1 U883 ( .A(n785), .ZN(n819) );
  NAND2_X1 U884 ( .A1(n996), .A2(n819), .ZN(n815) );
  NAND2_X1 U885 ( .A1(n786), .A2(n815), .ZN(n788) );
  XNOR2_X1 U886 ( .A(G1986), .B(G290), .ZN(n926) );
  AND2_X1 U887 ( .A1(n926), .A2(n819), .ZN(n787) );
  NOR2_X1 U888 ( .A1(n788), .A2(n787), .ZN(n791) );
  AND2_X1 U889 ( .A1(n937), .A2(n791), .ZN(n789) );
  NAND2_X1 U890 ( .A1(n790), .A2(n789), .ZN(n808) );
  INV_X1 U891 ( .A(n791), .ZN(n806) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n792) );
  XOR2_X1 U893 ( .A(n792), .B(KEYINPUT24), .Z(n793) );
  NOR2_X1 U894 ( .A1(n800), .A2(n793), .ZN(n804) );
  NOR2_X1 U895 ( .A1(G2090), .A2(G303), .ZN(n794) );
  XOR2_X1 U896 ( .A(KEYINPUT99), .B(n794), .Z(n795) );
  NAND2_X1 U897 ( .A1(G8), .A2(n795), .ZN(n799) );
  NAND2_X1 U898 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U900 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U901 ( .A(KEYINPUT100), .B(n802), .Z(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  OR2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  AND2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n822) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n866), .ZN(n989) );
  AND2_X1 U906 ( .A1(n1008), .A2(n865), .ZN(n975) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n809) );
  XOR2_X1 U908 ( .A(n809), .B(KEYINPUT101), .Z(n810) );
  NOR2_X1 U909 ( .A1(n975), .A2(n810), .ZN(n811) );
  NOR2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U911 ( .A1(n989), .A2(n813), .ZN(n814) );
  XNOR2_X1 U912 ( .A(n814), .B(KEYINPUT39), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n817), .A2(n891), .ZN(n993) );
  NAND2_X1 U915 ( .A1(n818), .A2(n993), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n825) );
  XOR2_X1 U918 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n823) );
  XNOR2_X1 U919 ( .A(KEYINPUT40), .B(n823), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n825), .B(n824), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U924 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U926 ( .A(n830), .ZN(G319) );
  XNOR2_X1 U927 ( .A(G1996), .B(G2474), .ZN(n840) );
  XOR2_X1 U928 ( .A(G1986), .B(G1991), .Z(n832) );
  XNOR2_X1 U929 ( .A(G1961), .B(G1956), .ZN(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U931 ( .A(G1966), .B(G1971), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1981), .B(G1976), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U934 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U935 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2090), .Z(n842) );
  XNOR2_X1 U939 ( .A(G2072), .B(G2084), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n843), .B(G2100), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2067), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U944 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U945 ( .A(KEYINPUT105), .B(G2678), .ZN(n846) );
  XNOR2_X1 U946 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U947 ( .A(n849), .B(n848), .Z(G227) );
  NAND2_X1 U948 ( .A1(G112), .A2(n877), .ZN(n856) );
  NAND2_X1 U949 ( .A1(G100), .A2(n880), .ZN(n851) );
  NAND2_X1 U950 ( .A1(G136), .A2(n881), .ZN(n850) );
  NAND2_X1 U951 ( .A1(n851), .A2(n850), .ZN(n854) );
  NAND2_X1 U952 ( .A1(n876), .A2(G124), .ZN(n852) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(n852), .Z(n853) );
  NOR2_X1 U954 ( .A1(n854), .A2(n853), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n857), .B(KEYINPUT107), .ZN(G162) );
  NAND2_X1 U957 ( .A1(G103), .A2(n880), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G139), .A2(n881), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G127), .A2(n876), .ZN(n861) );
  NAND2_X1 U961 ( .A1(G115), .A2(n877), .ZN(n860) );
  NAND2_X1 U962 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(KEYINPUT47), .B(n862), .Z(n863) );
  NOR2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n976) );
  XOR2_X1 U965 ( .A(n974), .B(n976), .Z(n868) );
  XOR2_X1 U966 ( .A(n866), .B(n865), .Z(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n875) );
  XOR2_X1 U968 ( .A(KEYINPUT48), .B(KEYINPUT109), .Z(n870) );
  XNOR2_X1 U969 ( .A(G164), .B(KEYINPUT110), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(n871), .B(KEYINPUT46), .Z(n873) );
  XNOR2_X1 U972 ( .A(G160), .B(KEYINPUT111), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U974 ( .A(n875), .B(n874), .Z(n890) );
  NAND2_X1 U975 ( .A1(G130), .A2(n876), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G118), .A2(n877), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n887) );
  NAND2_X1 U978 ( .A1(G106), .A2(n880), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G142), .A2(n881), .ZN(n882) );
  NAND2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U981 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  XNOR2_X1 U982 ( .A(KEYINPUT108), .B(n885), .ZN(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U984 ( .A(G162), .B(n888), .ZN(n889) );
  XNOR2_X1 U985 ( .A(n890), .B(n889), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n893) );
  NOR2_X1 U987 ( .A1(G37), .A2(n893), .ZN(G395) );
  XNOR2_X1 U988 ( .A(n894), .B(n922), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n895), .B(n925), .ZN(n897) );
  XNOR2_X1 U990 ( .A(G286), .B(G171), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(n899) );
  XNOR2_X1 U993 ( .A(KEYINPUT112), .B(n899), .ZN(G397) );
  XOR2_X1 U994 ( .A(G2438), .B(KEYINPUT104), .Z(n901) );
  XNOR2_X1 U995 ( .A(G2443), .B(G2430), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U997 ( .A(n902), .B(G2435), .Z(n904) );
  XNOR2_X1 U998 ( .A(G1341), .B(G1348), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1000 ( .A(G2451), .B(G2427), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G2454), .B(G2446), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1003 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1004 ( .A1(G14), .A2(n909), .ZN(n921) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n921), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  XNOR2_X1 U1011 ( .A(KEYINPUT113), .B(G225), .ZN(G308) );
  XNOR2_X1 U1013 ( .A(KEYINPUT80), .B(n915), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(G860), .A2(n916), .ZN(n917) );
  XOR2_X1 U1015 ( .A(n918), .B(n917), .Z(G145) );
  INV_X1 U1016 ( .A(G120), .ZN(G236) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1020 ( .A(G325), .ZN(G261) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  INV_X1 U1022 ( .A(n921), .ZN(G401) );
  XOR2_X1 U1023 ( .A(G16), .B(KEYINPUT56), .Z(n947) );
  XNOR2_X1 U1024 ( .A(G1341), .B(n922), .ZN(n945) );
  XNOR2_X1 U1025 ( .A(n957), .B(G171), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(n923), .B(KEYINPUT123), .ZN(n936) );
  XOR2_X1 U1027 ( .A(G1348), .B(KEYINPUT122), .Z(n924) );
  XNOR2_X1 U1028 ( .A(n925), .B(n924), .ZN(n929) );
  NOR2_X1 U1029 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(G1956), .B(n930), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(G1971), .A2(G303), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(G168), .B(G1966), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1038 ( .A(KEYINPUT57), .B(n939), .Z(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n1034) );
  XOR2_X1 U1043 ( .A(G16), .B(KEYINPUT124), .Z(n972) );
  XNOR2_X1 U1044 ( .A(G20), .B(n948), .ZN(n952) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G1341), .B(G19), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1049 ( .A(KEYINPUT59), .B(G1348), .Z(n953) );
  XNOR2_X1 U1050 ( .A(G4), .B(n953), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(KEYINPUT60), .B(n956), .ZN(n968) );
  XOR2_X1 U1053 ( .A(G1966), .B(G21), .Z(n959) );
  XNOR2_X1 U1054 ( .A(n957), .B(G5), .ZN(n958) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G1976), .B(G23), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G1971), .B(G22), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n963) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n962) );
  NAND2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n964), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(KEYINPUT61), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(n970), .B(KEYINPUT125), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT126), .B(n973), .ZN(n1032) );
  INV_X1 U1068 ( .A(KEYINPUT55), .ZN(n1000) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n987) );
  XNOR2_X1 U1070 ( .A(G2072), .B(n976), .ZN(n977) );
  XNOR2_X1 U1071 ( .A(n977), .B(KEYINPUT115), .ZN(n979) );
  XOR2_X1 U1072 ( .A(G2078), .B(G164), .Z(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1074 ( .A(KEYINPUT50), .B(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1076 ( .A(G2084), .B(G160), .Z(n983) );
  XNOR2_X1 U1077 ( .A(KEYINPUT114), .B(n983), .ZN(n984) );
  NOR2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n992) );
  XOR2_X1 U1080 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(KEYINPUT51), .B(n990), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT52), .B(KEYINPUT116), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n998), .B(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(G29), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(n1002), .B(KEYINPUT117), .ZN(n1030) );
  XNOR2_X1 U1091 ( .A(G32), .B(n1003), .ZN(n1005) );
  XOR2_X1 U1092 ( .A(G2067), .B(G26), .Z(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G33), .B(G2072), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1016) );
  XNOR2_X1 U1096 ( .A(n1008), .B(G25), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(G28), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT118), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(n1011), .B(G27), .Z(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT119), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1017), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(G34), .B(KEYINPUT120), .Z(n1019) );
  XNOR2_X1 U1105 ( .A(G2084), .B(KEYINPUT54), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(n1019), .B(n1018), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(G35), .B(G2090), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT55), .B(n1024), .ZN(n1026) );
  INV_X1 U1111 ( .A(G29), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(G11), .ZN(n1028) );
  XOR2_X1 U1114 ( .A(KEYINPUT121), .B(n1028), .Z(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .Z(n1036) );
  XNOR2_X1 U1119 ( .A(KEYINPUT127), .B(n1036), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

