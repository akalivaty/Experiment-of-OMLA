//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n598, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  AND3_X1   g032(.A1(new_n457), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n458));
  AOI21_X1  g033(.A(KEYINPUT70), .B1(new_n457), .B2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G101), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(new_n457), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(G137), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n460), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n473), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n465), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(G125), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n478), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(KEYINPUT68), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n472), .B1(new_n479), .B2(new_n486), .ZN(G160));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n467), .A2(G2105), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n467), .A2(new_n478), .ZN(new_n493));
  AOI211_X1 g068(.A(new_n490), .B(new_n492), .C1(G124), .C2(new_n493), .ZN(G162));
  NAND4_X1  g069(.A1(new_n469), .A2(KEYINPUT4), .A3(G138), .A4(new_n470), .ZN(new_n495));
  NAND2_X1  g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n469), .A2(G138), .A3(new_n470), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n482), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(new_n457), .B2(G114), .ZN(new_n503));
  NOR2_X1   g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT71), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(G114), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n506), .A2(new_n508), .A3(new_n509), .A4(G2104), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n499), .A2(new_n502), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(new_n518), .B1(new_n515), .B2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n522), .A2(G88), .B1(new_n524), .B2(G50), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(G166));
  NAND2_X1  g106(.A1(new_n524), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(G89), .B2(new_n522), .ZN(G168));
  AOI22_X1  g112(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n526), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n521), .A2(new_n540), .B1(new_n523), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT74), .B(G43), .Z(new_n545));
  OAI22_X1  g120(.A1(new_n521), .A2(new_n544), .B1(new_n523), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n519), .A2(G56), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n526), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  AOI22_X1  g131(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G91), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n557), .A2(new_n526), .B1(new_n558), .B2(new_n521), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n524), .A2(KEYINPUT9), .A3(G53), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n523), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND3_X1  g144(.A1(new_n520), .A2(G49), .A3(G543), .ZN(new_n570));
  XOR2_X1   g145(.A(new_n570), .B(KEYINPUT76), .Z(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n522), .A2(G87), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n526), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT77), .Z(new_n577));
  AOI22_X1  g152(.A1(new_n522), .A2(G86), .B1(new_n524), .B2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G305));
  XNOR2_X1  g154(.A(KEYINPUT78), .B(G85), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n522), .A2(new_n580), .B1(new_n524), .B2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n526), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n521), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n585), .A2(new_n588), .B1(G54), .B2(new_n524), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n519), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(KEYINPUT79), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(KEYINPUT79), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n591), .A2(G651), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n584), .B1(new_n595), .B2(G868), .ZN(G321));
  XNOR2_X1  g171(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g172(.A1(G286), .A2(G868), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G868), .B2(new_n565), .ZN(G280));
  XOR2_X1   g174(.A(G280), .B(KEYINPUT81), .Z(G297));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n595), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n595), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n491), .A2(G135), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n493), .A2(G123), .ZN(new_n608));
  OAI221_X1 g183(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n478), .C2(G111), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT83), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G2096), .ZN(new_n613));
  INV_X1    g188(.A(G2096), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n474), .B1(new_n458), .B2(new_n459), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XOR2_X1   g192(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n617), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n613), .A2(new_n615), .A3(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G2427), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n627), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G14), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n631), .A2(new_n634), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(KEYINPUT86), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT17), .Z(new_n647));
  INV_X1    g222(.A(new_n640), .ZN(new_n648));
  INV_X1    g223(.A(new_n639), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n642), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n641), .B1(new_n651), .B2(new_n639), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n645), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n614), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(G227));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT87), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1961), .B(G1966), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n658), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  INV_X1    g243(.A(G1981), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1991), .B(G1996), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT88), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  NOR2_X1   g250(.A1(G16), .A2(G22), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G166), .B2(G16), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(G1971), .Z(new_n678));
  NOR2_X1   g253(.A1(G6), .A2(G16), .ZN(new_n679));
  INV_X1    g254(.A(G305), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(G16), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT32), .B(G1981), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(G23), .B(G288), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT89), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n678), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(KEYINPUT34), .ZN(new_n690));
  MUX2_X1   g265(.A(G24), .B(G290), .S(G16), .Z(new_n691));
  INV_X1    g266(.A(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G25), .ZN(new_n695));
  OAI221_X1 g270(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n478), .C2(G107), .ZN(new_n696));
  INV_X1    g271(.A(new_n493), .ZN(new_n697));
  INV_X1    g272(.A(G119), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G131), .B2(new_n491), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n695), .B1(new_n700), .B2(new_n694), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n689), .A2(new_n690), .A3(new_n693), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT36), .ZN(new_n705));
  INV_X1    g280(.A(G16), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G4), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n595), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT90), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1348), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT25), .ZN(new_n711));
  NAND2_X1  g286(.A1(G103), .A2(G2104), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n485), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n478), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n713), .A2(new_n714), .B1(new_n491), .B2(G139), .ZN(new_n715));
  NAND2_X1  g290(.A1(G115), .A2(G2104), .ZN(new_n716));
  INV_X1    g291(.A(G127), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n482), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(new_n485), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT92), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(KEYINPUT92), .A3(new_n485), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n715), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G33), .B(new_n723), .S(G29), .Z(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT93), .Z(new_n725));
  INV_X1    g300(.A(G2072), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n694), .A2(G32), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n491), .A2(G141), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT94), .Z(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT26), .Z(new_n732));
  OAI21_X1  g307(.A(G105), .B1(new_n458), .B2(new_n459), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G129), .B2(new_n493), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n728), .B1(new_n737), .B2(new_n694), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT27), .B(G1996), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n725), .A2(new_n726), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT97), .B(KEYINPUT23), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n706), .A2(G20), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n565), .B2(new_n706), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n727), .A2(new_n740), .A3(new_n741), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n694), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n694), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT29), .B(G2090), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT31), .B(G11), .Z(new_n753));
  INV_X1    g328(.A(G28), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(KEYINPUT30), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT95), .ZN(new_n756));
  AOI21_X1  g331(.A(G29), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G168), .A2(new_n706), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n706), .B2(G21), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G27), .A2(G29), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G164), .B2(G29), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2078), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n752), .A2(new_n762), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n706), .A2(G5), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G171), .B2(new_n706), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n770), .C1(new_n694), .C2(new_n612), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n760), .A2(new_n761), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT96), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  INV_X1    g349(.A(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(G29), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n774), .B2(new_n775), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G160), .B2(new_n694), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n706), .A2(G19), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n550), .B2(new_n706), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1341), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n694), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT91), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  OAI221_X1 g361(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n478), .C2(G116), .ZN(new_n787));
  INV_X1    g362(.A(G128), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n697), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G140), .B2(new_n491), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n786), .B1(new_n790), .B2(new_n694), .ZN(new_n791));
  INV_X1    g366(.A(G2067), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n773), .A2(new_n780), .A3(new_n783), .A4(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n710), .A2(new_n748), .A3(new_n771), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n705), .A2(new_n795), .ZN(G150));
  INV_X1    g371(.A(G150), .ZN(G311));
  INV_X1    g372(.A(G93), .ZN(new_n798));
  INV_X1    g373(.A(G55), .ZN(new_n799));
  OAI22_X1  g374(.A1(new_n521), .A2(new_n798), .B1(new_n523), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n519), .A2(G67), .ZN(new_n801));
  NAND2_X1  g376(.A1(G80), .A2(G543), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n526), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n550), .B(new_n804), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT38), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n595), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n809));
  INV_X1    g384(.A(G860), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(KEYINPUT39), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n804), .A2(new_n810), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT37), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(G145));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n736), .B(G164), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n790), .B(KEYINPUT98), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n723), .A2(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT100), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(KEYINPUT100), .B2(new_n723), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(KEYINPUT100), .A3(new_n820), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n491), .A2(G142), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n493), .A2(G130), .ZN(new_n827));
  OAI221_X1 g402(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n478), .C2(G118), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n617), .B(new_n829), .Z(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(new_n700), .Z(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n816), .B1(new_n825), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g408(.A(KEYINPUT101), .B(new_n831), .C1(new_n823), .C2(new_n824), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n833), .A2(new_n834), .B1(new_n832), .B2(new_n825), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n611), .B(G160), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G162), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n825), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n839), .B2(new_n831), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n825), .A2(new_n832), .ZN(new_n841));
  AOI21_X1  g416(.A(G37), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n838), .A2(KEYINPUT102), .A3(new_n842), .ZN(new_n846));
  AND3_X1   g421(.A1(new_n845), .A2(KEYINPUT40), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT40), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(G395));
  NOR2_X1   g424(.A1(new_n804), .A2(G868), .ZN(new_n850));
  XNOR2_X1  g425(.A(G166), .B(G290), .ZN(new_n851));
  XNOR2_X1  g426(.A(G305), .B(G288), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT104), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT42), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n857), .B1(new_n853), .B2(KEYINPUT104), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n856), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n595), .A2(G299), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n594), .A2(new_n565), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT41), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(KEYINPUT103), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n860), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n864), .B1(new_n867), .B2(KEYINPUT41), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n603), .B(new_n805), .Z(new_n869));
  MUX2_X1   g444(.A(new_n863), .B(new_n868), .S(new_n869), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n859), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n859), .A2(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(G868), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n850), .B1(new_n874), .B2(KEYINPUT106), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(KEYINPUT106), .B2(new_n874), .ZN(G295));
  OAI21_X1  g451(.A(new_n875), .B1(KEYINPUT106), .B2(new_n874), .ZN(G331));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n878));
  NOR2_X1   g453(.A1(G301), .A2(KEYINPUT107), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n805), .B(new_n879), .Z(new_n880));
  AOI21_X1  g455(.A(G168), .B1(G301), .B2(KEYINPUT107), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n868), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(new_n862), .B2(new_n882), .ZN(new_n884));
  INV_X1    g459(.A(new_n853), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n887));
  AOI21_X1  g462(.A(G37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(KEYINPUT108), .A3(new_n885), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n882), .A2(KEYINPUT41), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n885), .B1(new_n891), .B2(new_n867), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n862), .B2(new_n891), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n884), .A2(new_n885), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n888), .A2(new_n897), .A3(new_n890), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n894), .A2(new_n895), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n878), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n889), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n888), .A2(new_n890), .A3(new_n893), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n889), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT44), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n906), .ZN(G397));
  INV_X1    g482(.A(G1384), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT45), .B1(new_n512), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n460), .B(G40), .C1(new_n467), .C2(new_n471), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n479), .B2(new_n486), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G1996), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n736), .B(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n790), .B(G2067), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n700), .A2(new_n702), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n700), .A2(new_n702), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(G290), .B(new_n692), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n912), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n908), .A2(KEYINPUT45), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n511), .A2(new_n502), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n467), .B1(new_n495), .B2(new_n496), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n911), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(new_n909), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n929), .A2(G1971), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n908), .B1(new_n925), .B2(new_n926), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT50), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n512), .A2(new_n933), .A3(new_n908), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n911), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(G2090), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n930), .B1(new_n936), .B2(KEYINPUT110), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(KEYINPUT110), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G8), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n529), .A2(G8), .A3(new_n530), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(KEYINPUT111), .B(G8), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n478), .A2(new_n474), .A3(G138), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n944), .A2(new_n500), .B1(new_n505), .B2(new_n510), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n945), .B2(new_n499), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n943), .B1(new_n911), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1976), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(G288), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT52), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT52), .B1(G288), .B2(new_n948), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n952), .B2(new_n949), .ZN(new_n953));
  INV_X1    g528(.A(new_n947), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n680), .A2(new_n669), .ZN(new_n955));
  NAND2_X1  g530(.A1(G305), .A2(G1981), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n955), .A2(KEYINPUT49), .A3(new_n956), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n953), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n943), .ZN(new_n962));
  INV_X1    g537(.A(new_n936), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(new_n930), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n941), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n942), .A2(new_n961), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT124), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(G168), .A2(new_n943), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n761), .B1(new_n928), .B2(new_n909), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT113), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n911), .B(new_n927), .C1(new_n946), .C2(KEYINPUT45), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT113), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n973), .A3(new_n761), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n932), .A2(new_n779), .A3(new_n934), .A4(new_n911), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n971), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n969), .B1(new_n976), .B2(G8), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT120), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n973), .B1(new_n972), .B2(new_n761), .ZN(new_n982));
  AND4_X1   g557(.A1(new_n779), .A2(new_n932), .A3(new_n911), .A4(new_n934), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n984), .B2(new_n974), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n980), .B(KEYINPUT51), .C1(new_n985), .C2(new_n969), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n976), .A2(new_n962), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n987), .B(new_n978), .C1(G168), .C2(new_n943), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n979), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT121), .ZN(new_n990));
  INV_X1    g565(.A(new_n987), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(G286), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n989), .B2(new_n992), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT62), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n992), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT121), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT62), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n989), .A2(new_n990), .A3(new_n992), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G2078), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n929), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT122), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n929), .A2(KEYINPUT122), .A3(new_n1001), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n1006), .A2(new_n1007), .B1(new_n769), .B2(new_n935), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1004), .B1(new_n1008), .B2(KEYINPUT123), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n935), .A2(new_n769), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n1010), .A2(KEYINPUT123), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(G171), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n995), .A2(new_n1000), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(G301), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT53), .B(new_n1001), .C1(new_n475), .C2(new_n478), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(new_n910), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n927), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1004), .B(new_n1011), .C1(new_n909), .C2(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1020), .A2(KEYINPUT125), .ZN(new_n1021));
  AOI21_X1  g596(.A(G301), .B1(new_n1020), .B2(KEYINPUT125), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1016), .A2(KEYINPUT54), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1020), .A2(G171), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(KEYINPUT54), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1013), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1348), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n935), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n911), .A2(new_n946), .A3(new_n792), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT60), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT60), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n594), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT58), .B(G1341), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n911), .B2(new_n946), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n1039));
  OAI22_X1  g614(.A1(new_n972), .A2(G1996), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n550), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g617(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1036), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n560), .A2(new_n1047), .A3(new_n563), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1047), .B1(new_n560), .B2(new_n563), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(new_n559), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT115), .B1(new_n1051), .B2(KEYINPUT57), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1050), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1048), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1053), .B(new_n1054), .C1(new_n1056), .C2(new_n559), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n565), .A2(KEYINPUT57), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1063));
  XNOR2_X1  g638(.A(new_n1063), .B(new_n726), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n929), .A2(new_n1064), .B1(new_n935), .B2(new_n746), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1068), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1067), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1071), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1046), .A2(new_n1069), .A3(new_n1070), .A4(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1031), .A2(new_n594), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1072), .B1(new_n1066), .B2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1024), .A2(new_n1027), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n994), .B2(new_n993), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n968), .B1(new_n1015), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT63), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n991), .A2(G168), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1081), .B1(new_n966), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n939), .A2(new_n941), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1082), .A2(new_n1081), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n942), .A2(new_n961), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n959), .A2(new_n960), .ZN(new_n1088));
  NOR2_X1   g663(.A1(G288), .A2(G1976), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1088), .A2(new_n1089), .B1(new_n669), .B2(new_n680), .ZN(new_n1090));
  INV_X1    g665(.A(new_n961), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1090), .A2(new_n954), .B1(new_n1091), .B2(new_n942), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1087), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n923), .B1(new_n1080), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n912), .B1(new_n915), .B2(new_n737), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT46), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n909), .A2(new_n913), .A3(new_n911), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1102));
  XOR2_X1   g677(.A(new_n1102), .B(KEYINPUT47), .Z(new_n1103));
  NOR2_X1   g678(.A1(new_n920), .A2(new_n912), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n912), .A2(G1986), .A3(G290), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(KEYINPUT48), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n917), .B(KEYINPUT126), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n916), .A2(new_n1107), .B1(new_n792), .B2(new_n790), .ZN(new_n1108));
  OAI22_X1  g683(.A1(new_n1104), .A2(new_n1106), .B1(new_n912), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1103), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1097), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT127), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1097), .A2(KEYINPUT127), .A3(new_n1110), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g690(.A1(new_n900), .A2(new_n901), .ZN(new_n1117));
  OAI21_X1  g691(.A(G319), .B1(new_n636), .B2(new_n637), .ZN(new_n1118));
  NOR3_X1   g692(.A1(G229), .A2(G227), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g693(.A(new_n846), .ZN(new_n1120));
  AOI21_X1  g694(.A(KEYINPUT102), .B1(new_n838), .B2(new_n842), .ZN(new_n1121));
  OAI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g696(.A1(new_n1117), .A2(new_n1122), .ZN(G308));
  OAI221_X1 g697(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .C1(new_n900), .C2(new_n901), .ZN(G225));
endmodule


