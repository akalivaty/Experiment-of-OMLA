

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773;

  XNOR2_X1 U379 ( .A(n383), .B(n671), .ZN(n672) );
  XNOR2_X1 U380 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X2 U381 ( .A1(n641), .A2(n434), .ZN(n433) );
  INV_X1 U382 ( .A(KEYINPUT70), .ZN(n356) );
  XNOR2_X2 U383 ( .A(n634), .B(KEYINPUT89), .ZN(n674) );
  NOR2_X1 U384 ( .A1(n613), .A2(n356), .ZN(n370) );
  XOR2_X1 U385 ( .A(n533), .B(KEYINPUT1), .Z(n357) );
  NAND2_X2 U386 ( .A1(n547), .A2(n375), .ZN(n408) );
  OR2_X2 U387 ( .A1(n363), .A2(n414), .ZN(n410) );
  AND2_X2 U388 ( .A1(n416), .A2(n412), .ZN(n411) );
  NAND2_X2 U389 ( .A1(n422), .A2(n369), .ZN(n399) );
  OR2_X2 U390 ( .A1(n660), .A2(G902), .ZN(n447) );
  NOR2_X2 U391 ( .A1(n716), .A2(n597), .ZN(n587) );
  OR2_X1 U392 ( .A1(n405), .A2(n358), .ZN(n716) );
  NOR2_X1 U393 ( .A1(G953), .A2(G237), .ZN(n477) );
  XNOR2_X1 U394 ( .A(n599), .B(n598), .ZN(n601) );
  NOR2_X1 U395 ( .A1(n424), .A2(n364), .ZN(n427) );
  NOR2_X1 U396 ( .A1(n726), .A2(n729), .ZN(n532) );
  XNOR2_X1 U397 ( .A(n405), .B(n404), .ZN(n421) );
  INV_X2 U398 ( .A(n586), .ZN(n358) );
  XNOR2_X1 U399 ( .A(n484), .B(n483), .ZN(n648) );
  NOR2_X1 U400 ( .A1(n606), .A2(n607), .ZN(n409) );
  NAND2_X1 U401 ( .A1(n367), .A2(n384), .ZN(n607) );
  NAND2_X1 U402 ( .A1(n601), .A2(n600), .ZN(n603) );
  OR2_X1 U403 ( .A1(n427), .A2(n430), .ZN(n395) );
  NAND2_X1 U404 ( .A1(n421), .A2(n594), .ZN(n420) );
  XNOR2_X1 U405 ( .A(n468), .B(n467), .ZN(n534) );
  NOR2_X2 U406 ( .A1(n648), .A2(G902), .ZN(n419) );
  XNOR2_X1 U407 ( .A(n475), .B(n454), .ZN(n761) );
  XNOR2_X1 U408 ( .A(KEYINPUT77), .B(KEYINPUT34), .ZN(n598) );
  OR2_X1 U409 ( .A1(n549), .A2(n414), .ZN(n359) );
  NAND2_X1 U410 ( .A1(n361), .A2(n362), .ZN(n360) );
  NAND2_X1 U411 ( .A1(n609), .A2(n381), .ZN(n361) );
  AND2_X1 U412 ( .A1(n615), .A2(n614), .ZN(n362) );
  XNOR2_X1 U413 ( .A(n587), .B(KEYINPUT31), .ZN(n695) );
  NOR2_X2 U414 ( .A1(n541), .A2(n540), .ZN(n550) );
  XNOR2_X1 U415 ( .A(n418), .B(n417), .ZN(n645) );
  NAND2_X1 U416 ( .A1(n411), .A2(n410), .ZN(n418) );
  XNOR2_X1 U417 ( .A(n560), .B(KEYINPUT1), .ZN(n585) );
  XNOR2_X1 U418 ( .A(n420), .B(KEYINPUT33), .ZN(n733) );
  XNOR2_X1 U419 ( .A(n619), .B(n618), .ZN(n627) );
  NOR2_X1 U420 ( .A1(n627), .A2(n622), .ZN(n397) );
  NAND2_X1 U421 ( .A1(n393), .A2(n390), .ZN(n363) );
  NAND2_X1 U422 ( .A1(n393), .A2(n390), .ZN(n544) );
  OR2_X2 U423 ( .A1(n383), .A2(n500), .ZN(n503) );
  XNOR2_X2 U424 ( .A(n497), .B(n442), .ZN(n475) );
  OR2_X1 U425 ( .A1(n530), .A2(n379), .ZN(n414) );
  INV_X1 U426 ( .A(KEYINPUT99), .ZN(n388) );
  NOR2_X1 U427 ( .A1(n639), .A2(KEYINPUT83), .ZN(n434) );
  XNOR2_X1 U428 ( .A(KEYINPUT67), .B(G101), .ZN(n476) );
  XNOR2_X1 U429 ( .A(n389), .B(n491), .ZN(n495) );
  XNOR2_X1 U430 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n491) );
  XNOR2_X1 U431 ( .A(KEYINPUT16), .B(G122), .ZN(n488) );
  INV_X1 U432 ( .A(G128), .ZN(n440) );
  XNOR2_X1 U433 ( .A(n515), .B(n514), .ZN(n631) );
  NAND2_X1 U434 ( .A1(n392), .A2(n391), .ZN(n390) );
  INV_X1 U435 ( .A(KEYINPUT85), .ZN(n381) );
  AND2_X1 U436 ( .A1(n386), .A2(n387), .ZN(n385) );
  INV_X1 U437 ( .A(n678), .ZN(n387) );
  OR2_X1 U438 ( .A1(n613), .A2(KEYINPUT66), .ZN(n384) );
  INV_X1 U439 ( .A(KEYINPUT69), .ZN(n407) );
  NAND2_X1 U440 ( .A1(n429), .A2(KEYINPUT30), .ZN(n428) );
  INV_X1 U441 ( .A(n535), .ZN(n431) );
  INV_X1 U442 ( .A(n375), .ZN(n429) );
  INV_X1 U443 ( .A(G953), .ZN(n492) );
  INV_X1 U444 ( .A(n530), .ZN(n723) );
  XNOR2_X1 U445 ( .A(G146), .B(G137), .ZN(n479) );
  XOR2_X1 U446 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n618) );
  XOR2_X1 U447 ( .A(G122), .B(G104), .Z(n510) );
  XNOR2_X1 U448 ( .A(G113), .B(G143), .ZN(n509) );
  XNOR2_X1 U449 ( .A(G131), .B(G140), .ZN(n504) );
  INV_X1 U450 ( .A(KEYINPUT79), .ZN(n620) );
  INV_X1 U451 ( .A(KEYINPUT100), .ZN(n404) );
  NAND2_X1 U452 ( .A1(G234), .A2(G237), .ZN(n470) );
  OR2_X1 U453 ( .A1(n552), .A2(n545), .ZN(n726) );
  INV_X1 U454 ( .A(G237), .ZN(n487) );
  INV_X1 U455 ( .A(G902), .ZN(n527) );
  INV_X1 U456 ( .A(G953), .ZN(n764) );
  XNOR2_X1 U457 ( .A(G119), .B(KEYINPUT24), .ZN(n456) );
  XNOR2_X1 U458 ( .A(G128), .B(G110), .ZN(n455) );
  XNOR2_X1 U459 ( .A(G116), .B(G107), .ZN(n519) );
  XOR2_X1 U460 ( .A(KEYINPUT7), .B(G122), .Z(n520) );
  XNOR2_X1 U461 ( .A(n499), .B(n498), .ZN(n383) );
  NAND2_X1 U462 ( .A1(n530), .A2(n379), .ZN(n415) );
  INV_X1 U463 ( .A(KEYINPUT0), .ZN(n398) );
  XOR2_X1 U464 ( .A(KEYINPUT62), .B(n648), .Z(n649) );
  NAND2_X1 U465 ( .A1(n570), .A2(n423), .ZN(n639) );
  INV_X1 U466 ( .A(KEYINPUT40), .ZN(n417) );
  NOR2_X1 U467 ( .A1(n568), .A2(n423), .ZN(n558) );
  NAND2_X1 U468 ( .A1(n372), .A2(n764), .ZN(n742) );
  AND2_X1 U469 ( .A1(n586), .A2(n373), .ZN(n364) );
  AND2_X1 U470 ( .A1(n733), .A2(n720), .ZN(n365) );
  XOR2_X1 U471 ( .A(n502), .B(KEYINPUT92), .Z(n366) );
  AND2_X1 U472 ( .A1(n604), .A2(n385), .ZN(n367) );
  NOR2_X1 U473 ( .A1(n710), .A2(n534), .ZN(n368) );
  NOR2_X1 U474 ( .A1(n357), .A2(n582), .ZN(n369) );
  AND2_X1 U475 ( .A1(n639), .A2(KEYINPUT83), .ZN(n371) );
  NOR2_X1 U476 ( .A1(n741), .A2(n365), .ZN(n372) );
  AND2_X1 U477 ( .A1(n375), .A2(n426), .ZN(n373) );
  NOR2_X1 U478 ( .A1(n707), .A2(n583), .ZN(n374) );
  NAND2_X1 U479 ( .A1(n501), .A2(G214), .ZN(n375) );
  AND2_X1 U480 ( .A1(n416), .A2(n415), .ZN(n376) );
  AND2_X1 U481 ( .A1(n357), .A2(n595), .ZN(n377) );
  AND2_X1 U482 ( .A1(n431), .A2(n428), .ZN(n378) );
  XNOR2_X1 U483 ( .A(KEYINPUT71), .B(KEYINPUT39), .ZN(n379) );
  XOR2_X1 U484 ( .A(n580), .B(KEYINPUT22), .Z(n380) );
  INV_X1 U485 ( .A(KEYINPUT76), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n603), .B(KEYINPUT35), .ZN(n609) );
  XNOR2_X1 U487 ( .A(n603), .B(n602), .ZN(n612) );
  NOR2_X1 U488 ( .A1(n743), .A2(n742), .ZN(n744) );
  AND2_X1 U489 ( .A1(n629), .A2(n705), .ZN(n382) );
  AND2_X2 U490 ( .A1(n629), .A2(n705), .ZN(n670) );
  XNOR2_X1 U491 ( .A(n761), .B(n446), .ZN(n660) );
  BUF_X1 U492 ( .A(n627), .Z(n745) );
  INV_X1 U493 ( .A(n588), .ZN(n392) );
  NAND2_X1 U494 ( .A1(n588), .A2(KEYINPUT76), .ZN(n394) );
  XNOR2_X2 U495 ( .A(n469), .B(KEYINPUT96), .ZN(n588) );
  XNOR2_X2 U496 ( .A(n584), .B(KEYINPUT86), .ZN(n613) );
  XNOR2_X1 U497 ( .A(n593), .B(n388), .ZN(n386) );
  XNOR2_X1 U498 ( .A(n461), .B(n389), .ZN(n759) );
  XNOR2_X2 U499 ( .A(G146), .B(G125), .ZN(n389) );
  AND2_X1 U500 ( .A1(n427), .A2(n430), .ZN(n391) );
  AND2_X2 U501 ( .A1(n394), .A2(n395), .ZN(n393) );
  NAND2_X1 U502 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U503 ( .A1(n397), .A2(n396), .ZN(n621) );
  XNOR2_X1 U504 ( .A(n700), .B(KEYINPUT74), .ZN(n396) );
  NAND2_X1 U505 ( .A1(n544), .A2(n379), .ZN(n416) );
  BUF_X1 U506 ( .A(n612), .Z(n644) );
  NAND2_X1 U507 ( .A1(n585), .A2(n368), .ZN(n405) );
  XNOR2_X1 U508 ( .A(n490), .B(n753), .ZN(n499) );
  INV_X1 U509 ( .A(n590), .ZN(n597) );
  NAND2_X1 U510 ( .A1(n590), .A2(n438), .ZN(n581) );
  XNOR2_X2 U511 ( .A(n577), .B(n398), .ZN(n590) );
  NAND2_X1 U512 ( .A1(n644), .A2(n370), .ZN(n611) );
  NAND2_X1 U513 ( .A1(n643), .A2(n640), .ZN(n584) );
  XNOR2_X2 U514 ( .A(n399), .B(KEYINPUT32), .ZN(n643) );
  XNOR2_X2 U515 ( .A(n581), .B(n380), .ZN(n422) );
  XNOR2_X2 U516 ( .A(n489), .B(n488), .ZN(n753) );
  XNOR2_X2 U517 ( .A(n401), .B(n400), .ZN(n489) );
  XNOR2_X2 U518 ( .A(G110), .B(KEYINPUT90), .ZN(n400) );
  XNOR2_X2 U519 ( .A(G107), .B(G104), .ZN(n401) );
  XNOR2_X2 U520 ( .A(n751), .B(n476), .ZN(n490) );
  XNOR2_X2 U521 ( .A(n403), .B(n402), .ZN(n751) );
  XNOR2_X2 U522 ( .A(KEYINPUT3), .B(G119), .ZN(n402) );
  XNOR2_X2 U523 ( .A(G116), .B(G113), .ZN(n403) );
  NOR2_X2 U524 ( .A1(n432), .A2(n436), .ZN(n700) );
  NOR2_X2 U525 ( .A1(n645), .A2(n773), .ZN(n543) );
  NAND2_X1 U526 ( .A1(n565), .A2(n406), .ZN(n567) );
  XNOR2_X1 U527 ( .A(n564), .B(n407), .ZN(n406) );
  XNOR2_X2 U528 ( .A(n408), .B(KEYINPUT19), .ZN(n576) );
  NAND2_X1 U529 ( .A1(n409), .A2(n617), .ZN(n619) );
  NOR2_X1 U530 ( .A1(n613), .A2(n609), .ZN(n605) );
  NAND2_X1 U531 ( .A1(n376), .A2(n359), .ZN(n571) );
  NOR2_X1 U532 ( .A1(n413), .A2(n692), .ZN(n412) );
  INV_X1 U533 ( .A(n415), .ZN(n413) );
  XNOR2_X2 U534 ( .A(n419), .B(n486), .ZN(n586) );
  NAND2_X1 U535 ( .A1(n733), .A2(n590), .ZN(n599) );
  NAND2_X1 U536 ( .A1(n422), .A2(n374), .ZN(n640) );
  AND2_X1 U537 ( .A1(n422), .A2(n377), .ZN(n678) );
  XNOR2_X1 U538 ( .A(n547), .B(KEYINPUT38), .ZN(n530) );
  INV_X1 U539 ( .A(n547), .ZN(n423) );
  XNOR2_X2 U540 ( .A(n503), .B(n366), .ZN(n547) );
  NAND2_X1 U541 ( .A1(n425), .A2(n378), .ZN(n424) );
  NAND2_X1 U542 ( .A1(n358), .A2(KEYINPUT30), .ZN(n425) );
  INV_X1 U543 ( .A(KEYINPUT30), .ZN(n426) );
  XNOR2_X1 U544 ( .A(n567), .B(n566), .ZN(n437) );
  NAND2_X1 U545 ( .A1(n437), .A2(n371), .ZN(n435) );
  NAND2_X1 U546 ( .A1(n435), .A2(n433), .ZN(n432) );
  NOR2_X1 U547 ( .A1(n437), .A2(KEYINPUT83), .ZN(n436) );
  BUF_X1 U548 ( .A(n560), .Z(n533) );
  AND2_X1 U549 ( .A1(n579), .A2(n578), .ZN(n438) );
  AND2_X1 U550 ( .A1(n610), .A2(KEYINPUT66), .ZN(n439) );
  XNOR2_X1 U551 ( .A(n513), .B(n512), .ZN(n514) );
  BUF_X1 U552 ( .A(n700), .Z(n763) );
  INV_X1 U553 ( .A(KEYINPUT41), .ZN(n531) );
  BUF_X1 U554 ( .A(n660), .Z(n665) );
  INV_X1 U555 ( .A(KEYINPUT60), .ZN(n636) );
  XNOR2_X2 U556 ( .A(G143), .B(KEYINPUT65), .ZN(n441) );
  XNOR2_X2 U557 ( .A(n441), .B(n440), .ZN(n524) );
  XNOR2_X2 U558 ( .A(n524), .B(KEYINPUT4), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G134), .B(G131), .ZN(n442) );
  XNOR2_X1 U560 ( .A(G140), .B(G137), .ZN(n454) );
  NAND2_X1 U561 ( .A1(n764), .A2(G227), .ZN(n443) );
  XNOR2_X1 U562 ( .A(n443), .B(G146), .ZN(n444) );
  XNOR2_X1 U563 ( .A(n444), .B(n476), .ZN(n445) );
  XNOR2_X1 U564 ( .A(n489), .B(n445), .ZN(n446) );
  XNOR2_X2 U565 ( .A(n447), .B(G469), .ZN(n560) );
  XNOR2_X2 U566 ( .A(G902), .B(KEYINPUT15), .ZN(n622) );
  NAND2_X1 U567 ( .A1(G234), .A2(n622), .ZN(n448) );
  XNOR2_X1 U568 ( .A(KEYINPUT20), .B(n448), .ZN(n451) );
  AND2_X1 U569 ( .A1(n451), .A2(G221), .ZN(n450) );
  INV_X1 U570 ( .A(KEYINPUT21), .ZN(n449) );
  XNOR2_X1 U571 ( .A(n450), .B(n449), .ZN(n710) );
  AND2_X1 U572 ( .A1(n451), .A2(G217), .ZN(n452) );
  XNOR2_X1 U573 ( .A(n452), .B(KEYINPUT95), .ZN(n453) );
  XNOR2_X1 U574 ( .A(n453), .B(KEYINPUT25), .ZN(n468) );
  XNOR2_X1 U575 ( .A(n455), .B(n454), .ZN(n459) );
  XOR2_X1 U576 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n457) );
  XNOR2_X1 U577 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U578 ( .A(n459), .B(n458), .ZN(n466) );
  INV_X1 U579 ( .A(KEYINPUT68), .ZN(n460) );
  XNOR2_X1 U580 ( .A(n460), .B(KEYINPUT10), .ZN(n461) );
  XOR2_X1 U581 ( .A(KEYINPUT78), .B(KEYINPUT8), .Z(n463) );
  NAND2_X1 U582 ( .A1(G234), .A2(n492), .ZN(n462) );
  XNOR2_X1 U583 ( .A(n463), .B(n462), .ZN(n518) );
  AND2_X1 U584 ( .A1(G221), .A2(n518), .ZN(n464) );
  XNOR2_X1 U585 ( .A(n759), .B(n464), .ZN(n465) );
  XNOR2_X1 U586 ( .A(n466), .B(n465), .ZN(n654) );
  NAND2_X1 U587 ( .A1(n654), .A2(n527), .ZN(n467) );
  NAND2_X1 U588 ( .A1(n560), .A2(n368), .ZN(n469) );
  XNOR2_X1 U589 ( .A(n470), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U590 ( .A1(G902), .A2(n473), .ZN(n572) );
  NOR2_X1 U591 ( .A1(G900), .A2(n572), .ZN(n471) );
  NAND2_X1 U592 ( .A1(G953), .A2(n471), .ZN(n472) );
  XNOR2_X1 U593 ( .A(n472), .B(KEYINPUT102), .ZN(n474) );
  NAND2_X1 U594 ( .A1(G952), .A2(n473), .ZN(n740) );
  OR2_X1 U595 ( .A1(n740), .A2(G953), .ZN(n574) );
  AND2_X1 U596 ( .A1(n474), .A2(n574), .ZN(n535) );
  INV_X1 U597 ( .A(n475), .ZN(n484) );
  INV_X1 U598 ( .A(n477), .ZN(n478) );
  XNOR2_X1 U599 ( .A(KEYINPUT75), .B(n478), .ZN(n511) );
  NAND2_X1 U600 ( .A1(n511), .A2(G210), .ZN(n481) );
  XNOR2_X1 U601 ( .A(n479), .B(KEYINPUT5), .ZN(n480) );
  XNOR2_X1 U602 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U603 ( .A(n490), .B(n482), .ZN(n483) );
  INV_X1 U604 ( .A(KEYINPUT72), .ZN(n485) );
  XNOR2_X1 U605 ( .A(n485), .B(G472), .ZN(n486) );
  NAND2_X1 U606 ( .A1(n527), .A2(n487), .ZN(n501) );
  NAND2_X1 U607 ( .A1(n492), .A2(G224), .ZN(n493) );
  XNOR2_X1 U608 ( .A(n493), .B(KEYINPUT91), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U610 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U611 ( .A(n622), .ZN(n500) );
  NAND2_X1 U612 ( .A1(n501), .A2(G210), .ZN(n502) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n508) );
  XOR2_X1 U614 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n505) );
  XNOR2_X1 U615 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U616 ( .A(n759), .B(n506), .ZN(n507) );
  XNOR2_X1 U617 ( .A(n508), .B(n507), .ZN(n515) );
  XOR2_X1 U618 ( .A(n510), .B(n509), .Z(n513) );
  NAND2_X1 U619 ( .A1(G214), .A2(n511), .ZN(n512) );
  NAND2_X1 U620 ( .A1(n631), .A2(n527), .ZN(n517) );
  XOR2_X1 U621 ( .A(KEYINPUT13), .B(G475), .Z(n516) );
  XNOR2_X1 U622 ( .A(n517), .B(n516), .ZN(n552) );
  AND2_X1 U623 ( .A1(n518), .A2(G217), .ZN(n523) );
  XNOR2_X1 U624 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U625 ( .A(n521), .B(KEYINPUT9), .Z(n522) );
  XNOR2_X1 U626 ( .A(n523), .B(n522), .ZN(n526) );
  XNOR2_X1 U627 ( .A(n524), .B(G134), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n526), .B(n525), .ZN(n658) );
  NAND2_X1 U629 ( .A1(n658), .A2(n527), .ZN(n529) );
  INV_X1 U630 ( .A(G478), .ZN(n528) );
  XNOR2_X1 U631 ( .A(n529), .B(n528), .ZN(n551) );
  NAND2_X1 U632 ( .A1(n552), .A2(n551), .ZN(n692) );
  INV_X1 U633 ( .A(n551), .ZN(n545) );
  NAND2_X1 U634 ( .A1(n723), .A2(n375), .ZN(n729) );
  XNOR2_X1 U635 ( .A(n532), .B(n531), .ZN(n720) );
  XNOR2_X1 U636 ( .A(n533), .B(KEYINPUT103), .ZN(n541) );
  BUF_X2 U637 ( .A(n534), .Z(n709) );
  NOR2_X1 U638 ( .A1(n710), .A2(n535), .ZN(n536) );
  NAND2_X1 U639 ( .A1(n709), .A2(n536), .ZN(n554) );
  NOR2_X1 U640 ( .A1(n358), .A2(n554), .ZN(n539) );
  XOR2_X1 U641 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n537) );
  XOR2_X1 U642 ( .A(n537), .B(KEYINPUT28), .Z(n538) );
  XNOR2_X1 U643 ( .A(n539), .B(n538), .ZN(n540) );
  NAND2_X1 U644 ( .A1(n720), .A2(n550), .ZN(n542) );
  XOR2_X1 U645 ( .A(KEYINPUT42), .B(n542), .Z(n773) );
  XNOR2_X1 U646 ( .A(n543), .B(KEYINPUT46), .ZN(n565) );
  BUF_X1 U647 ( .A(n363), .Z(n549) );
  NAND2_X1 U648 ( .A1(n552), .A2(n545), .ZN(n546) );
  XNOR2_X1 U649 ( .A(n546), .B(KEYINPUT101), .ZN(n600) );
  NAND2_X1 U650 ( .A1(n600), .A2(n547), .ZN(n548) );
  NOR2_X1 U651 ( .A1(n549), .A2(n548), .ZN(n638) );
  NAND2_X1 U652 ( .A1(n550), .A2(n576), .ZN(n690) );
  OR2_X1 U653 ( .A1(n552), .A2(n551), .ZN(n696) );
  AND2_X1 U654 ( .A1(n692), .A2(n696), .ZN(n728) );
  NOR2_X1 U655 ( .A1(n690), .A2(n728), .ZN(n553) );
  XNOR2_X1 U656 ( .A(n553), .B(KEYINPUT47), .ZN(n562) );
  XNOR2_X1 U657 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n559) );
  INV_X1 U658 ( .A(n554), .ZN(n555) );
  NAND2_X1 U659 ( .A1(n555), .A2(n375), .ZN(n556) );
  NOR2_X1 U660 ( .A1(n692), .A2(n556), .ZN(n557) );
  XNOR2_X1 U661 ( .A(n358), .B(KEYINPUT6), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n557), .A2(n594), .ZN(n568) );
  XOR2_X1 U663 ( .A(n559), .B(n558), .Z(n561) );
  INV_X1 U664 ( .A(n357), .ZN(n707) );
  NAND2_X1 U665 ( .A1(n561), .A2(n707), .ZN(n698) );
  NAND2_X1 U666 ( .A1(n562), .A2(n698), .ZN(n563) );
  NOR2_X1 U667 ( .A1(n638), .A2(n563), .ZN(n564) );
  INV_X1 U668 ( .A(KEYINPUT48), .ZN(n566) );
  NOR2_X1 U669 ( .A1(n707), .A2(n568), .ZN(n569) );
  XOR2_X1 U670 ( .A(KEYINPUT43), .B(n569), .Z(n570) );
  NOR2_X1 U671 ( .A1(n571), .A2(n696), .ZN(n641) );
  XNOR2_X1 U672 ( .A(G898), .B(KEYINPUT93), .ZN(n748) );
  NAND2_X1 U673 ( .A1(G953), .A2(n748), .ZN(n754) );
  OR2_X1 U674 ( .A1(n572), .A2(n754), .ZN(n573) );
  NAND2_X1 U675 ( .A1(n574), .A2(n573), .ZN(n575) );
  INV_X1 U676 ( .A(n726), .ZN(n579) );
  INV_X1 U677 ( .A(n710), .ZN(n578) );
  INV_X1 U678 ( .A(KEYINPUT73), .ZN(n580) );
  INV_X1 U679 ( .A(n594), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n596), .A2(n709), .ZN(n582) );
  NAND2_X1 U681 ( .A1(n358), .A2(n709), .ZN(n583) );
  NOR2_X1 U682 ( .A1(n588), .A2(n586), .ZN(n589) );
  NAND2_X1 U683 ( .A1(n590), .A2(n589), .ZN(n684) );
  NAND2_X1 U684 ( .A1(n695), .A2(n684), .ZN(n592) );
  INV_X1 U685 ( .A(n728), .ZN(n591) );
  NAND2_X1 U686 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U687 ( .A1(n594), .A2(n709), .ZN(n595) );
  INV_X1 U688 ( .A(KEYINPUT35), .ZN(n602) );
  NAND2_X1 U689 ( .A1(n612), .A2(KEYINPUT85), .ZN(n604) );
  NOR2_X1 U690 ( .A1(n605), .A2(KEYINPUT70), .ZN(n606) );
  NOR2_X1 U691 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n439), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n613), .A2(KEYINPUT66), .ZN(n615) );
  AND2_X1 U694 ( .A1(KEYINPUT70), .A2(KEYINPUT44), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n616), .A2(n360), .ZN(n617) );
  XNOR2_X1 U696 ( .A(n621), .B(n620), .ZN(n625) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT81), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n623), .A2(KEYINPUT2), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U700 ( .A1(n700), .A2(KEYINPUT2), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT82), .B(n626), .Z(n628) );
  INV_X1 U702 ( .A(n745), .ZN(n701) );
  NAND2_X1 U703 ( .A1(n628), .A2(n701), .ZN(n705) );
  NAND2_X1 U704 ( .A1(n670), .A2(G475), .ZN(n633) );
  XOR2_X1 U705 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n630) );
  XNOR2_X1 U706 ( .A(n633), .B(n632), .ZN(n635) );
  NOR2_X1 U707 ( .A1(n764), .A2(G952), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n674), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(G60) );
  XOR2_X1 U710 ( .A(G143), .B(n638), .Z(G45) );
  XNOR2_X1 U711 ( .A(n639), .B(G140), .ZN(G42) );
  XNOR2_X1 U712 ( .A(n640), .B(G110), .ZN(G12) );
  XOR2_X1 U713 ( .A(G134), .B(n641), .Z(G36) );
  XNOR2_X1 U714 ( .A(G119), .B(KEYINPUT126), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n643), .B(n642), .ZN(G21) );
  XNOR2_X1 U716 ( .A(n644), .B(G122), .ZN(G24) );
  BUF_X1 U717 ( .A(n645), .Z(n646) );
  XNOR2_X1 U718 ( .A(G131), .B(KEYINPUT127), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n646), .B(n647), .ZN(G33) );
  NAND2_X1 U720 ( .A1(n670), .A2(G472), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n651), .A2(n674), .ZN(n653) );
  XNOR2_X1 U723 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(G57) );
  NAND2_X1 U725 ( .A1(n382), .A2(G217), .ZN(n655) );
  XOR2_X1 U726 ( .A(n654), .B(n655), .Z(n656) );
  INV_X1 U727 ( .A(n674), .ZN(n668) );
  NOR2_X1 U728 ( .A1(n656), .A2(n668), .ZN(G66) );
  NAND2_X1 U729 ( .A1(n382), .A2(G478), .ZN(n657) );
  XOR2_X1 U730 ( .A(n658), .B(n657), .Z(n659) );
  NOR2_X1 U731 ( .A1(n659), .A2(n668), .ZN(G63) );
  NAND2_X1 U732 ( .A1(n382), .A2(G469), .ZN(n667) );
  XNOR2_X1 U733 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n661), .B(KEYINPUT117), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n662) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n667), .B(n666), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n669), .A2(n668), .ZN(G54) );
  NAND2_X1 U740 ( .A1(n670), .A2(G210), .ZN(n673) );
  XNOR2_X1 U741 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n675) );
  NAND2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n677) );
  XOR2_X1 U744 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n676) );
  XNOR2_X1 U745 ( .A(n677), .B(n676), .ZN(G51) );
  XOR2_X1 U746 ( .A(G101), .B(n678), .Z(G3) );
  NOR2_X1 U747 ( .A1(n684), .A2(n692), .ZN(n680) );
  XNOR2_X1 U748 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U750 ( .A(G104), .B(n681), .ZN(G6) );
  XOR2_X1 U751 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n683) );
  XNOR2_X1 U752 ( .A(G107), .B(KEYINPUT108), .ZN(n682) );
  XNOR2_X1 U753 ( .A(n683), .B(n682), .ZN(n686) );
  NOR2_X1 U754 ( .A1(n684), .A2(n696), .ZN(n685) );
  XOR2_X1 U755 ( .A(n686), .B(n685), .Z(G9) );
  NOR2_X1 U756 ( .A1(n690), .A2(n696), .ZN(n688) );
  XNOR2_X1 U757 ( .A(KEYINPUT109), .B(KEYINPUT29), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n688), .B(n687), .ZN(n689) );
  XOR2_X1 U759 ( .A(G128), .B(n689), .Z(G30) );
  NOR2_X1 U760 ( .A1(n690), .A2(n692), .ZN(n691) );
  XOR2_X1 U761 ( .A(G146), .B(n691), .Z(G48) );
  NOR2_X1 U762 ( .A1(n692), .A2(n695), .ZN(n693) );
  XOR2_X1 U763 ( .A(KEYINPUT110), .B(n693), .Z(n694) );
  XNOR2_X1 U764 ( .A(G113), .B(n694), .ZN(G15) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U766 ( .A(G116), .B(n697), .Z(G18) );
  XOR2_X1 U767 ( .A(G125), .B(n698), .Z(n699) );
  XNOR2_X1 U768 ( .A(n699), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U769 ( .A1(n763), .A2(n701), .ZN(n703) );
  INV_X1 U770 ( .A(KEYINPUT2), .ZN(n702) );
  NAND2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U773 ( .A(KEYINPUT80), .B(n706), .Z(n743) );
  NOR2_X1 U774 ( .A1(n368), .A2(n707), .ZN(n708) );
  XNOR2_X1 U775 ( .A(n708), .B(KEYINPUT50), .ZN(n715) );
  NAND2_X1 U776 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT111), .ZN(n712) );
  XNOR2_X1 U778 ( .A(KEYINPUT49), .B(n712), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n713), .A2(n358), .ZN(n714) );
  NOR2_X1 U780 ( .A1(n715), .A2(n714), .ZN(n718) );
  INV_X1 U781 ( .A(n716), .ZN(n717) );
  NOR2_X1 U782 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n719), .ZN(n721) );
  NAND2_X1 U784 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U785 ( .A(n722), .B(KEYINPUT112), .ZN(n736) );
  NOR2_X1 U786 ( .A1(n723), .A2(n375), .ZN(n724) );
  XOR2_X1 U787 ( .A(KEYINPUT113), .B(n724), .Z(n725) );
  NOR2_X1 U788 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U789 ( .A(n727), .B(KEYINPUT114), .ZN(n731) );
  NOR2_X1 U790 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U791 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U792 ( .A(KEYINPUT115), .B(n732), .ZN(n734) );
  NAND2_X1 U793 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U794 ( .A1(n736), .A2(n735), .ZN(n738) );
  XOR2_X1 U795 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n737) );
  XNOR2_X1 U796 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U797 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U798 ( .A(n744), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U799 ( .A1(n745), .A2(G953), .ZN(n750) );
  NAND2_X1 U800 ( .A1(G953), .A2(G224), .ZN(n746) );
  XOR2_X1 U801 ( .A(KEYINPUT61), .B(n746), .Z(n747) );
  NOR2_X1 U802 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n757) );
  XOR2_X1 U804 ( .A(n751), .B(G101), .Z(n752) );
  XNOR2_X1 U805 ( .A(n753), .B(n752), .ZN(n755) );
  NAND2_X1 U806 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U807 ( .A(n757), .B(n756), .Z(n758) );
  XNOR2_X1 U808 ( .A(KEYINPUT121), .B(n758), .ZN(G69) );
  XNOR2_X1 U809 ( .A(n759), .B(KEYINPUT122), .ZN(n760) );
  XNOR2_X1 U810 ( .A(n761), .B(n760), .ZN(n767) );
  XNOR2_X1 U811 ( .A(n767), .B(KEYINPUT123), .ZN(n762) );
  XNOR2_X1 U812 ( .A(n763), .B(n762), .ZN(n765) );
  NAND2_X1 U813 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U814 ( .A(KEYINPUT124), .B(n766), .ZN(n772) );
  XNOR2_X1 U815 ( .A(G227), .B(n767), .ZN(n768) );
  NAND2_X1 U816 ( .A1(n768), .A2(G900), .ZN(n769) );
  NAND2_X1 U817 ( .A1(n769), .A2(G953), .ZN(n770) );
  XOR2_X1 U818 ( .A(KEYINPUT125), .B(n770), .Z(n771) );
  NAND2_X1 U819 ( .A1(n772), .A2(n771), .ZN(G72) );
  XOR2_X1 U820 ( .A(G137), .B(n773), .Z(G39) );
endmodule

