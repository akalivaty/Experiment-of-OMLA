//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  NOR2_X1   g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT14), .ZN(new_n203));
  NAND2_X1  g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n204), .A2(KEYINPUT87), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(KEYINPUT87), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n203), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT15), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT14), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n202), .B(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(new_n205), .A3(new_n206), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n211), .B1(new_n209), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT88), .A2(G1gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(KEYINPUT16), .A3(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n225), .B(KEYINPUT89), .C1(G1gat), .C2(new_n224), .ZN(new_n226));
  INV_X1    g025(.A(G8gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n220), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(KEYINPUT17), .B1(new_n213), .B2(new_n219), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n209), .A2(new_n218), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n210), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n236), .A2(new_n237), .A3(new_n212), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n234), .A2(new_n238), .A3(new_n228), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT91), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT18), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n240), .B1(KEYINPUT90), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n229), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n239), .A2(new_n242), .A3(new_n243), .A4(new_n231), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n241), .ZN(new_n245));
  AND4_X1   g044(.A1(new_n245), .A2(new_n239), .A3(new_n243), .A4(new_n231), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n233), .B(new_n244), .C1(new_n246), .C2(new_n242), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G197gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT11), .ZN(new_n250));
  INV_X1    g049(.A(G169gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n247), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G230gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT10), .ZN(new_n258));
  XNOR2_X1  g057(.A(G57gat), .B(G64gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G71gat), .B(G78gat), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT95), .B(G85gat), .ZN(new_n264));
  INV_X1    g063(.A(G92gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(KEYINPUT7), .ZN(new_n268));
  INV_X1    g067(.A(G99gat), .ZN(new_n269));
  INV_X1    g068(.A(G106gat), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT8), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G99gat), .B(G106gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n266), .A2(new_n268), .A3(new_n273), .A4(new_n271), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n263), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(KEYINPUT96), .A3(new_n276), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT96), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n272), .A2(new_n279), .A3(new_n274), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n258), .B(new_n277), .C1(new_n281), .C2(new_n263), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT98), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n263), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n257), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G120gat), .B(G148gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT100), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(G176gat), .ZN(new_n290));
  INV_X1    g089(.A(G204gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n277), .B1(new_n281), .B2(new_n263), .ZN(new_n293));
  INV_X1    g092(.A(new_n257), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT99), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n287), .B(new_n298), .C1(new_n297), .C2(new_n296), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n294), .B1(new_n282), .B2(new_n284), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n292), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(G197gat), .A2(G204gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT22), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G211gat), .ZN(new_n306));
  INV_X1    g105(.A(G218gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n307), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT22), .ZN(new_n314));
  OAI22_X1  g113(.A1(new_n314), .A2(new_n308), .B1(new_n304), .B2(new_n303), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n305), .A2(new_n309), .A3(KEYINPUT69), .A4(new_n310), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  OAI21_X1  g118(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NOR3_X1   g120(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g122(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n318), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n319), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330));
  INV_X1    g129(.A(G176gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n251), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n329), .B1(new_n332), .B2(new_n320), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT64), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT64), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G190gat), .ZN(new_n337));
  AOI21_X1  g136(.A(G183gat), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT24), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n333), .B(KEYINPUT25), .C1(new_n338), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT27), .B(G183gat), .Z(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT64), .B(G190gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT28), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n335), .A2(new_n337), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT27), .B(G183gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OR3_X1    g151(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n319), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n348), .A2(new_n352), .A3(new_n339), .A4(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n345), .A2(KEYINPUT71), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT71), .B1(new_n345), .B2(new_n356), .ZN(new_n358));
  INV_X1    g157(.A(G226gat), .ZN(new_n359));
  INV_X1    g158(.A(G233gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NOR3_X1   g161(.A1(new_n357), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n356), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n361), .A2(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n317), .B1(new_n363), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n317), .B(KEYINPUT70), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n365), .B1(new_n357), .B2(new_n358), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n364), .A2(new_n362), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(G64gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(G92gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n368), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT37), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n368), .B2(new_n374), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT82), .B(KEYINPUT37), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n368), .A2(new_n374), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n374), .A3(KEYINPUT83), .A4(new_n381), .ZN(new_n385));
  AOI211_X1 g184(.A(new_n377), .B(new_n380), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT38), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n378), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n390));
  INV_X1    g189(.A(G148gat), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(G141gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(G141gat), .ZN(new_n393));
  INV_X1    g192(.A(G141gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G155gat), .A2(G162gat), .ZN(new_n397));
  INV_X1    g196(.A(G155gat), .ZN(new_n398));
  INV_X1    g197(.A(G162gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n397), .B1(new_n400), .B2(KEYINPUT2), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(G155gat), .A2(G162gat), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT73), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT73), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n400), .A2(new_n406), .A3(new_n397), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n394), .A2(G148gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n393), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n397), .A2(KEYINPUT2), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n405), .A2(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(new_n402), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  NOR3_X1   g212(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT73), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n406), .B1(new_n400), .B2(new_n397), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n401), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G120gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G113gat), .ZN(new_n421));
  INV_X1    g220(.A(G113gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G120gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT1), .ZN(new_n425));
  XNOR2_X1  g224(.A(G127gat), .B(G134gat), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(KEYINPUT65), .ZN(new_n427));
  INV_X1    g226(.A(G127gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(G134gat), .ZN(new_n429));
  INV_X1    g228(.A(G134gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G127gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(KEYINPUT65), .ZN(new_n433));
  XNOR2_X1  g232(.A(G113gat), .B(G120gat), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n432), .B(new_n433), .C1(new_n434), .C2(KEYINPUT1), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n427), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n412), .A2(new_n419), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n418), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n438), .A2(KEYINPUT4), .A3(new_n436), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n427), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n405), .A2(new_n407), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n442), .A2(new_n413), .B1(new_n396), .B2(new_n401), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n389), .B(new_n437), .C1(new_n439), .C2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT75), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n441), .B2(new_n443), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n450), .B1(new_n441), .B2(new_n443), .ZN(new_n451));
  INV_X1    g250(.A(new_n389), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n438), .A2(new_n449), .A3(new_n436), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT4), .B1(new_n438), .B2(new_n436), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n441), .A2(new_n440), .A3(new_n443), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(new_n389), .A3(new_n437), .A4(new_n446), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n448), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT0), .ZN(new_n461));
  XNOR2_X1  g260(.A(G57gat), .B(G85gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n463), .B(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n459), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n448), .A2(new_n466), .A3(new_n454), .A4(new_n458), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n470), .A2(new_n469), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n470), .A2(new_n469), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n474), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n384), .A2(new_n385), .ZN(new_n479));
  INV_X1    g278(.A(new_n365), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT71), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n364), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n345), .A2(KEYINPUT71), .A3(new_n356), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n369), .B1(new_n484), .B2(new_n372), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n361), .A3(new_n483), .ZN(new_n486));
  INV_X1    g285(.A(new_n317), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n366), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n379), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n377), .B(KEYINPUT72), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n489), .A2(KEYINPUT38), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n479), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n475), .A2(new_n478), .A3(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n388), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT79), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n487), .A2(new_n496), .A3(KEYINPUT29), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT29), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT79), .B1(new_n317), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n497), .A2(KEYINPUT3), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT80), .B1(new_n500), .B2(new_n443), .ZN(new_n501));
  INV_X1    g300(.A(G228gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(new_n360), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT80), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n499), .A2(KEYINPUT3), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n504), .B(new_n438), .C1(new_n505), .C2(new_n497), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n419), .A2(new_n498), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n370), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n501), .A2(new_n503), .A3(new_n506), .A4(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT31), .B(G50gat), .Z(new_n510));
  XNOR2_X1  g309(.A(G78gat), .B(G106gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT81), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(G22gat), .Z(new_n514));
  OR2_X1    g313(.A1(new_n512), .A2(KEYINPUT81), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT29), .B1(new_n311), .B2(new_n315), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n438), .B1(new_n516), .B2(KEYINPUT3), .ZN(new_n517));
  INV_X1    g316(.A(new_n507), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n317), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n519), .B1(new_n502), .B2(new_n360), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n509), .A2(new_n514), .A3(new_n515), .A4(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n509), .A2(new_n515), .A3(new_n520), .ZN(new_n522));
  INV_X1    g321(.A(new_n514), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n368), .A2(new_n374), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n490), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT30), .A3(new_n378), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n378), .A2(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n457), .A2(new_n437), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(new_n452), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(KEYINPUT39), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(new_n466), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n451), .A2(new_n453), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n530), .B(KEYINPUT39), .C1(new_n533), .C2(new_n452), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(KEYINPUT40), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n527), .A2(new_n528), .A3(new_n470), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT40), .B1(new_n532), .B2(new_n534), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n521), .B(new_n524), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT85), .B1(new_n495), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n527), .A2(new_n528), .B1(new_n471), .B2(new_n472), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n540), .B1(new_n521), .B2(new_n524), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT36), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n364), .A2(new_n436), .ZN(new_n543));
  NAND2_X1  g342(.A1(G227gat), .A2(G233gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n345), .A2(new_n441), .A3(new_n356), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT34), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n547), .B1(new_n544), .B2(KEYINPUT68), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n546), .B(new_n548), .Z(new_n549));
  AOI21_X1  g348(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(KEYINPUT33), .ZN(new_n551));
  XNOR2_X1  g350(.A(G15gat), .B(G43gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G71gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(new_n269), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT66), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n550), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n544), .ZN(new_n558));
  INV_X1    g357(.A(new_n545), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n441), .B1(new_n345), .B2(new_n356), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT66), .B1(new_n561), .B2(KEYINPUT32), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n551), .B(new_n554), .C1(new_n557), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT67), .ZN(new_n564));
  INV_X1    g363(.A(new_n554), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n555), .B1(new_n550), .B2(new_n556), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(KEYINPUT66), .A3(KEYINPUT32), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT67), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n551), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n554), .A2(KEYINPUT33), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n561), .A2(KEYINPUT32), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n549), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n549), .ZN(new_n576));
  AOI211_X1 g375(.A(new_n576), .B(new_n573), .C1(new_n564), .C2(new_n570), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n542), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT67), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n569), .B1(new_n568), .B2(new_n551), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n576), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n571), .A2(new_n574), .A3(new_n549), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n582), .A2(KEYINPUT36), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n541), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n538), .ZN(new_n586));
  INV_X1    g385(.A(new_n380), .ZN(new_n587));
  INV_X1    g386(.A(new_n377), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n479), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT38), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n590), .A2(new_n378), .A3(new_n591), .A4(new_n493), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT85), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n586), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n539), .A2(new_n585), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n524), .A2(new_n521), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n596), .A2(new_n582), .A3(new_n540), .A4(new_n583), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT35), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n575), .A2(new_n577), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT35), .ZN(new_n600));
  INV_X1    g399(.A(new_n591), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n596), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n527), .A2(new_n528), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n598), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n256), .B(new_n302), .C1(new_n595), .C2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n263), .A2(KEYINPUT21), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n263), .A2(KEYINPUT21), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n228), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n228), .B2(new_n608), .ZN(new_n611));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT20), .ZN(new_n617));
  XNOR2_X1  g416(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n615), .B(new_n619), .ZN(new_n620));
  OAI22_X1  g419(.A1(new_n213), .A2(new_n219), .B1(KEYINPUT97), .B2(KEYINPUT17), .ZN(new_n621));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n621), .A2(new_n281), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n281), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n234), .A2(new_n238), .A3(KEYINPUT97), .A4(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n626), .A3(new_n334), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n334), .B1(new_n624), .B2(new_n626), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n307), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(G190gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n632), .A2(G218gat), .A3(new_n627), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n630), .A2(new_n633), .A3(KEYINPUT94), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT93), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n630), .A2(new_n633), .A3(KEYINPUT94), .A4(new_n638), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n620), .A2(new_n642), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n606), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n473), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g446(.A1(new_n644), .A2(new_n604), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT16), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT42), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n649), .B2(KEYINPUT42), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n227), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(KEYINPUT42), .B2(new_n648), .ZN(G1325gat));
  AOI21_X1  g454(.A(G15gat), .B1(new_n644), .B2(new_n599), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n578), .A2(new_n584), .A3(G15gat), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n644), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n524), .A2(new_n521), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT43), .B(G22gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  NAND3_X1  g461(.A1(new_n606), .A2(new_n620), .A3(new_n642), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n663), .A2(G29gat), .A3(new_n473), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT45), .Z(new_n665));
  NAND2_X1  g464(.A1(new_n595), .A2(new_n605), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n642), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n620), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n302), .B(KEYINPUT102), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n640), .A2(new_n641), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n595), .B2(new_n605), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(KEYINPUT44), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n669), .A2(new_n255), .A3(new_n672), .A4(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n473), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n665), .A2(new_n677), .ZN(G1328gat));
  NOR3_X1   g477(.A1(new_n663), .A2(G36gat), .A3(new_n603), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT46), .ZN(new_n680));
  OAI21_X1  g479(.A(G36gat), .B1(new_n676), .B2(new_n603), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1329gat));
  NAND2_X1  g481(.A1(new_n578), .A2(new_n584), .ZN(new_n683));
  OAI21_X1  g482(.A(G43gat), .B1(new_n676), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n599), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n663), .A2(G43gat), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g487(.A(G50gat), .B1(new_n676), .B2(new_n596), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n596), .A2(G50gat), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n606), .A2(new_n620), .A3(new_n642), .A4(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT48), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT44), .B1(new_n666), .B2(new_n642), .ZN(new_n696));
  AOI211_X1 g495(.A(new_n668), .B(new_n673), .C1(new_n595), .C2(new_n605), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n698), .A2(new_n255), .A3(new_n659), .A4(new_n672), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n699), .A2(G50gat), .B1(KEYINPUT103), .B2(new_n691), .ZN(new_n700));
  INV_X1    g499(.A(new_n302), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n666), .A2(new_n620), .A3(new_n255), .A4(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n690), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n702), .A2(new_n673), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n693), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n695), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT103), .ZN(new_n708));
  AND4_X1   g507(.A1(new_n695), .A2(new_n689), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n694), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT105), .B(new_n694), .C1(new_n707), .C2(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1331gat));
  INV_X1    g513(.A(new_n671), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n715), .B1(new_n595), .B2(new_n605), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n620), .A2(new_n642), .A3(new_n255), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n645), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n603), .ZN(new_n722));
  NOR2_X1   g521(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n723));
  AND2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n722), .B2(new_n723), .ZN(G1333gat));
  NOR2_X1   g525(.A1(new_n718), .A2(new_n685), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n578), .A2(new_n584), .A3(G71gat), .ZN(new_n728));
  OAI22_X1  g527(.A1(new_n727), .A2(G71gat), .B1(new_n718), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT106), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g530(.A1(new_n719), .A2(new_n659), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n670), .A2(new_n255), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n674), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n737), .A2(KEYINPUT107), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n736), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n473), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n743), .A2(new_n264), .A3(new_n302), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n698), .A2(new_n302), .A3(new_n734), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n473), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n264), .B2(new_n746), .ZN(G1336gat));
  INV_X1    g546(.A(new_n745), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n265), .B1(new_n748), .B2(new_n604), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(KEYINPUT52), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n715), .A2(G92gat), .A3(new_n603), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n742), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n741), .B(KEYINPUT108), .Z(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n740), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n749), .B1(new_n756), .B2(new_n751), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n754), .B2(new_n757), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n745), .B2(new_n683), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n742), .A2(G99gat), .A3(new_n685), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n760), .B2(new_n701), .ZN(G1338gat));
  AOI21_X1  g560(.A(new_n270), .B1(new_n748), .B2(new_n659), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(KEYINPUT53), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n715), .A2(G106gat), .A3(new_n596), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n742), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n756), .B2(new_n764), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(G1339gat));
  NOR2_X1   g568(.A1(new_n247), .A2(new_n254), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n239), .A2(new_n243), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n771), .A2(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n252), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n302), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n282), .A2(new_n294), .A3(new_n284), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n287), .A2(KEYINPUT54), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  INV_X1    g579(.A(new_n292), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n300), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n780), .B1(new_n779), .B2(new_n783), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n299), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n774), .B1(new_n256), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n673), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n785), .A2(new_n786), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(new_n642), .A3(new_n299), .A4(new_n773), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n792), .A2(new_n620), .B1(new_n701), .B2(new_n717), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n685), .A2(new_n659), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n604), .A2(new_n473), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n256), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n255), .A2(new_n422), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT111), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n799), .B2(new_n802), .ZN(G1340gat));
  OAI21_X1  g602(.A(G120gat), .B1(new_n799), .B2(new_n715), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n798), .A2(new_n420), .A3(new_n302), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1341gat));
  NAND2_X1  g605(.A1(new_n798), .A2(new_n670), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g607(.A1(new_n798), .A2(new_n430), .A3(new_n642), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n642), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(G134gat), .ZN(new_n815));
  AOI211_X1 g614(.A(KEYINPUT112), .B(new_n430), .C1(new_n798), .C2(new_n642), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n811), .A2(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT113), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819));
  OAI221_X1 g618(.A(new_n819), .B1(new_n815), .B2(new_n816), .C1(new_n811), .C2(new_n812), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1343gat));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n792), .A2(new_n620), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n717), .A2(new_n701), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(KEYINPUT57), .A3(new_n659), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n793), .B2(new_n596), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n683), .A2(new_n797), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n255), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G141gat), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n825), .A2(new_n659), .ZN(new_n834));
  NOR4_X1   g633(.A1(new_n834), .A2(G141gat), .A3(new_n256), .A4(new_n830), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n822), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n830), .B1(new_n826), .B2(new_n828), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n394), .B1(new_n838), .B2(new_n255), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(KEYINPUT115), .A3(new_n835), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT58), .B1(new_n839), .B2(KEYINPUT114), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT115), .B1(new_n839), .B2(new_n835), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n833), .A2(new_n822), .A3(new_n836), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n833), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n843), .A2(new_n844), .B1(new_n846), .B2(KEYINPUT58), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n842), .A2(new_n847), .ZN(G1344gat));
  NOR2_X1   g647(.A1(new_n793), .A2(new_n596), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n830), .A2(new_n701), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n391), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n853), .B1(new_n673), .B2(new_n787), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n790), .A2(KEYINPUT116), .A3(new_n642), .A4(new_n299), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n773), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n789), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n789), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n620), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n596), .B1(new_n861), .B2(new_n824), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n826), .B1(new_n862), .B2(KEYINPUT57), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n850), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n391), .B1(new_n864), .B2(KEYINPUT118), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(new_n866), .A3(new_n850), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n852), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AOI211_X1 g667(.A(KEYINPUT59), .B(new_n391), .C1(new_n838), .C2(new_n302), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n851), .B1(new_n868), .B2(new_n869), .ZN(G1345gat));
  NOR2_X1   g669(.A1(new_n834), .A2(new_n830), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n670), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT119), .Z(new_n873));
  NOR2_X1   g672(.A1(new_n620), .A2(new_n398), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT120), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n873), .A2(new_n398), .B1(new_n838), .B2(new_n875), .ZN(G1346gat));
  AOI21_X1  g675(.A(new_n399), .B1(new_n838), .B2(new_n642), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n673), .A2(G162gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n871), .B2(new_n878), .ZN(new_n879));
  XOR2_X1   g678(.A(new_n879), .B(KEYINPUT121), .Z(G1347gat));
  NOR2_X1   g679(.A1(new_n645), .A2(new_n603), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT122), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n796), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n256), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n796), .A2(new_n881), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n251), .A3(new_n255), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n886), .B2(new_n302), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n715), .A2(new_n331), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n883), .B2(new_n890), .ZN(G1349gat));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n825), .A2(new_n670), .A3(new_n794), .A4(new_n882), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(KEYINPUT123), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n796), .A2(new_n895), .A3(new_n670), .A4(new_n882), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n896), .A3(G183gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n886), .A2(new_n670), .A3(new_n350), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n898), .A3(new_n892), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n900), .A2(KEYINPUT60), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT60), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n642), .A3(new_n349), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n883), .A2(new_n642), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(G190gat), .ZN(new_n908));
  AOI211_X1 g707(.A(KEYINPUT61), .B(new_n334), .C1(new_n883), .C2(new_n642), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n910), .B(new_n911), .ZN(G1351gat));
  AND3_X1   g711(.A1(new_n849), .A2(new_n683), .A3(new_n881), .ZN(new_n913));
  INV_X1    g712(.A(G197gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n255), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT126), .Z(new_n916));
  NAND3_X1  g715(.A1(new_n863), .A2(new_n683), .A3(new_n882), .ZN(new_n917));
  OAI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n256), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1352gat));
  NAND3_X1  g718(.A1(new_n913), .A2(new_n291), .A3(new_n302), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n913), .A2(new_n922), .A3(new_n291), .A4(new_n302), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n921), .A2(KEYINPUT62), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT62), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G204gat), .B1(new_n917), .B2(new_n715), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n913), .A2(new_n306), .A3(new_n670), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n863), .A2(new_n670), .A3(new_n683), .A4(new_n882), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n307), .A3(new_n673), .ZN(new_n934));
  AOI21_X1  g733(.A(G218gat), .B1(new_n913), .B2(new_n642), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(G1355gat));
endmodule


