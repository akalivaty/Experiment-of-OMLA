

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739;

  AND2_X1 U371 ( .A1(n541), .A2(n405), .ZN(n630) );
  XNOR2_X1 U372 ( .A(n443), .B(n444), .ZN(n715) );
  XNOR2_X2 U373 ( .A(n412), .B(KEYINPUT36), .ZN(n411) );
  NOR2_X2 U374 ( .A1(n630), .A2(n523), .ZN(n525) );
  XNOR2_X2 U375 ( .A(KEYINPUT38), .B(n540), .ZN(n648) );
  INV_X1 U376 ( .A(n521), .ZN(n633) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n503) );
  NOR2_X1 U378 ( .A1(n658), .A2(n376), .ZN(n584) );
  NOR2_X1 U379 ( .A1(n686), .A2(n685), .ZN(n687) );
  AND2_X2 U380 ( .A1(n381), .A2(n380), .ZN(n705) );
  NOR2_X1 U381 ( .A1(n537), .A2(n536), .ZN(n538) );
  AND2_X1 U382 ( .A1(n737), .A2(n738), .ZN(n551) );
  XNOR2_X1 U383 ( .A(n410), .B(KEYINPUT112), .ZN(n735) );
  XNOR2_X1 U384 ( .A(n542), .B(KEYINPUT39), .ZN(n559) );
  XNOR2_X1 U385 ( .A(n578), .B(n577), .ZN(n591) );
  NOR2_X1 U386 ( .A1(n658), .A2(n659), .ZN(n595) );
  XNOR2_X1 U387 ( .A(n471), .B(n470), .ZN(n544) );
  XNOR2_X1 U388 ( .A(n447), .B(n446), .ZN(n526) );
  XNOR2_X1 U389 ( .A(n460), .B(n459), .ZN(n543) );
  XOR2_X1 U390 ( .A(n696), .B(KEYINPUT59), .Z(n698) );
  XNOR2_X1 U391 ( .A(n409), .B(KEYINPUT84), .ZN(n609) );
  XNOR2_X1 U392 ( .A(G902), .B(KEYINPUT15), .ZN(n409) );
  XNOR2_X1 U393 ( .A(G137), .B(G131), .ZN(n494) );
  XNOR2_X2 U394 ( .A(n722), .B(n498), .ZN(n515) );
  NAND2_X1 U395 ( .A1(n541), .A2(n648), .ZN(n542) );
  NOR2_X1 U396 ( .A1(n641), .A2(n560), .ZN(n561) );
  INV_X1 U397 ( .A(KEYINPUT45), .ZN(n354) );
  AND2_X1 U398 ( .A1(n527), .A2(n416), .ZN(n398) );
  NAND2_X1 U399 ( .A1(n663), .A2(n662), .ZN(n659) );
  INV_X1 U400 ( .A(G472), .ZN(n390) );
  OR2_X2 U401 ( .A1(n614), .A2(G902), .ZN(n391) );
  BUF_X1 U402 ( .A(n612), .Z(n710) );
  INV_X1 U403 ( .A(n720), .ZN(n414) );
  INV_X1 U404 ( .A(KEYINPUT0), .ZN(n420) );
  INV_X1 U405 ( .A(KEYINPUT103), .ZN(n602) );
  NOR2_X1 U406 ( .A1(n601), .A2(n652), .ZN(n603) );
  XNOR2_X1 U407 ( .A(G119), .B(KEYINPUT5), .ZN(n500) );
  XOR2_X1 U408 ( .A(KEYINPUT70), .B(KEYINPUT93), .Z(n501) );
  INV_X1 U409 ( .A(G134), .ZN(n432) );
  XNOR2_X1 U410 ( .A(n493), .B(n417), .ZN(n527) );
  INV_X1 U411 ( .A(KEYINPUT67), .ZN(n417) );
  XNOR2_X1 U412 ( .A(n600), .B(n374), .ZN(n520) );
  INV_X1 U413 ( .A(KEYINPUT109), .ZN(n374) );
  NOR2_X1 U414 ( .A1(n694), .A2(G902), .ZN(n516) );
  XNOR2_X1 U415 ( .A(n389), .B(n402), .ZN(n663) );
  XNOR2_X1 U416 ( .A(n404), .B(n403), .ZN(n402) );
  NAND2_X1 U417 ( .A1(n401), .A2(n400), .ZN(n389) );
  INV_X1 U418 ( .A(KEYINPUT25), .ZN(n403) );
  INV_X1 U419 ( .A(n642), .ZN(n372) );
  XOR2_X1 U420 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n474) );
  XNOR2_X1 U421 ( .A(G137), .B(G128), .ZN(n472) );
  XOR2_X1 U422 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n453) );
  XNOR2_X1 U423 ( .A(KEYINPUT10), .B(G140), .ZN(n415) );
  XNOR2_X1 U424 ( .A(G131), .B(G143), .ZN(n449) );
  XOR2_X1 U425 ( .A(KEYINPUT95), .B(G104), .Z(n450) );
  XNOR2_X1 U426 ( .A(n455), .B(n385), .ZN(n384) );
  INV_X1 U427 ( .A(KEYINPUT96), .ZN(n385) );
  XNOR2_X1 U428 ( .A(G113), .B(G122), .ZN(n455) );
  INV_X1 U429 ( .A(KEYINPUT18), .ZN(n435) );
  NAND2_X1 U430 ( .A1(n595), .A2(n590), .ZN(n570) );
  XNOR2_X1 U431 ( .A(n369), .B(n611), .ZN(n613) );
  INV_X1 U432 ( .A(KEYINPUT79), .ZN(n611) );
  NAND2_X1 U433 ( .A1(n394), .A2(n349), .ZN(n393) );
  BUF_X1 U434 ( .A(n526), .Z(n558) );
  NOR2_X1 U435 ( .A1(n544), .A2(n543), .ZN(n571) );
  NOR2_X1 U436 ( .A1(n659), .A2(n530), .ZN(n600) );
  INV_X1 U437 ( .A(KEYINPUT89), .ZN(n428) );
  BUF_X1 U438 ( .A(n666), .Z(n370) );
  XNOR2_X1 U439 ( .A(n499), .B(n512), .ZN(n443) );
  XNOR2_X1 U440 ( .A(n439), .B(n463), .ZN(n444) );
  XNOR2_X1 U441 ( .A(n477), .B(n364), .ZN(n439) );
  INV_X1 U442 ( .A(KEYINPUT46), .ZN(n550) );
  OR2_X1 U443 ( .A1(n652), .A2(n627), .ZN(n535) );
  INV_X1 U444 ( .A(KEYINPUT82), .ZN(n357) );
  NAND2_X1 U445 ( .A1(n606), .A2(n605), .ZN(n358) );
  NAND2_X1 U446 ( .A1(G237), .A2(G234), .ZN(n485) );
  XOR2_X1 U447 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n486) );
  OR2_X1 U448 ( .A1(G902), .A2(G237), .ZN(n508) );
  NAND2_X1 U449 ( .A1(n395), .A2(KEYINPUT108), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n515), .B(n506), .ZN(n614) );
  XNOR2_X1 U451 ( .A(n365), .B(KEYINPUT68), .ZN(n364) );
  INV_X1 U452 ( .A(KEYINPUT16), .ZN(n365) );
  INV_X1 U453 ( .A(G146), .ZN(n498) );
  NOR2_X1 U454 ( .A1(n643), .A2(KEYINPUT2), .ZN(n644) );
  XNOR2_X1 U455 ( .A(n528), .B(n360), .ZN(n529) );
  XNOR2_X1 U456 ( .A(KEYINPUT110), .B(KEYINPUT28), .ZN(n360) );
  XNOR2_X1 U457 ( .A(n546), .B(n545), .ZN(n682) );
  AND2_X1 U458 ( .A1(n520), .A2(n519), .ZN(n408) );
  INV_X1 U459 ( .A(KEYINPUT30), .ZN(n407) );
  BUF_X1 U460 ( .A(n663), .Z(n376) );
  AND2_X1 U461 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U462 ( .A(n413), .B(n481), .ZN(n707) );
  XNOR2_X1 U463 ( .A(n467), .B(n387), .ZN(n701) );
  XNOR2_X1 U464 ( .A(n469), .B(n351), .ZN(n387) );
  XNOR2_X1 U465 ( .A(n454), .B(n384), .ZN(n456) );
  NAND2_X1 U466 ( .A1(n371), .A2(n353), .ZN(n381) );
  XNOR2_X1 U467 ( .A(n515), .B(n429), .ZN(n694) );
  XNOR2_X1 U468 ( .A(n431), .B(n430), .ZN(n429) );
  XNOR2_X1 U469 ( .A(n514), .B(n513), .ZN(n430) );
  XNOR2_X1 U470 ( .A(n511), .B(n512), .ZN(n431) );
  XNOR2_X1 U471 ( .A(n437), .B(n445), .ZN(n425) );
  NOR2_X1 U472 ( .A1(G952), .A2(n728), .ZN(n709) );
  NAND2_X1 U473 ( .A1(n399), .A2(n396), .ZN(n555) );
  AND2_X1 U474 ( .A1(n392), .A2(n399), .ZN(n412) );
  INV_X1 U475 ( .A(KEYINPUT34), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n424), .B(n422), .ZN(n733) );
  XNOR2_X1 U477 ( .A(n588), .B(n423), .ZN(n422) );
  OR2_X1 U478 ( .A1(n591), .A2(n587), .ZN(n424) );
  INV_X1 U479 ( .A(KEYINPUT32), .ZN(n423) );
  AND2_X1 U480 ( .A1(n571), .A2(n558), .ZN(n405) );
  NOR2_X1 U481 ( .A1(n368), .A2(n370), .ZN(n367) );
  INV_X1 U482 ( .A(n600), .ZN(n368) );
  INV_X1 U483 ( .A(KEYINPUT53), .ZN(n377) );
  AND2_X1 U484 ( .A1(n558), .A2(n647), .ZN(n349) );
  NAND2_X1 U485 ( .A1(n394), .A2(n647), .ZN(n350) );
  INV_X1 U486 ( .A(n558), .ZN(n540) );
  XOR2_X1 U487 ( .A(n462), .B(n461), .Z(n351) );
  OR2_X1 U488 ( .A1(n607), .A2(KEYINPUT44), .ZN(n352) );
  NAND2_X1 U489 ( .A1(G214), .A2(n508), .ZN(n647) );
  INV_X1 U490 ( .A(KEYINPUT108), .ZN(n416) );
  OR2_X1 U491 ( .A1(n610), .A2(n609), .ZN(n353) );
  XNOR2_X2 U492 ( .A(n355), .B(n354), .ZN(n612) );
  NAND2_X1 U493 ( .A1(n356), .A2(n352), .ZN(n355) );
  XNOR2_X1 U494 ( .A(n358), .B(n357), .ZN(n356) );
  XNOR2_X1 U495 ( .A(n715), .B(n359), .ZN(n688) );
  XNOR2_X1 U496 ( .A(n438), .B(n425), .ZN(n359) );
  INV_X1 U497 ( .A(n645), .ZN(n380) );
  INV_X2 U498 ( .A(n440), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n697), .B(n698), .ZN(n699) );
  XNOR2_X1 U500 ( .A(n361), .B(KEYINPUT124), .ZN(G66) );
  NOR2_X2 U501 ( .A1(n708), .A2(n709), .ZN(n361) );
  XNOR2_X1 U502 ( .A(n362), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U503 ( .A1(n691), .A2(n709), .ZN(n362) );
  XNOR2_X1 U504 ( .A(n363), .B(KEYINPUT19), .ZN(n569) );
  NAND2_X1 U505 ( .A1(n526), .A2(n647), .ZN(n363) );
  XNOR2_X2 U506 ( .A(KEYINPUT3), .B(G116), .ZN(n441) );
  XNOR2_X1 U507 ( .A(n576), .B(n428), .ZN(n599) );
  XNOR2_X2 U508 ( .A(n442), .B(n441), .ZN(n499) );
  NAND2_X1 U509 ( .A1(n705), .A2(G217), .ZN(n706) );
  INV_X1 U510 ( .A(G902), .ZN(n400) );
  XNOR2_X1 U511 ( .A(n375), .B(KEYINPUT40), .ZN(n737) );
  NOR2_X2 U512 ( .A1(n612), .A2(n609), .ZN(n608) );
  XNOR2_X1 U513 ( .A(n366), .B(n618), .ZN(G57) );
  NOR2_X2 U514 ( .A1(n617), .A2(n709), .ZN(n366) );
  AND2_X1 U515 ( .A1(n599), .A2(n367), .ZN(n624) );
  XNOR2_X1 U516 ( .A(n608), .B(KEYINPUT78), .ZN(n373) );
  NOR2_X2 U517 ( .A1(n699), .A2(n709), .ZN(n700) );
  INV_X1 U518 ( .A(n517), .ZN(n666) );
  XNOR2_X2 U519 ( .A(n391), .B(n390), .ZN(n517) );
  XNOR2_X1 U520 ( .A(n518), .B(n407), .ZN(n406) );
  NAND2_X1 U521 ( .A1(n559), .A2(n633), .ZN(n375) );
  NAND2_X1 U522 ( .A1(n726), .A2(KEYINPUT2), .ZN(n369) );
  NAND2_X1 U523 ( .A1(n373), .A2(n372), .ZN(n371) );
  INV_X1 U524 ( .A(n707), .ZN(n401) );
  XNOR2_X1 U525 ( .A(n378), .B(n377), .ZN(G75) );
  NAND2_X1 U526 ( .A1(n388), .A2(n728), .ZN(n378) );
  NOR2_X1 U527 ( .A1(n642), .A2(n612), .ZN(n643) );
  NOR2_X1 U528 ( .A1(n732), .A2(n734), .ZN(n589) );
  XNOR2_X2 U529 ( .A(n530), .B(KEYINPUT1), .ZN(n658) );
  INV_X2 U530 ( .A(G128), .ZN(n382) );
  NAND2_X1 U531 ( .A1(n688), .A2(n609), .ZN(n447) );
  XNOR2_X1 U532 ( .A(n573), .B(KEYINPUT35), .ZN(n732) );
  XNOR2_X1 U533 ( .A(n427), .B(n426), .ZN(n572) );
  INV_X2 U534 ( .A(n379), .ZN(n477) );
  XNOR2_X2 U535 ( .A(G110), .B(G119), .ZN(n379) );
  XNOR2_X1 U536 ( .A(n464), .B(KEYINPUT4), .ZN(n434) );
  XNOR2_X2 U537 ( .A(n382), .B(G143), .ZN(n464) );
  XNOR2_X1 U538 ( .A(n383), .B(KEYINPUT77), .ZN(n523) );
  NAND2_X1 U539 ( .A1(n652), .A2(KEYINPUT47), .ZN(n383) );
  XNOR2_X2 U540 ( .A(n666), .B(KEYINPUT106), .ZN(n580) );
  NOR2_X1 U541 ( .A1(n696), .A2(G902), .ZN(n460) );
  XNOR2_X1 U542 ( .A(n692), .B(n386), .ZN(n695) );
  XNOR2_X1 U543 ( .A(n694), .B(n693), .ZN(n386) );
  AND2_X2 U544 ( .A1(n408), .A2(n406), .ZN(n541) );
  XNOR2_X1 U545 ( .A(n687), .B(KEYINPUT122), .ZN(n388) );
  XNOR2_X1 U546 ( .A(n476), .B(n414), .ZN(n413) );
  NOR2_X1 U547 ( .A1(n646), .A2(n645), .ZN(n686) );
  XNOR2_X2 U548 ( .A(n517), .B(n507), .ZN(n590) );
  OR2_X1 U549 ( .A1(n418), .A2(n416), .ZN(n399) );
  NOR2_X1 U550 ( .A1(n397), .A2(n393), .ZN(n392) );
  AND2_X1 U551 ( .A1(n418), .A2(n398), .ZN(n397) );
  INV_X1 U552 ( .A(n527), .ZN(n395) );
  NOR2_X1 U553 ( .A1(n397), .A2(n350), .ZN(n396) );
  NAND2_X1 U554 ( .A1(n483), .A2(G217), .ZN(n404) );
  NAND2_X1 U555 ( .A1(n411), .A2(n579), .ZN(n410) );
  XNOR2_X2 U556 ( .A(n448), .B(n415), .ZN(n720) );
  NOR2_X1 U557 ( .A1(n521), .A2(n419), .ZN(n418) );
  INV_X1 U558 ( .A(n590), .ZN(n419) );
  XNOR2_X2 U559 ( .A(n421), .B(n420), .ZN(n576) );
  NAND2_X1 U560 ( .A1(n569), .A2(n568), .ZN(n421) );
  INV_X1 U561 ( .A(n576), .ZN(n596) );
  INV_X1 U562 ( .A(n681), .ZN(n655) );
  NAND2_X1 U563 ( .A1(n599), .A2(n681), .ZN(n427) );
  XNOR2_X2 U564 ( .A(n570), .B(KEYINPUT33), .ZN(n681) );
  XNOR2_X2 U565 ( .A(n497), .B(n496), .ZN(n722) );
  XNOR2_X2 U566 ( .A(n464), .B(n432), .ZN(n497) );
  XOR2_X2 U567 ( .A(G125), .B(G146), .Z(n448) );
  NOR2_X1 U568 ( .A1(n663), .A2(n492), .ZN(n493) );
  XNOR2_X1 U569 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n433) );
  INV_X1 U570 ( .A(KEYINPUT75), .ZN(n524) );
  XNOR2_X1 U571 ( .A(n436), .B(n435), .ZN(n437) );
  INV_X1 U572 ( .A(n640), .ZN(n560) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U574 ( .A(KEYINPUT41), .ZN(n545) );
  XNOR2_X1 U575 ( .A(n458), .B(G475), .ZN(n459) );
  XNOR2_X1 U576 ( .A(n614), .B(KEYINPUT62), .ZN(n615) );
  INV_X2 U577 ( .A(G953), .ZN(n728) );
  XNOR2_X1 U578 ( .A(n434), .B(n448), .ZN(n438) );
  AND2_X1 U579 ( .A1(G224), .A2(n728), .ZN(n436) );
  XOR2_X1 U580 ( .A(G107), .B(G122), .Z(n463) );
  XNOR2_X2 U581 ( .A(G101), .B(G113), .ZN(n440) );
  XOR2_X1 U582 ( .A(KEYINPUT85), .B(G104), .Z(n512) );
  XOR2_X1 U583 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n445) );
  AND2_X1 U584 ( .A1(G210), .A2(n508), .ZN(n446) );
  XNOR2_X1 U585 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U586 ( .A(n720), .B(n451), .ZN(n457) );
  NAND2_X1 U587 ( .A1(G214), .A2(n503), .ZN(n452) );
  XNOR2_X1 U588 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U589 ( .A(n457), .B(n456), .ZN(n696) );
  XNOR2_X1 U590 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n458) );
  XOR2_X1 U591 ( .A(KEYINPUT98), .B(n543), .Z(n522) );
  XNOR2_X1 U592 ( .A(KEYINPUT102), .B(G478), .ZN(n471) );
  XOR2_X1 U593 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n462) );
  XNOR2_X1 U594 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n461) );
  XOR2_X1 U595 ( .A(KEYINPUT101), .B(n463), .Z(n466) );
  XNOR2_X1 U596 ( .A(n497), .B(G116), .ZN(n465) );
  XNOR2_X1 U597 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U598 ( .A1(G234), .A2(n728), .ZN(n468) );
  XOR2_X1 U599 ( .A(KEYINPUT8), .B(n468), .Z(n478) );
  NAND2_X1 U600 ( .A1(G217), .A2(n478), .ZN(n469) );
  NOR2_X1 U601 ( .A1(G902), .A2(n701), .ZN(n470) );
  NAND2_X1 U602 ( .A1(n522), .A2(n544), .ZN(n521) );
  XOR2_X1 U603 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n473) );
  XNOR2_X1 U604 ( .A(n473), .B(n472), .ZN(n475) );
  XOR2_X1 U605 ( .A(n477), .B(KEYINPUT71), .Z(n480) );
  NAND2_X1 U606 ( .A1(G221), .A2(n478), .ZN(n479) );
  XNOR2_X1 U607 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U608 ( .A1(n609), .A2(G234), .ZN(n482) );
  XNOR2_X1 U609 ( .A(n482), .B(KEYINPUT20), .ZN(n483) );
  NAND2_X1 U610 ( .A1(n483), .A2(G221), .ZN(n484) );
  XOR2_X1 U611 ( .A(KEYINPUT21), .B(n484), .Z(n662) );
  XNOR2_X1 U612 ( .A(n486), .B(n485), .ZN(n488) );
  NAND2_X1 U613 ( .A1(G952), .A2(n488), .ZN(n679) );
  NOR2_X1 U614 ( .A1(G953), .A2(n679), .ZN(n487) );
  XOR2_X1 U615 ( .A(KEYINPUT87), .B(n487), .Z(n567) );
  INV_X1 U616 ( .A(n567), .ZN(n491) );
  NAND2_X1 U617 ( .A1(G902), .A2(n488), .ZN(n563) );
  NOR2_X1 U618 ( .A1(G900), .A2(n563), .ZN(n489) );
  NAND2_X1 U619 ( .A1(G953), .A2(n489), .ZN(n490) );
  NAND2_X1 U620 ( .A1(n491), .A2(n490), .ZN(n519) );
  NAND2_X1 U621 ( .A1(n662), .A2(n519), .ZN(n492) );
  XNOR2_X1 U622 ( .A(KEYINPUT6), .B(KEYINPUT104), .ZN(n507) );
  XOR2_X1 U623 ( .A(KEYINPUT4), .B(KEYINPUT66), .Z(n495) );
  XNOR2_X1 U624 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U625 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U626 ( .A(n499), .B(n502), .Z(n505) );
  NAND2_X1 U627 ( .A1(n503), .A2(G210), .ZN(n504) );
  XNOR2_X1 U628 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U629 ( .A(KEYINPUT72), .B(KEYINPUT90), .ZN(n514) );
  XOR2_X1 U630 ( .A(G107), .B(G101), .Z(n510) );
  XNOR2_X1 U631 ( .A(G110), .B(G140), .ZN(n509) );
  XNOR2_X1 U632 ( .A(n510), .B(n509), .ZN(n511) );
  NAND2_X1 U633 ( .A1(G227), .A2(n728), .ZN(n513) );
  XNOR2_X2 U634 ( .A(n516), .B(G469), .ZN(n530) );
  INV_X1 U635 ( .A(n658), .ZN(n579) );
  XNOR2_X1 U636 ( .A(n735), .B(KEYINPUT80), .ZN(n539) );
  NAND2_X1 U637 ( .A1(n580), .A2(n647), .ZN(n518) );
  NOR2_X1 U638 ( .A1(n544), .A2(n522), .ZN(n636) );
  NOR2_X2 U639 ( .A1(n633), .A2(n636), .ZN(n652) );
  XNOR2_X1 U640 ( .A(n525), .B(n524), .ZN(n533) );
  BUF_X1 U641 ( .A(n569), .Z(n531) );
  NAND2_X1 U642 ( .A1(n580), .A2(n527), .ZN(n528) );
  NOR2_X1 U643 ( .A1(n530), .A2(n529), .ZN(n547) );
  NAND2_X1 U644 ( .A1(n531), .A2(n547), .ZN(n627) );
  NAND2_X1 U645 ( .A1(n627), .A2(KEYINPUT47), .ZN(n532) );
  NAND2_X1 U646 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U647 ( .A(n534), .B(KEYINPUT76), .ZN(n537) );
  NOR2_X1 U648 ( .A1(KEYINPUT47), .A2(n535), .ZN(n536) );
  NAND2_X1 U649 ( .A1(n539), .A2(n538), .ZN(n553) );
  XOR2_X1 U650 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n549) );
  NAND2_X1 U651 ( .A1(n544), .A2(n543), .ZN(n650) );
  NAND2_X1 U652 ( .A1(n648), .A2(n647), .ZN(n651) );
  NOR2_X1 U653 ( .A1(n650), .A2(n651), .ZN(n546) );
  NAND2_X1 U654 ( .A1(n547), .A2(n682), .ZN(n548) );
  XNOR2_X1 U655 ( .A(n549), .B(n548), .ZN(n738) );
  XNOR2_X1 U656 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X2 U657 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U658 ( .A(n554), .B(KEYINPUT48), .ZN(n562) );
  NOR2_X1 U659 ( .A1(n579), .A2(n555), .ZN(n556) );
  XNOR2_X1 U660 ( .A(n556), .B(KEYINPUT43), .ZN(n557) );
  NOR2_X1 U661 ( .A1(n558), .A2(n557), .ZN(n641) );
  NAND2_X1 U662 ( .A1(n636), .A2(n559), .ZN(n640) );
  AND2_X2 U663 ( .A1(n562), .A2(n561), .ZN(n726) );
  INV_X1 U664 ( .A(n726), .ZN(n642) );
  INV_X1 U665 ( .A(n563), .ZN(n564) );
  NOR2_X1 U666 ( .A1(G898), .A2(n728), .ZN(n717) );
  NAND2_X1 U667 ( .A1(n564), .A2(n717), .ZN(n565) );
  XOR2_X1 U668 ( .A(KEYINPUT88), .B(n565), .Z(n566) );
  OR2_X1 U669 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U670 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U671 ( .A(n650), .ZN(n574) );
  AND2_X1 U672 ( .A1(n574), .A2(n662), .ZN(n575) );
  XNOR2_X1 U673 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n577) );
  NOR2_X1 U674 ( .A1(n591), .A2(n579), .ZN(n582) );
  NOR2_X1 U675 ( .A1(n376), .A2(n580), .ZN(n581) );
  NAND2_X1 U676 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U677 ( .A(n583), .B(KEYINPUT107), .ZN(n734) );
  INV_X1 U678 ( .A(KEYINPUT64), .ZN(n588) );
  XNOR2_X1 U679 ( .A(n584), .B(KEYINPUT105), .ZN(n585) );
  NOR2_X1 U680 ( .A1(n590), .A2(n585), .ZN(n586) );
  XNOR2_X1 U681 ( .A(n586), .B(KEYINPUT73), .ZN(n587) );
  NAND2_X1 U682 ( .A1(n589), .A2(n733), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n607), .A2(KEYINPUT44), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n658), .A2(n376), .ZN(n594) );
  NOR2_X1 U685 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U686 ( .A(n592), .B(KEYINPUT81), .ZN(n593) );
  NOR2_X1 U687 ( .A1(n594), .A2(n593), .ZN(n619) );
  NAND2_X1 U688 ( .A1(n370), .A2(n595), .ZN(n669) );
  NOR2_X1 U689 ( .A1(n669), .A2(n596), .ZN(n598) );
  XOR2_X1 U690 ( .A(KEYINPUT94), .B(KEYINPUT31), .Z(n597) );
  XNOR2_X1 U691 ( .A(n598), .B(n597), .ZN(n637) );
  NOR2_X1 U692 ( .A1(n637), .A2(n624), .ZN(n601) );
  XNOR2_X1 U693 ( .A(n603), .B(n602), .ZN(n604) );
  NOR2_X1 U694 ( .A1(n619), .A2(n604), .ZN(n605) );
  INV_X1 U695 ( .A(KEYINPUT2), .ZN(n610) );
  NOR2_X2 U696 ( .A1(n613), .A2(n710), .ZN(n645) );
  NAND2_X1 U697 ( .A1(n705), .A2(G472), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U699 ( .A(KEYINPUT63), .B(KEYINPUT83), .ZN(n618) );
  XOR2_X1 U700 ( .A(G101), .B(n619), .Z(G3) );
  NAND2_X1 U701 ( .A1(n624), .A2(n633), .ZN(n620) );
  XNOR2_X1 U702 ( .A(n620), .B(G104), .ZN(G6) );
  XOR2_X1 U703 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n622) );
  XNOR2_X1 U704 ( .A(G107), .B(KEYINPUT26), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n622), .B(n621), .ZN(n623) );
  XOR2_X1 U706 ( .A(KEYINPUT113), .B(n623), .Z(n626) );
  NAND2_X1 U707 ( .A1(n624), .A2(n636), .ZN(n625) );
  XNOR2_X1 U708 ( .A(n626), .B(n625), .ZN(G9) );
  XOR2_X1 U709 ( .A(G128), .B(KEYINPUT29), .Z(n629) );
  INV_X1 U710 ( .A(n627), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n631), .A2(n636), .ZN(n628) );
  XNOR2_X1 U712 ( .A(n629), .B(n628), .ZN(G30) );
  XOR2_X1 U713 ( .A(G143), .B(n630), .Z(G45) );
  NAND2_X1 U714 ( .A1(n631), .A2(n633), .ZN(n632) );
  XNOR2_X1 U715 ( .A(n632), .B(G146), .ZN(G48) );
  XOR2_X1 U716 ( .A(G113), .B(KEYINPUT115), .Z(n635) );
  NAND2_X1 U717 ( .A1(n633), .A2(n637), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n635), .B(n634), .ZN(G15) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n638), .B(KEYINPUT116), .ZN(n639) );
  XNOR2_X1 U721 ( .A(G116), .B(n639), .ZN(G18) );
  XNOR2_X1 U722 ( .A(G134), .B(n640), .ZN(G36) );
  XOR2_X1 U723 ( .A(G140), .B(n641), .Z(G42) );
  XNOR2_X1 U724 ( .A(n644), .B(KEYINPUT74), .ZN(n646) );
  NOR2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  NOR2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT119), .B(n657), .ZN(n675) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U732 ( .A(KEYINPUT50), .B(n660), .Z(n661) );
  XNOR2_X1 U733 ( .A(n661), .B(KEYINPUT117), .ZN(n668) );
  NOR2_X1 U734 ( .A1(n376), .A2(n662), .ZN(n664) );
  XOR2_X1 U735 ( .A(KEYINPUT49), .B(n664), .Z(n665) );
  NOR2_X1 U736 ( .A1(n370), .A2(n665), .ZN(n667) );
  NAND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U739 ( .A(KEYINPUT51), .B(n671), .Z(n672) );
  NAND2_X1 U740 ( .A1(n682), .A2(n672), .ZN(n673) );
  XNOR2_X1 U741 ( .A(KEYINPUT118), .B(n673), .ZN(n674) );
  NAND2_X1 U742 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U743 ( .A(n676), .B(KEYINPUT120), .ZN(n677) );
  XOR2_X1 U744 ( .A(KEYINPUT52), .B(n677), .Z(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U746 ( .A(n680), .B(KEYINPUT121), .ZN(n684) );
  NAND2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U749 ( .A1(n705), .A2(G210), .ZN(n690) );
  XNOR2_X1 U750 ( .A(n688), .B(n433), .ZN(n689) );
  XNOR2_X1 U751 ( .A(n690), .B(n689), .ZN(n691) );
  XOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n693) );
  NAND2_X1 U753 ( .A1(n705), .A2(G469), .ZN(n692) );
  NOR2_X1 U754 ( .A1(n709), .A2(n695), .ZN(G54) );
  NAND2_X1 U755 ( .A1(n705), .A2(G475), .ZN(n697) );
  XNOR2_X1 U756 ( .A(n700), .B(KEYINPUT60), .ZN(G60) );
  XOR2_X1 U757 ( .A(n701), .B(KEYINPUT123), .Z(n703) );
  NAND2_X1 U758 ( .A1(n705), .A2(G478), .ZN(n702) );
  XNOR2_X1 U759 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n709), .A2(n704), .ZN(G63) );
  XNOR2_X1 U761 ( .A(n706), .B(n707), .ZN(n708) );
  OR2_X1 U762 ( .A1(G953), .A2(n710), .ZN(n714) );
  NAND2_X1 U763 ( .A1(G953), .A2(G224), .ZN(n711) );
  XNOR2_X1 U764 ( .A(KEYINPUT61), .B(n711), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n712), .A2(G898), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n714), .A2(n713), .ZN(n719) );
  XOR2_X1 U767 ( .A(n715), .B(KEYINPUT125), .Z(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(G69) );
  XOR2_X1 U770 ( .A(n720), .B(KEYINPUT90), .Z(n721) );
  XOR2_X1 U771 ( .A(n722), .B(n721), .Z(n727) );
  XOR2_X1 U772 ( .A(n727), .B(KEYINPUT126), .Z(n723) );
  XNOR2_X1 U773 ( .A(G227), .B(n723), .ZN(n724) );
  NAND2_X1 U774 ( .A1(G900), .A2(n724), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(G953), .ZN(n731) );
  XNOR2_X1 U776 ( .A(n727), .B(n372), .ZN(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U779 ( .A(n732), .B(G122), .Z(G24) );
  XNOR2_X1 U780 ( .A(G119), .B(n733), .ZN(G21) );
  XOR2_X1 U781 ( .A(n734), .B(G110), .Z(G12) );
  XOR2_X1 U782 ( .A(n735), .B(G125), .Z(n736) );
  XNOR2_X1 U783 ( .A(KEYINPUT37), .B(n736), .ZN(G27) );
  XNOR2_X1 U784 ( .A(n737), .B(G131), .ZN(G33) );
  XOR2_X1 U785 ( .A(G137), .B(n738), .Z(n739) );
  XNOR2_X1 U786 ( .A(KEYINPUT127), .B(n739), .ZN(G39) );
endmodule

