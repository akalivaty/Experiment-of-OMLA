

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XOR2_X2 U323 ( .A(n440), .B(n439), .Z(n574) );
  NOR2_X1 U324 ( .A1(n565), .A2(n543), .ZN(n545) );
  XOR2_X1 U325 ( .A(n435), .B(KEYINPUT88), .Z(n291) );
  XOR2_X1 U326 ( .A(G64GAT), .B(KEYINPUT85), .Z(n292) );
  XOR2_X1 U327 ( .A(KEYINPUT74), .B(KEYINPUT13), .Z(n293) );
  NOR2_X1 U328 ( .A1(n552), .A2(n566), .ZN(n496) );
  NOR2_X1 U329 ( .A1(n498), .A2(n497), .ZN(n500) );
  NOR2_X1 U330 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U331 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U332 ( .A(n349), .B(n348), .ZN(n353) );
  XNOR2_X1 U333 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n447) );
  XOR2_X1 U334 ( .A(KEYINPUT97), .B(KEYINPUT6), .Z(n295) );
  XNOR2_X1 U335 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n313) );
  XOR2_X1 U337 ( .A(G85GAT), .B(G162GAT), .Z(n297) );
  XNOR2_X1 U338 ( .A(G29GAT), .B(G141GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U340 ( .A(KEYINPUT5), .B(G57GAT), .Z(n299) );
  XNOR2_X1 U341 ( .A(G1GAT), .B(G155GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U343 ( .A(n301), .B(n300), .Z(n311) );
  XNOR2_X1 U344 ( .A(G127GAT), .B(G134GAT), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n302), .B(KEYINPUT0), .ZN(n303) );
  XOR2_X1 U346 ( .A(n303), .B(KEYINPUT90), .Z(n305) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G120GAT), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n305), .B(n304), .ZN(n386) );
  XNOR2_X1 U349 ( .A(G148GAT), .B(KEYINPUT3), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n306), .B(KEYINPUT2), .ZN(n365) );
  XOR2_X1 U351 ( .A(n365), .B(KEYINPUT98), .Z(n308) );
  NAND2_X1 U352 ( .A1(G225GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U354 ( .A(n386), .B(n309), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U356 ( .A(n313), .B(n312), .Z(n482) );
  XOR2_X1 U357 ( .A(KEYINPUT29), .B(KEYINPUT71), .Z(n315) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(G8GAT), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U360 ( .A(n316), .B(G197GAT), .Z(n318) );
  XOR2_X1 U361 ( .A(G15GAT), .B(G1GAT), .Z(n430) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(n430), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n333) );
  XOR2_X1 U364 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n320) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U367 ( .A(G141GAT), .B(G22GAT), .Z(n359) );
  XOR2_X1 U368 ( .A(n321), .B(n359), .Z(n331) );
  XOR2_X1 U369 ( .A(G43GAT), .B(G29GAT), .Z(n323) );
  XNOR2_X1 U370 ( .A(KEYINPUT8), .B(G50GAT), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U372 ( .A(n324), .B(KEYINPUT7), .Z(n326) );
  XNOR2_X1 U373 ( .A(G36GAT), .B(KEYINPUT70), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n422) );
  XOR2_X1 U375 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n328) );
  XNOR2_X1 U376 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U378 ( .A(n422), .B(n329), .ZN(n330) );
  XNOR2_X1 U379 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U380 ( .A(n333), .B(n332), .ZN(n566) );
  XNOR2_X1 U381 ( .A(KEYINPUT73), .B(n566), .ZN(n549) );
  XOR2_X1 U382 ( .A(KEYINPUT79), .B(G64GAT), .Z(n335) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(G78GAT), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U385 ( .A(G148GAT), .B(G92GAT), .Z(n336) );
  XNOR2_X1 U386 ( .A(n337), .B(n336), .ZN(n345) );
  XNOR2_X1 U387 ( .A(KEYINPUT32), .B(KEYINPUT78), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n338), .B(KEYINPUT31), .ZN(n339) );
  XOR2_X1 U389 ( .A(n339), .B(KEYINPUT80), .Z(n343) );
  XNOR2_X1 U390 ( .A(G71GAT), .B(G57GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n293), .B(n340), .ZN(n427) );
  XNOR2_X1 U392 ( .A(G176GAT), .B(G204GAT), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n341), .B(KEYINPUT77), .ZN(n389) );
  XNOR2_X1 U394 ( .A(n427), .B(n389), .ZN(n342) );
  XNOR2_X1 U395 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n349) );
  NAND2_X1 U397 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  INV_X1 U398 ( .A(KEYINPUT75), .ZN(n346) );
  XOR2_X1 U399 ( .A(KEYINPUT76), .B(G85GAT), .Z(n351) );
  XNOR2_X1 U400 ( .A(G99GAT), .B(G106GAT), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n410) );
  XNOR2_X1 U402 ( .A(n410), .B(KEYINPUT33), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n570) );
  NAND2_X1 U404 ( .A1(n549), .A2(n570), .ZN(n459) );
  XOR2_X1 U405 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n355) );
  XNOR2_X1 U406 ( .A(KEYINPUT95), .B(KEYINPUT93), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n371) );
  XOR2_X1 U408 ( .A(G155GAT), .B(G78GAT), .Z(n429) );
  XOR2_X1 U409 ( .A(G106GAT), .B(n429), .Z(n357) );
  XOR2_X1 U410 ( .A(G218GAT), .B(G162GAT), .Z(n411) );
  XNOR2_X1 U411 ( .A(G50GAT), .B(n411), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n369) );
  XOR2_X1 U414 ( .A(KEYINPUT24), .B(G204GAT), .Z(n361) );
  NAND2_X1 U415 ( .A1(G228GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U417 ( .A(n362), .B(KEYINPUT22), .Z(n367) );
  XOR2_X1 U418 ( .A(G211GAT), .B(KEYINPUT21), .Z(n364) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(KEYINPUT94), .ZN(n363) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n390) );
  XNOR2_X1 U421 ( .A(n365), .B(n390), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n543) );
  XOR2_X1 U425 ( .A(G99GAT), .B(G190GAT), .Z(n373) );
  NAND2_X1 U426 ( .A1(G227GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n376) );
  XOR2_X1 U428 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n375) );
  XNOR2_X1 U429 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n391) );
  XOR2_X1 U431 ( .A(n376), .B(n391), .Z(n384) );
  XOR2_X1 U432 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n378) );
  XNOR2_X1 U433 ( .A(G43GAT), .B(KEYINPUT91), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U435 ( .A(G71GAT), .B(G176GAT), .Z(n380) );
  XNOR2_X1 U436 ( .A(G15GAT), .B(G183GAT), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(n386), .B(n385), .Z(n507) );
  NAND2_X1 U441 ( .A1(n543), .A2(n507), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n387), .B(KEYINPUT26), .ZN(n564) );
  XNOR2_X1 U443 ( .A(G190GAT), .B(G92GAT), .ZN(n388) );
  XNOR2_X1 U444 ( .A(n388), .B(KEYINPUT83), .ZN(n414) );
  XOR2_X1 U445 ( .A(n389), .B(n414), .Z(n393) );
  XNOR2_X1 U446 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n399) );
  XNOR2_X1 U448 ( .A(G8GAT), .B(G183GAT), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n292), .B(n394), .ZN(n435) );
  XOR2_X1 U450 ( .A(G218GAT), .B(G36GAT), .Z(n396) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U453 ( .A(n435), .B(n397), .Z(n398) );
  XOR2_X1 U454 ( .A(n399), .B(n398), .Z(n485) );
  XOR2_X1 U455 ( .A(KEYINPUT27), .B(n485), .Z(n405) );
  NOR2_X1 U456 ( .A1(n564), .A2(n405), .ZN(n523) );
  INV_X1 U457 ( .A(n485), .ZN(n538) );
  NOR2_X1 U458 ( .A1(n507), .A2(n538), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n543), .A2(n400), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n401), .B(KEYINPUT25), .ZN(n402) );
  XNOR2_X1 U461 ( .A(KEYINPUT99), .B(n402), .ZN(n403) );
  NOR2_X1 U462 ( .A1(n523), .A2(n403), .ZN(n404) );
  NOR2_X1 U463 ( .A1(n482), .A2(n404), .ZN(n409) );
  XOR2_X1 U464 ( .A(KEYINPUT28), .B(n543), .Z(n466) );
  INV_X1 U465 ( .A(n466), .ZN(n490) );
  INV_X1 U466 ( .A(n482), .ZN(n540) );
  NOR2_X1 U467 ( .A1(n490), .A2(n540), .ZN(n407) );
  INV_X1 U468 ( .A(n405), .ZN(n406) );
  NAND2_X1 U469 ( .A1(n407), .A2(n406), .ZN(n509) );
  INV_X1 U470 ( .A(n507), .ZN(n546) );
  NOR2_X1 U471 ( .A1(n509), .A2(n546), .ZN(n408) );
  NOR2_X1 U472 ( .A1(n409), .A2(n408), .ZN(n455) );
  XOR2_X1 U473 ( .A(KEYINPUT16), .B(KEYINPUT89), .Z(n443) );
  XOR2_X1 U474 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n413) );
  XNOR2_X1 U475 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n418) );
  XOR2_X1 U477 ( .A(n414), .B(KEYINPUT65), .Z(n416) );
  NAND2_X1 U478 ( .A1(G232GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U480 ( .A(n418), .B(n417), .Z(n424) );
  XOR2_X1 U481 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n420) );
  XNOR2_X1 U482 ( .A(G134GAT), .B(KEYINPUT82), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U484 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n534) );
  XNOR2_X1 U486 ( .A(n534), .B(KEYINPUT84), .ZN(n559) );
  XOR2_X1 U487 ( .A(KEYINPUT87), .B(KEYINPUT14), .Z(n426) );
  XNOR2_X1 U488 ( .A(KEYINPUT86), .B(KEYINPUT12), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n440) );
  XOR2_X1 U493 ( .A(KEYINPUT15), .B(G211GAT), .Z(n434) );
  XNOR2_X1 U494 ( .A(G22GAT), .B(G127GAT), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n438) );
  NAND2_X1 U496 ( .A1(G231GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n291), .B(n436), .ZN(n437) );
  XOR2_X1 U498 ( .A(n438), .B(n437), .Z(n439) );
  INV_X1 U499 ( .A(n574), .ZN(n441) );
  NAND2_X1 U500 ( .A1(n559), .A2(n441), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  OR2_X1 U502 ( .A1(n455), .A2(n444), .ZN(n470) );
  NOR2_X1 U503 ( .A1(n459), .A2(n470), .ZN(n445) );
  XNOR2_X1 U504 ( .A(KEYINPUT100), .B(n445), .ZN(n452) );
  NAND2_X1 U505 ( .A1(n482), .A2(n452), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(G1324GAT) );
  NAND2_X1 U507 ( .A1(n485), .A2(n452), .ZN(n448) );
  XNOR2_X1 U508 ( .A(G8GAT), .B(n448), .ZN(G1325GAT) );
  XOR2_X1 U509 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n450) );
  NAND2_X1 U510 ( .A1(n452), .A2(n546), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U512 ( .A(G15GAT), .B(n451), .Z(G1326GAT) );
  NAND2_X1 U513 ( .A1(n452), .A2(n490), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(KEYINPUT102), .ZN(n454) );
  XNOR2_X1 U515 ( .A(G22GAT), .B(n454), .ZN(G1327GAT) );
  XNOR2_X1 U516 ( .A(KEYINPUT36), .B(n559), .ZN(n580) );
  NOR2_X1 U517 ( .A1(n580), .A2(n455), .ZN(n456) );
  NAND2_X1 U518 ( .A1(n574), .A2(n456), .ZN(n457) );
  XNOR2_X1 U519 ( .A(KEYINPUT37), .B(n457), .ZN(n458) );
  XNOR2_X1 U520 ( .A(KEYINPUT103), .B(n458), .ZN(n480) );
  NOR2_X1 U521 ( .A1(n480), .A2(n459), .ZN(n460) );
  XOR2_X1 U522 ( .A(KEYINPUT38), .B(n460), .Z(n467) );
  NOR2_X1 U523 ( .A1(n467), .A2(n540), .ZN(n462) );
  XNOR2_X1 U524 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n461) );
  XNOR2_X1 U525 ( .A(n462), .B(n461), .ZN(G1328GAT) );
  NOR2_X1 U526 ( .A1(n467), .A2(n538), .ZN(n463) );
  XOR2_X1 U527 ( .A(G36GAT), .B(n463), .Z(G1329GAT) );
  NOR2_X1 U528 ( .A1(n507), .A2(n467), .ZN(n464) );
  XOR2_X1 U529 ( .A(KEYINPUT40), .B(n464), .Z(n465) );
  XNOR2_X1 U530 ( .A(G43GAT), .B(n465), .ZN(G1330GAT) );
  NOR2_X1 U531 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U532 ( .A(G50GAT), .B(n468), .Z(G1331GAT) );
  XNOR2_X1 U533 ( .A(KEYINPUT41), .B(n570), .ZN(n511) );
  NAND2_X1 U534 ( .A1(n511), .A2(n566), .ZN(n469) );
  XNOR2_X1 U535 ( .A(n469), .B(KEYINPUT104), .ZN(n481) );
  NOR2_X1 U536 ( .A1(n481), .A2(n470), .ZN(n471) );
  XOR2_X1 U537 ( .A(KEYINPUT105), .B(n471), .Z(n477) );
  NAND2_X1 U538 ( .A1(n477), .A2(n482), .ZN(n472) );
  XNOR2_X1 U539 ( .A(n472), .B(KEYINPUT42), .ZN(n473) );
  XNOR2_X1 U540 ( .A(G57GAT), .B(n473), .ZN(G1332GAT) );
  NAND2_X1 U541 ( .A1(n477), .A2(n485), .ZN(n474) );
  XNOR2_X1 U542 ( .A(n474), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U543 ( .A1(n546), .A2(n477), .ZN(n475) );
  XNOR2_X1 U544 ( .A(n475), .B(KEYINPUT106), .ZN(n476) );
  XNOR2_X1 U545 ( .A(G71GAT), .B(n476), .ZN(G1334GAT) );
  XOR2_X1 U546 ( .A(G78GAT), .B(KEYINPUT43), .Z(n479) );
  NAND2_X1 U547 ( .A1(n477), .A2(n490), .ZN(n478) );
  XNOR2_X1 U548 ( .A(n479), .B(n478), .ZN(G1335GAT) );
  XOR2_X1 U549 ( .A(G85GAT), .B(KEYINPUT107), .Z(n484) );
  NOR2_X1 U550 ( .A1(n481), .A2(n480), .ZN(n491) );
  NAND2_X1 U551 ( .A1(n491), .A2(n482), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n484), .B(n483), .ZN(G1336GAT) );
  NAND2_X1 U553 ( .A1(n491), .A2(n485), .ZN(n486) );
  XNOR2_X1 U554 ( .A(n486), .B(KEYINPUT108), .ZN(n487) );
  XNOR2_X1 U555 ( .A(G92GAT), .B(n487), .ZN(G1337GAT) );
  XOR2_X1 U556 ( .A(G99GAT), .B(KEYINPUT109), .Z(n489) );
  NAND2_X1 U557 ( .A1(n491), .A2(n546), .ZN(n488) );
  XNOR2_X1 U558 ( .A(n489), .B(n488), .ZN(G1338GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n493) );
  NAND2_X1 U560 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U561 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U562 ( .A(G106GAT), .B(n494), .Z(G1339GAT) );
  INV_X1 U563 ( .A(n511), .ZN(n552) );
  XNOR2_X1 U564 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n495) );
  XNOR2_X1 U565 ( .A(n496), .B(n495), .ZN(n498) );
  XOR2_X1 U566 ( .A(KEYINPUT111), .B(n574), .Z(n557) );
  NAND2_X1 U567 ( .A1(n557), .A2(n534), .ZN(n497) );
  XNOR2_X1 U568 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n499) );
  XNOR2_X1 U569 ( .A(n500), .B(n499), .ZN(n505) );
  NOR2_X1 U570 ( .A1(n574), .A2(n580), .ZN(n501) );
  XNOR2_X1 U571 ( .A(KEYINPUT45), .B(n501), .ZN(n502) );
  NAND2_X1 U572 ( .A1(n570), .A2(n502), .ZN(n503) );
  NOR2_X1 U573 ( .A1(n549), .A2(n503), .ZN(n504) );
  NOR2_X1 U574 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U575 ( .A(KEYINPUT48), .B(n506), .ZN(n537) );
  OR2_X1 U576 ( .A1(n537), .A2(n507), .ZN(n508) );
  NOR2_X1 U577 ( .A1(n509), .A2(n508), .ZN(n514) );
  NAND2_X1 U578 ( .A1(n549), .A2(n514), .ZN(n510) );
  XNOR2_X1 U579 ( .A(G113GAT), .B(n510), .ZN(G1340GAT) );
  XOR2_X1 U580 ( .A(G120GAT), .B(KEYINPUT49), .Z(n513) );
  NAND2_X1 U581 ( .A1(n514), .A2(n511), .ZN(n512) );
  XNOR2_X1 U582 ( .A(n513), .B(n512), .ZN(G1341GAT) );
  INV_X1 U583 ( .A(n514), .ZN(n518) );
  NOR2_X1 U584 ( .A1(n557), .A2(n518), .ZN(n516) );
  XNOR2_X1 U585 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n515) );
  XNOR2_X1 U586 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U587 ( .A(G127GAT), .B(n517), .Z(G1342GAT) );
  NOR2_X1 U588 ( .A1(n559), .A2(n518), .ZN(n520) );
  XNOR2_X1 U589 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n519) );
  XNOR2_X1 U590 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U591 ( .A(G134GAT), .B(n521), .Z(G1343GAT) );
  NOR2_X1 U592 ( .A1(n540), .A2(n537), .ZN(n522) );
  NAND2_X1 U593 ( .A1(n523), .A2(n522), .ZN(n533) );
  NOR2_X1 U594 ( .A1(n566), .A2(n533), .ZN(n524) );
  XOR2_X1 U595 ( .A(KEYINPUT116), .B(n524), .Z(n525) );
  XNOR2_X1 U596 ( .A(G141GAT), .B(n525), .ZN(G1344GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n527) );
  XNOR2_X1 U598 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n526) );
  XNOR2_X1 U599 ( .A(n527), .B(n526), .ZN(n531) );
  NOR2_X1 U600 ( .A1(n552), .A2(n533), .ZN(n529) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n528) );
  XNOR2_X1 U602 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U603 ( .A(n531), .B(n530), .Z(G1345GAT) );
  NOR2_X1 U604 ( .A1(n574), .A2(n533), .ZN(n532) );
  XOR2_X1 U605 ( .A(G155GAT), .B(n532), .Z(G1346GAT) );
  NOR2_X1 U606 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U607 ( .A(KEYINPUT120), .B(n535), .Z(n536) );
  XNOR2_X1 U608 ( .A(G162GAT), .B(n536), .ZN(G1347GAT) );
  XNOR2_X1 U609 ( .A(n539), .B(KEYINPUT54), .ZN(n541) );
  NAND2_X1 U610 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n542), .B(KEYINPUT64), .ZN(n565) );
  XNOR2_X1 U612 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT122), .ZN(n560) );
  INV_X1 U616 ( .A(n560), .ZN(n550) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G169GAT), .ZN(G1348GAT) );
  OR2_X1 U619 ( .A1(n560), .A2(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT56), .Z(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n560), .ZN(n558) );
  XOR2_X1 U625 ( .A(G183GAT), .B(n558), .Z(G1350GAT) );
  INV_X1 U626 ( .A(KEYINPUT58), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(n563), .ZN(G1351GAT) );
  OR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n579) );
  NOR2_X1 U631 ( .A1(n566), .A2(n579), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n579), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n579), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n582) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(n582), .B(n581), .Z(G1355GAT) );
endmodule

