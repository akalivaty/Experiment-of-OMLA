//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n437, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT70), .B(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n466), .A2(KEYINPUT71), .A3(G137), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n472), .A2(G137), .A3(new_n467), .A4(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT71), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n468), .A2(new_n477), .B1(G101), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT69), .B1(new_n464), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n474), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(G113), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2105), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n479), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT72), .ZN(G160));
  NAND2_X1  g066(.A1(new_n472), .A2(new_n474), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(new_n467), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT73), .Z(new_n495));
  NOR2_X1   g070(.A1(new_n492), .A2(G2105), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G136), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n467), .A2(G112), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n495), .A2(new_n500), .ZN(G162));
  AND2_X1   g076(.A1(KEYINPUT74), .A2(G114), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT74), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(G2105), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n504), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n472), .A2(G126), .A3(G2105), .A4(new_n474), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n505), .B2(new_n506), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND3_X1   g085(.A1(new_n474), .A2(new_n483), .A3(new_n484), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n484), .B1(new_n474), .B2(new_n483), .ZN(new_n512));
  OAI211_X1 g087(.A(G138), .B(new_n467), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT4), .A2(G138), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n496), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n510), .A2(new_n518), .ZN(G164));
  AOI21_X1  g094(.A(KEYINPUT78), .B1(KEYINPUT77), .B2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT78), .A2(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT6), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(G651), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT76), .B1(new_n528), .B2(KEYINPUT6), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(new_n531), .A3(G651), .ZN(new_n535));
  AOI211_X1 g110(.A(new_n530), .B(new_n532), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G50), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n526), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n529), .A2(new_n541), .ZN(G166));
  INV_X1    g117(.A(KEYINPUT79), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n536), .B(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G51), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n526), .A2(new_n538), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G89), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT7), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g126(.A1(new_n545), .A2(new_n547), .A3(new_n551), .ZN(G168));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n524), .A2(new_n525), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n536), .B(KEYINPUT79), .ZN(new_n559));
  INV_X1    g134(.A(G52), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n557), .B1(new_n558), .B2(new_n539), .C1(new_n559), .C2(new_n560), .ZN(G301));
  INV_X1    g136(.A(G301), .ZN(G171));
  NAND2_X1  g137(.A1(new_n544), .A2(G43), .ZN(new_n563));
  NAND2_X1  g138(.A1(G68), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G56), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n554), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n546), .A2(G81), .B1(new_n566), .B2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n554), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n546), .A2(G91), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n538), .A2(KEYINPUT80), .A3(G53), .A4(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G299));
  NAND3_X1  g157(.A1(new_n545), .A2(new_n547), .A3(new_n551), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  NAND2_X1  g159(.A1(new_n546), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n536), .A2(G49), .ZN(new_n587));
  AND3_X1   g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G288));
  NAND4_X1  g164(.A1(new_n526), .A2(KEYINPUT81), .A3(G86), .A4(new_n538), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n538), .A2(new_n524), .A3(G86), .A4(new_n525), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n530), .B1(KEYINPUT78), .B2(KEYINPUT5), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n525), .B(G61), .C1(new_n595), .C2(new_n520), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n536), .B2(G48), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n594), .A2(new_n599), .ZN(G305));
  AND2_X1   g175(.A1(new_n544), .A2(G47), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n602), .A2(new_n528), .B1(new_n603), .B2(new_n539), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n526), .A2(G92), .A3(new_n538), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT82), .B(G66), .Z(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n554), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n544), .A2(G54), .B1(G651), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G868), .ZN(G284));
  OAI21_X1  g190(.A(new_n607), .B1(new_n614), .B2(G868), .ZN(G321));
  XOR2_X1   g191(.A(G299), .B(KEYINPUT83), .Z(new_n617));
  MUX2_X1   g192(.A(new_n617), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g193(.A(new_n617), .B(G286), .S(G868), .Z(G280));
  XOR2_X1   g194(.A(KEYINPUT84), .B(G559), .Z(new_n620));
  OAI21_X1  g195(.A(new_n614), .B1(G860), .B2(new_n620), .ZN(G148));
  NAND2_X1  g196(.A1(new_n614), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g200(.A1(new_n511), .A2(new_n512), .ZN(new_n626));
  OR3_X1    g201(.A1(new_n626), .A2(G2105), .A3(new_n465), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2100), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n496), .A2(G135), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT85), .ZN(new_n633));
  OR2_X1    g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n634), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n493), .A2(G123), .ZN(new_n636));
  AND3_X1   g211(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n631), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT86), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2072), .B(G2078), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT87), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2084), .B(G2090), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n662), .B1(new_n659), .B2(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n660), .B2(new_n661), .ZN(new_n665));
  INV_X1    g240(.A(new_n661), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n666), .A2(new_n662), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT18), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT89), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT90), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n679), .A2(new_n680), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n676), .A2(new_n677), .A3(new_n681), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n678), .A2(new_n687), .ZN(new_n690));
  NAND4_X1  g265(.A1(new_n685), .A2(new_n686), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  MUX2_X1   g274(.A(G6), .B(G305), .S(G16), .Z(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT32), .B(G1981), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n703), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(G23), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n588), .B2(new_n703), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AND3_X1   g286(.A1(new_n702), .A2(new_n707), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT93), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n496), .A2(G131), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n493), .A2(G119), .ZN(new_n720));
  OR2_X1    g295(.A1(G95), .A2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G2104), .C1(G107), .C2(new_n467), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(new_n717), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n605), .A2(G16), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G16), .B2(G24), .ZN(new_n730));
  INV_X1    g305(.A(G1986), .ZN(new_n731));
  AOI21_X1  g306(.A(KEYINPUT94), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n731), .B2(new_n730), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n728), .B(new_n733), .C1(new_n712), .C2(new_n713), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n716), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n716), .A2(KEYINPUT36), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n496), .A2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n493), .A2(G128), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n467), .A2(G116), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G29), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n717), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT97), .B(G2067), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n703), .A2(G19), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n569), .B2(new_n703), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1341), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n703), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n703), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n750), .B(new_n753), .C1(G1966), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n703), .A2(G20), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT23), .Z(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G299), .B2(G16), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1956), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n496), .A2(G141), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n493), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT26), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n478), .A2(G105), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n761), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G32), .B(new_n768), .S(G29), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT27), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1996), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n703), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G171), .B2(new_n703), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1961), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT31), .B(G11), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT30), .B(G28), .Z(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n637), .B2(G29), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n755), .B2(G1966), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n756), .A2(new_n760), .A3(new_n771), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G29), .A2(G35), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G162), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(G2090), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(G2090), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n717), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n717), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(G2078), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n703), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n614), .B2(new_n703), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT95), .B(G1348), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n786), .A2(new_n787), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  AND2_X1   g370(.A1(KEYINPUT24), .A2(G34), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n717), .B1(KEYINPUT24), .B2(G34), .ZN(new_n797));
  OAI22_X1  g372(.A1(G160), .A2(new_n717), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2084), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n717), .A2(G33), .ZN(new_n800));
  NAND2_X1  g375(.A1(G115), .A2(G2104), .ZN(new_n801));
  INV_X1    g376(.A(G127), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n626), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n467), .B1(new_n803), .B2(KEYINPUT99), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(KEYINPUT99), .B2(new_n803), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT25), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(KEYINPUT25), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n808), .A2(new_n809), .B1(G139), .B2(new_n496), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n800), .B1(new_n813), .B2(new_n717), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G2072), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n781), .A2(new_n795), .A3(new_n799), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n737), .A2(new_n738), .A3(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NAND2_X1  g393(.A1(new_n614), .A2(G559), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n554), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G651), .ZN(new_n825));
  INV_X1    g400(.A(G93), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n539), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G55), .B2(new_n544), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n569), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G55), .ZN(new_n830));
  OAI221_X1 g405(.A(new_n825), .B1(new_n826), .B2(new_n539), .C1(new_n559), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(new_n568), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n821), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n831), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT103), .Z(G145));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n743), .B(new_n768), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n813), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n811), .B(KEYINPUT100), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n505), .A2(new_n506), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n515), .A2(new_n849), .A3(new_n517), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n845), .A2(new_n847), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n628), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n496), .A2(G142), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n493), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n467), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n854), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n854), .A2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n723), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n628), .B(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n724), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n851), .A2(new_n853), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n853), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n852), .B1(new_n845), .B2(new_n847), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n851), .A2(new_n853), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(new_n865), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n868), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G160), .B(new_n637), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n842), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(KEYINPUT105), .B1(new_n869), .B2(new_n870), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n851), .A2(new_n881), .A3(new_n853), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n882), .A3(new_n866), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n874), .B1(new_n873), .B2(new_n865), .ZN(new_n884));
  AOI211_X1 g459(.A(KEYINPUT104), .B(new_n866), .C1(new_n851), .C2(new_n853), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n883), .B(new_n878), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n879), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n867), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(new_n878), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT40), .B1(new_n892), .B2(new_n886), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n889), .A2(new_n893), .ZN(G395));
  XNOR2_X1  g469(.A(new_n605), .B(G305), .ZN(new_n895));
  XNOR2_X1  g470(.A(G303), .B(new_n588), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT42), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n614), .A2(G299), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n609), .A2(new_n613), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n581), .A3(new_n579), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT41), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(KEYINPUT41), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n833), .B(new_n622), .ZN(new_n907));
  MUX2_X1   g482(.A(new_n906), .B(new_n902), .S(new_n907), .Z(new_n908));
  XNOR2_X1  g483(.A(new_n898), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(G868), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(G868), .B2(new_n828), .ZN(G295));
  OAI21_X1  g486(.A(new_n910), .B1(G868), .B2(new_n828), .ZN(G331));
  NAND2_X1  g487(.A1(G171), .A2(G168), .ZN(new_n913));
  NAND2_X1  g488(.A1(G301), .A2(G286), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n833), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n913), .A2(new_n829), .A3(new_n832), .A4(new_n914), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n906), .A2(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n917), .A2(new_n902), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(KEYINPUT106), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT106), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(new_n833), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n924), .A3(new_n897), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n842), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n897), .B1(new_n919), .B2(new_n924), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n921), .A2(new_n923), .A3(new_n917), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n930), .A2(new_n906), .B1(new_n916), .B2(new_n920), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n842), .B(new_n925), .C1(new_n931), .C2(new_n897), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n928), .B2(new_n933), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n926), .C2(new_n927), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n932), .B2(KEYINPUT43), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n931), .A2(new_n897), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n925), .A2(new_n842), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n942), .A3(KEYINPUT108), .A4(new_n933), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n937), .A2(new_n938), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n935), .B1(new_n944), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g520(.A(KEYINPUT51), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n468), .A2(new_n477), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n478), .A2(G101), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n489), .A3(G40), .A4(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G40), .ZN(new_n953));
  OAI21_X1  g528(.A(G125), .B1(new_n511), .B2(new_n512), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n487), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n955), .B2(G2105), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(KEYINPUT109), .A3(new_n479), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n850), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n952), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n514), .A2(new_n513), .B1(new_n496), .B2(new_n516), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n509), .B2(new_n508), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n958), .B1(new_n963), .B2(new_n959), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n961), .A2(new_n964), .A3(G2084), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n952), .A2(new_n957), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT45), .B1(new_n850), .B2(new_n959), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n968), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n970), .A2(KEYINPUT115), .A3(new_n952), .A4(new_n957), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(G1966), .ZN(new_n974));
  AOI211_X1 g549(.A(G286), .B(new_n965), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G8), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n947), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n946), .B1(new_n977), .B2(KEYINPUT122), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n974), .ZN(new_n979));
  INV_X1    g554(.A(new_n965), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(G168), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(KEYINPUT122), .A3(new_n946), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n980), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(KEYINPUT123), .B2(G286), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n976), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT62), .B1(new_n978), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT123), .B1(new_n981), .B2(G8), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT122), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT51), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT62), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n965), .B1(new_n973), .B2(new_n974), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n991), .B1(new_n947), .B2(G168), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n946), .A2(KEYINPUT122), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n991), .B2(G168), .ZN(new_n994));
  OAI21_X1  g569(.A(G8), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n989), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  NOR2_X1   g572(.A1(G288), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n962), .B2(new_n849), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n952), .A2(new_n1001), .A3(new_n957), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1002), .A2(KEYINPUT112), .A3(G8), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT112), .B1(new_n1002), .B2(G8), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n999), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(KEYINPUT112), .A3(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n998), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1005), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n594), .A2(new_n1015), .A3(new_n599), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n598), .A2(G651), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n536), .A2(G48), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n591), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G1981), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1020), .A3(KEYINPUT49), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT49), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1016), .A2(new_n1020), .A3(KEYINPUT113), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT114), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1022), .A2(new_n1028), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n956), .A2(KEYINPUT109), .A3(new_n479), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT109), .B1(new_n956), .B2(new_n479), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n959), .B1(new_n510), .B2(new_n518), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n850), .A2(KEYINPUT45), .A3(new_n959), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1037), .A2(new_n706), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n850), .A2(new_n959), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n958), .B(new_n959), .C1(new_n510), .C2(new_n518), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(new_n952), .A4(new_n957), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1042), .A2(G2090), .ZN(new_n1043));
  OAI21_X1  g618(.A(G8), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G303), .A2(G8), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1045), .B(KEYINPUT55), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1037), .A2(new_n706), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1032), .A2(new_n1049), .A3(new_n960), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(G2090), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1046), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1052), .A3(G8), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1013), .A2(new_n1029), .A3(new_n1047), .A4(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1032), .A2(KEYINPUT119), .A3(new_n1049), .A4(new_n960), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(new_n961), .B2(new_n964), .ZN(new_n1057));
  INV_X1    g632(.A(G1961), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1037), .B2(G2078), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(G2078), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n969), .A2(new_n971), .A3(new_n972), .A4(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G171), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1054), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n986), .A2(new_n996), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n989), .A2(new_n995), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT54), .B1(new_n1064), .B2(G171), .ZN(new_n1069));
  INV_X1    g644(.A(new_n950), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n970), .A2(new_n1070), .A3(new_n1062), .A4(new_n1036), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1061), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1059), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1059), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1069), .B1(new_n1076), .B2(G171), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(new_n1054), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n952), .A2(new_n957), .A3(new_n1036), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n963), .B2(new_n959), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT120), .B(G1996), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT58), .B(G1341), .Z(new_n1083));
  AND2_X1   g658(.A1(new_n1002), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n569), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1086));
  NAND2_X1  g661(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1055), .A2(new_n1057), .A3(new_n793), .ZN(new_n1089));
  INV_X1    g664(.A(G2067), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n952), .A2(new_n1090), .A3(new_n1001), .A4(new_n957), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1091), .B(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1002), .A2(new_n1083), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1037), .B2(new_n1081), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1097), .A2(KEYINPUT121), .A3(KEYINPUT59), .A4(new_n569), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1088), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1089), .A2(new_n1093), .A3(new_n900), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n900), .B1(new_n1089), .B2(new_n1093), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1956), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1042), .A2(new_n1103), .ZN(new_n1104));
  AND3_X1   g679(.A1(G299), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .A4(new_n1108), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1104), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT61), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1107), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1104), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1099), .A2(new_n1102), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1111), .B1(new_n1101), .B2(new_n1117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1065), .B1(new_n1076), .B2(G171), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT54), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1068), .A2(new_n1078), .A3(new_n1122), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1053), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(new_n1013), .A3(new_n1029), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1016), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(G1976), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1129), .B1(new_n1029), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1014), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n983), .A2(G8), .A3(G168), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1054), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1051), .A2(G8), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT116), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1051), .A2(new_n1139), .A3(G8), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1046), .A3(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1012), .B1(new_n1028), .B2(new_n1022), .ZN(new_n1142));
  NOR4_X1   g717(.A1(new_n991), .A2(new_n1134), .A3(new_n976), .A4(G286), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1141), .A2(new_n1142), .A3(new_n1053), .A4(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1133), .B1(new_n1136), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1067), .A2(new_n1126), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n967), .A2(new_n970), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT111), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(G1996), .A3(new_n768), .ZN(new_n1149));
  INV_X1    g724(.A(G1996), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1151), .A2(new_n768), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n743), .B(G2067), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1148), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1149), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1148), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n724), .A2(new_n727), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n724), .A2(new_n727), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1155), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(G290), .A2(G1986), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(KEYINPUT110), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(KEYINPUT110), .B2(new_n1163), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1165), .A2(new_n970), .A3(new_n967), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1146), .A2(new_n1167), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n743), .A2(G2067), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1156), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1171), .A2(KEYINPUT125), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1171), .A2(KEYINPUT125), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1161), .A2(new_n1147), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT48), .Z(new_n1175));
  OAI21_X1  g750(.A(new_n1148), .B1(new_n768), .B2(new_n1153), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1151), .B(KEYINPUT46), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1178), .A2(KEYINPUT47), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1178), .A2(KEYINPUT47), .ZN(new_n1180));
  OAI22_X1  g755(.A1(new_n1160), .A2(new_n1175), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1172), .A2(new_n1173), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1168), .A2(new_n1182), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g758(.A1(G227), .A2(new_n461), .ZN(new_n1185));
  AND2_X1   g759(.A1(new_n656), .A2(new_n1185), .ZN(new_n1186));
  OR2_X1    g760(.A1(new_n1186), .A2(KEYINPUT126), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT126), .ZN(new_n1188));
  AND3_X1   g762(.A1(new_n698), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  OAI21_X1  g763(.A(new_n1189), .B1(new_n879), .B2(new_n887), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1190), .A2(new_n944), .ZN(G308));
  NAND2_X1  g765(.A1(new_n892), .A2(new_n886), .ZN(new_n1192));
  AND2_X1   g766(.A1(new_n937), .A2(new_n938), .ZN(new_n1193));
  AND2_X1   g767(.A1(new_n940), .A2(new_n943), .ZN(new_n1194));
  OAI211_X1 g768(.A(new_n1192), .B(new_n1189), .C1(new_n1193), .C2(new_n1194), .ZN(G225));
endmodule


