//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1305, new_n1306, new_n1307, new_n1308, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n213));
  NAND3_X1  g0013(.A1(new_n212), .A2(G50), .A3(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n206), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT66), .Z(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n218), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n206), .B1(new_n201), .B2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n206), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n248), .A2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT8), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT8), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI211_X1 g0057(.A(new_n247), .B(new_n251), .C1(new_n252), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n216), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n205), .A2(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G50), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n265), .A2(new_n268), .B1(new_n246), .B2(new_n264), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(new_n276), .A3(G274), .ZN(new_n277));
  INV_X1    g0077(.A(G226), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT3), .B(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G222), .A2(G1698), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(G223), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n276), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n281), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(G169), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n271), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n257), .A2(new_n298), .B1(G20), .B2(G77), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT68), .ZN(new_n300));
  INV_X1    g0100(.A(new_n252), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT15), .B(G87), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n299), .A2(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n299), .A2(new_n300), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n260), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n291), .B1(new_n205), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n265), .A2(new_n306), .B1(new_n291), .B2(new_n264), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n282), .A2(G238), .A3(G1698), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n282), .A2(G232), .A3(new_n284), .ZN(new_n312));
  INV_X1    g0112(.A(G107), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n311), .B(new_n312), .C1(new_n313), .C2(new_n282), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n280), .ZN(new_n317));
  INV_X1    g0117(.A(G274), .ZN(new_n318));
  INV_X1    g0118(.A(new_n216), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(new_n275), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n317), .A2(G244), .B1(new_n320), .B2(new_n274), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n309), .B1(new_n310), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n322), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n297), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n305), .A2(new_n307), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n324), .A2(new_n294), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G68), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n264), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT71), .ZN(new_n336));
  OR3_X1    g0136(.A1(new_n335), .A2(new_n336), .A3(KEYINPUT12), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n335), .A2(KEYINPUT12), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n336), .B1(new_n335), .B2(KEYINPUT12), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n265), .A2(G68), .A3(new_n266), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n298), .A2(G50), .B1(G20), .B2(new_n334), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n301), .B2(new_n291), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT11), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(new_n260), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n344), .B1(new_n343), .B2(new_n260), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n340), .B(new_n341), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n278), .A2(new_n284), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n230), .A2(G1698), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n282), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n315), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT13), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n317), .A2(G238), .B1(new_n320), .B2(new_n274), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n276), .B1(new_n351), .B2(new_n352), .ZN(new_n358));
  INV_X1    g0158(.A(G238), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n277), .B1(new_n359), .B2(new_n280), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT13), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(KEYINPUT70), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT70), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(KEYINPUT13), .C1(new_n358), .C2(new_n360), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n357), .A2(G190), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n348), .B1(new_n362), .B2(new_n325), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n357), .A2(G179), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n328), .B1(new_n357), .B2(new_n361), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n366), .A2(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n347), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(KEYINPUT9), .B(new_n269), .C1(new_n258), .C2(new_n261), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT69), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n271), .A2(KEYINPUT9), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n293), .A2(G190), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n325), .B2(new_n293), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT10), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n377), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI221_X1 g0183(.A(new_n379), .B1(new_n325), .B2(new_n293), .C1(new_n271), .C2(KEYINPUT9), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT10), .B1(new_n384), .B2(new_n376), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n333), .A2(new_n368), .A3(new_n374), .A4(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(G1698), .ZN(new_n388));
  AND2_X1   g0188(.A1(KEYINPUT4), .A2(G244), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n287), .A2(new_n289), .A3(new_n389), .A4(new_n284), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G283), .ZN(new_n391));
  AND3_X1   g0191(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT4), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT72), .B1(new_n288), .B2(G33), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT72), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(new_n248), .A3(KEYINPUT3), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n394), .A2(new_n396), .A3(new_n284), .A4(new_n289), .ZN(new_n397));
  INV_X1    g0197(.A(G244), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n276), .B1(new_n392), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n273), .A2(G1), .ZN(new_n401));
  XNOR2_X1  g0201(.A(KEYINPUT5), .B(G41), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n315), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G257), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n402), .A2(G274), .A3(new_n276), .A4(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(G169), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  AND2_X1   g0207(.A1(KEYINPUT5), .A2(G41), .ZN(new_n408));
  NOR2_X1   g0208(.A1(KEYINPUT5), .A2(G41), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n401), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n403), .A2(G257), .B1(new_n411), .B2(new_n320), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n388), .A2(new_n390), .A3(new_n391), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n288), .A2(KEYINPUT72), .A3(G33), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n248), .A2(KEYINPUT3), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n416), .A2(G244), .A3(new_n284), .A4(new_n394), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(new_n393), .ZN(new_n418));
  OAI211_X1 g0218(.A(G179), .B(new_n412), .C1(new_n418), .C2(new_n276), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n407), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT81), .ZN(new_n421));
  NAND2_X1  g0221(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n282), .B2(G20), .ZN(new_n423));
  XNOR2_X1  g0223(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n290), .A2(new_n424), .A3(new_n206), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G107), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n249), .A2(new_n291), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT6), .ZN(new_n429));
  INV_X1    g0229(.A(G97), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n313), .ZN(new_n431));
  NOR2_X1   g0231(.A1(G97), .A2(G107), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n429), .A2(new_n430), .A3(G107), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n428), .B1(new_n436), .B2(G20), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n261), .B1(new_n427), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n263), .A2(G97), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n205), .A2(G33), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n261), .A2(new_n263), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n441), .B2(G97), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n421), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g0244(.A(G97), .B(G107), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n434), .B1(new_n445), .B2(new_n429), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n446), .A2(new_n206), .B1(new_n291), .B2(new_n249), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n313), .B1(new_n423), .B2(new_n425), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n260), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(KEYINPUT81), .A3(new_n442), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n420), .A2(new_n444), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT82), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT82), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n420), .A2(new_n444), .A3(new_n453), .A4(new_n450), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n400), .A2(new_n406), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT80), .B1(new_n455), .B2(new_n325), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT80), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n457), .B(G200), .C1(new_n400), .C2(new_n406), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n449), .A2(new_n442), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(G190), .B2(new_n455), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n452), .A2(new_n454), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n394), .A2(new_n396), .A3(new_n289), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(G257), .A3(new_n284), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT84), .ZN(new_n465));
  AND2_X1   g0265(.A1(G264), .A2(G1698), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n290), .A2(G303), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n394), .A2(new_n396), .A3(new_n289), .A4(new_n466), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT84), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n410), .A2(G270), .A3(new_n276), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n405), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT83), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT83), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n475), .A3(new_n405), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n471), .A2(new_n315), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G190), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n469), .B(new_n465), .ZN(new_n479));
  INV_X1    g0279(.A(new_n397), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(G257), .B1(G303), .B2(new_n290), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n276), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n476), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n475), .B1(new_n472), .B2(new_n405), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(G200), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n391), .B(new_n206), .C1(G33), .C2(new_n430), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n260), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT20), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n263), .A2(G116), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n493), .B1(new_n441), .B2(G116), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n478), .A2(new_n486), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n490), .B(KEYINPUT20), .ZN(new_n499));
  INV_X1    g0299(.A(new_n493), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n265), .A2(new_n440), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(new_n488), .ZN(new_n502));
  OAI21_X1  g0302(.A(G169), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n498), .B1(new_n477), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n477), .A2(G179), .A3(new_n495), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n328), .B1(new_n492), .B2(new_n494), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n506), .B(KEYINPUT21), .C1(new_n482), .C2(new_n485), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n206), .B1(new_n352), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(G87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n432), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n206), .A2(G33), .A3(G97), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n510), .A2(new_n512), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n394), .A2(new_n396), .A3(new_n206), .A4(new_n289), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n514), .B1(new_n334), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(new_n260), .B1(new_n264), .B2(new_n302), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n501), .A2(new_n302), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n276), .A2(G274), .A3(new_n401), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n205), .A2(G45), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n276), .A2(G250), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n394), .A2(new_n396), .A3(new_n289), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n398), .A2(G1698), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(G238), .B2(G1698), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n523), .A2(new_n525), .B1(new_n248), .B2(new_n488), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n522), .B1(new_n526), .B2(new_n315), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n517), .A2(new_n518), .B1(new_n527), .B2(new_n294), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n315), .ZN(new_n529));
  INV_X1    g0329(.A(new_n522), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n328), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n516), .A2(new_n260), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n302), .A2(new_n264), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n441), .A2(G87), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(G200), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n527), .A2(G190), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n533), .A2(new_n540), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n497), .A2(new_n508), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n410), .A2(G264), .A3(new_n276), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT86), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT86), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n410), .A2(new_n545), .A3(G264), .A4(new_n276), .ZN(new_n546));
  INV_X1    g0346(.A(G257), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G1698), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G250), .B2(G1698), .ZN(new_n549));
  INV_X1    g0349(.A(G294), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n523), .A2(new_n549), .B1(new_n248), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n544), .A2(new_n546), .B1(new_n551), .B2(new_n315), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n552), .A2(new_n294), .A3(new_n405), .ZN(new_n553));
  AOI21_X1  g0353(.A(G169), .B1(new_n552), .B2(new_n405), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(KEYINPUT22), .B1(new_n515), .B2(new_n511), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n511), .A2(KEYINPUT22), .A3(G20), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n282), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT85), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n282), .A2(KEYINPUT85), .A3(new_n557), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n556), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n248), .A2(new_n488), .A3(G20), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n206), .B2(G107), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n313), .A2(KEYINPUT23), .A3(G20), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n562), .A2(new_n570), .A3(new_n567), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n261), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n313), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT25), .B1(new_n264), .B2(new_n313), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n501), .A2(new_n313), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n555), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT87), .ZN(new_n578));
  AND3_X1   g0378(.A1(new_n562), .A2(new_n570), .A3(new_n567), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n570), .B1(new_n562), .B2(new_n567), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n260), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n544), .A2(new_n546), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n551), .A2(new_n315), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n405), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n325), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n552), .A2(new_n310), .A3(new_n405), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n576), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n581), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n577), .A2(new_n578), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n578), .B1(new_n577), .B2(new_n589), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n462), .B(new_n542), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n265), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n257), .A2(new_n266), .ZN(new_n594));
  OAI22_X1  g0394(.A1(new_n593), .A2(new_n594), .B1(new_n263), .B2(new_n257), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT74), .ZN(new_n596));
  INV_X1    g0396(.A(G159), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n249), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G58), .A2(G68), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n202), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n596), .B(new_n599), .C1(new_n601), .C2(new_n206), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n206), .B1(new_n202), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT74), .B1(new_n603), .B2(new_n598), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n523), .A2(new_n206), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT7), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n523), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(KEYINPUT73), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT7), .B1(new_n523), .B2(new_n206), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT73), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n334), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n605), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n261), .B1(new_n614), .B2(KEYINPUT16), .ZN(new_n615));
  XNOR2_X1  g0415(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n334), .B1(new_n423), .B2(new_n425), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n616), .B1(new_n605), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n595), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT77), .ZN(new_n620));
  NOR2_X1   g0420(.A1(G223), .A2(G1698), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n278), .B2(G1698), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n416), .A2(new_n394), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(G33), .A2(G87), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n620), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n278), .A2(G1698), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(G223), .B2(G1698), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n620), .B(new_n624), .C1(new_n523), .C2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n315), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(KEYINPUT78), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n276), .A2(G232), .A3(new_n279), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n277), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(KEYINPUT79), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(KEYINPUT79), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n635), .A2(new_n636), .A3(G179), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n624), .B1(new_n523), .B2(new_n627), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT77), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n628), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT78), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n315), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n631), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n630), .A2(new_n634), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n328), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT18), .B1(new_n619), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT17), .ZN(new_n648));
  AOI21_X1  g0448(.A(G200), .B1(new_n630), .B2(new_n634), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n641), .B1(new_n640), .B2(new_n315), .ZN(new_n650));
  AOI211_X1 g0450(.A(KEYINPUT78), .B(new_n276), .C1(new_n639), .C2(new_n628), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n635), .A2(new_n636), .A3(G190), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n602), .A2(new_n604), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n523), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n656), .A2(new_n611), .A3(new_n612), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n606), .A2(new_n612), .A3(new_n607), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G68), .ZN(new_n659));
  OAI211_X1 g0459(.A(KEYINPUT16), .B(new_n655), .C1(new_n657), .C2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(new_n260), .A3(new_n618), .ZN(new_n661));
  INV_X1    g0461(.A(new_n595), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n648), .B1(new_n654), .B2(new_n663), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n652), .A2(new_n637), .B1(new_n644), .B2(new_n328), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT18), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n663), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n631), .A2(new_n653), .A3(new_n642), .ZN(new_n668));
  INV_X1    g0468(.A(new_n649), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n619), .A2(new_n670), .A3(KEYINPUT17), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n647), .A2(new_n664), .A3(new_n667), .A4(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n387), .A2(new_n592), .A3(new_n672), .ZN(G372));
  INV_X1    g0473(.A(new_n297), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n647), .A2(new_n667), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n368), .A2(new_n332), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n374), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT91), .Z(new_n678));
  NAND2_X1  g0478(.A1(new_n664), .A2(new_n671), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT92), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n386), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT92), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n674), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n387), .A2(new_n672), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT26), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n420), .A2(KEYINPUT90), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n407), .A2(new_n419), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n460), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT88), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n522), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT88), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n693), .A2(new_n694), .B1(new_n526), .B2(new_n315), .ZN(new_n695));
  OAI21_X1  g0495(.A(KEYINPUT89), .B1(new_n695), .B2(G169), .ZN(new_n696));
  INV_X1    g0496(.A(new_n694), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT88), .B1(new_n519), .B2(new_n521), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n529), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT89), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(new_n328), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n528), .A3(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n537), .B(new_n539), .C1(new_n325), .C2(new_n695), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n687), .B1(new_n691), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n533), .A2(new_n540), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n452), .A2(KEYINPUT26), .A3(new_n706), .A4(new_n454), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n452), .A2(new_n454), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n459), .A2(new_n461), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n702), .A2(new_n703), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n584), .A2(new_n328), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n552), .A2(new_n294), .A3(new_n405), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n581), .B2(new_n588), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n712), .B(new_n589), .C1(new_n716), .C2(new_n508), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n702), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n686), .B1(new_n708), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n685), .A2(new_n719), .ZN(G369));
  NOR2_X1   g0520(.A1(new_n572), .A2(new_n576), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  OAI21_X1  g0523(.A(G213), .B1(new_n722), .B2(KEYINPUT27), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G343), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n590), .A2(new_n591), .B1(new_n721), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT94), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n716), .A2(new_n729), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n497), .A2(new_n508), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n730), .A2(new_n496), .ZN(new_n738));
  MUX2_X1   g0538(.A(new_n737), .B(new_n508), .S(new_n738), .Z(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n716), .A2(new_n730), .ZN(new_n743));
  INV_X1    g0543(.A(new_n508), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n729), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n733), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(G399));
  NAND2_X1  g0547(.A1(new_n209), .A2(new_n272), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n512), .A2(G116), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n748), .A2(G1), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n214), .B2(new_n748), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT28), .ZN(new_n752));
  INV_X1    g0552(.A(G330), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT96), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(KEYINPUT30), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n552), .A2(KEYINPUT95), .A3(new_n527), .ZN(new_n756));
  AOI21_X1  g0556(.A(KEYINPUT95), .B1(new_n552), .B2(new_n527), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n477), .A2(G179), .A3(new_n455), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n695), .B(KEYINPUT97), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n477), .A2(new_n455), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n761), .A2(new_n762), .A3(new_n294), .A4(new_n584), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT95), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n582), .A2(new_n583), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n765), .B2(new_n531), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n552), .A2(KEYINPUT95), .A3(new_n527), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n482), .A2(new_n485), .A3(new_n294), .ZN(new_n769));
  INV_X1    g0569(.A(new_n755), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n768), .A2(new_n769), .A3(new_n455), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n760), .A2(new_n763), .A3(new_n771), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n772), .A2(KEYINPUT31), .A3(new_n729), .ZN(new_n773));
  AOI21_X1  g0573(.A(KEYINPUT31), .B1(new_n772), .B2(new_n729), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g0575(.A1(new_n581), .A2(new_n587), .A3(new_n588), .ZN(new_n776));
  OAI21_X1  g0576(.A(KEYINPUT87), .B1(new_n776), .B2(new_n716), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n577), .A2(new_n578), .A3(new_n589), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n779), .A2(new_n462), .A3(new_n542), .A4(new_n730), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n753), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n711), .A2(KEYINPUT98), .ZN(new_n782));
  INV_X1    g0582(.A(new_n717), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT98), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n462), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(KEYINPUT26), .B1(new_n691), .B2(new_n704), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n452), .A2(new_n687), .A3(new_n706), .A4(new_n454), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n787), .A2(new_n788), .A3(new_n702), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n729), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT29), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n730), .B1(new_n718), .B2(new_n708), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT29), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n781), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n752), .B1(new_n796), .B2(G1), .ZN(G364));
  INV_X1    g0597(.A(new_n748), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n206), .A2(G13), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n205), .B1(new_n799), .B2(G45), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n741), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G330), .B2(new_n739), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n216), .B1(G20), .B2(new_n328), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n206), .A2(G179), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(new_n310), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G107), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G179), .A2(G200), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n206), .B1(new_n811), .B2(G190), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n206), .A2(G190), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n811), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n597), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT32), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n810), .B1(new_n430), .B2(new_n812), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n206), .A2(new_n294), .A3(G190), .A4(G200), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR4_X1   g0619(.A1(new_n206), .A2(new_n294), .A3(new_n310), .A4(G200), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n282), .B1(new_n819), .B2(new_n291), .C1(new_n821), .C2(new_n253), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n815), .A2(new_n816), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n807), .A2(G190), .A3(G200), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n511), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n817), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n827));
  OR2_X1    g0627(.A1(new_n827), .A2(KEYINPUT100), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(KEYINPUT100), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n828), .A2(G190), .A3(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n828), .A2(new_n310), .A3(new_n829), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G50), .A2(new_n831), .B1(new_n833), .B2(G68), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT33), .B(G317), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G326), .A2(new_n831), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n282), .B1(new_n820), .B2(G322), .ZN(new_n837));
  INV_X1    g0637(.A(new_n814), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G329), .B1(new_n818), .B2(G311), .ZN(new_n839));
  INV_X1    g0639(.A(G283), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n808), .A2(new_n840), .B1(new_n812), .B2(new_n550), .ZN(new_n841));
  INV_X1    g0641(.A(new_n824), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(G303), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n836), .A2(new_n837), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT101), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n826), .A2(new_n834), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n806), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n209), .A2(new_n282), .ZN(new_n849));
  INV_X1    g0649(.A(G355), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n850), .B1(G116), .B2(new_n209), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n244), .A2(G45), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT99), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n209), .A2(new_n523), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n215), .B2(new_n273), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n851), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(G13), .A2(G33), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(G20), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n805), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n802), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n848), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n859), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n739), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n804), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G396));
  NOR2_X1   g0667(.A1(new_n808), .A2(new_n511), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n869), .B1(new_n430), .B2(new_n812), .C1(new_n313), .C2(new_n824), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n290), .B1(new_n819), .B2(new_n488), .ZN(new_n871));
  INV_X1    g0671(.A(G311), .ZN(new_n872));
  OAI22_X1  g0672(.A1(new_n821), .A2(new_n550), .B1(new_n814), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G303), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n840), .A2(new_n832), .B1(new_n830), .B2(new_n874), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n870), .A2(new_n871), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT102), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n820), .A2(G143), .B1(new_n818), .B2(G159), .ZN(new_n878));
  INV_X1    g0678(.A(G137), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n878), .B1(new_n879), .B2(new_n830), .C1(new_n250), .C2(new_n832), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT34), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n881), .ZN(new_n883));
  INV_X1    g0683(.A(G132), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n463), .B1(new_n884), .B2(new_n814), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n808), .A2(new_n334), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n824), .A2(new_n246), .B1(new_n812), .B2(new_n253), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n882), .A2(new_n883), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n805), .B1(new_n877), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n802), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n805), .A2(new_n857), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n291), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n331), .A2(new_n729), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n323), .A2(new_n326), .B1(new_n309), .B2(new_n730), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n895), .B2(new_n331), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n890), .B(new_n893), .C1(new_n896), .C2(new_n858), .ZN(new_n897));
  INV_X1    g0697(.A(new_n896), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n793), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n730), .B(new_n896), .C1(new_n718), .C2(new_n708), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n781), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n781), .A3(new_n900), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n891), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(G384));
  OAI21_X1  g0706(.A(new_n655), .B1(new_n657), .B2(new_n659), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n616), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n595), .B1(new_n615), .B2(new_n908), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n663), .A2(new_n654), .B1(new_n909), .B2(new_n727), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n646), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n665), .A2(new_n663), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n619), .A2(new_n670), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  INV_X1    g0715(.A(new_n727), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n663), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n913), .A2(new_n914), .A3(new_n915), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n909), .A2(new_n727), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n672), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n913), .A2(new_n914), .A3(new_n917), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  INV_X1    g0724(.A(new_n917), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n924), .A2(new_n918), .B1(new_n672), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n922), .B1(KEYINPUT38), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT39), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n374), .A2(new_n729), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n919), .A2(new_n921), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(KEYINPUT39), .A3(new_n922), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n675), .A2(new_n916), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n922), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n374), .A2(new_n368), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n729), .A2(new_n347), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT104), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT104), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n939), .B(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(new_n374), .A3(new_n368), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n894), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n900), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n936), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n935), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n792), .A2(new_n686), .A3(new_n795), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n685), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n941), .A2(new_n896), .A3(new_n944), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n775), .B2(new_n780), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n919), .A2(KEYINPUT38), .A3(new_n921), .ZN(new_n955));
  AOI21_X1  g0755(.A(KEYINPUT38), .B1(new_n919), .B2(new_n921), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT40), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n958), .B(new_n953), .C1(new_n775), .C2(new_n780), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n957), .A2(new_n958), .B1(new_n927), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n772), .A2(new_n729), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT31), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n772), .A2(KEYINPUT31), .A3(new_n729), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n592), .C2(new_n729), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n686), .ZN(new_n967));
  OAI21_X1  g0767(.A(G330), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n967), .B2(new_n961), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n952), .A2(new_n969), .B1(new_n205), .B2(new_n799), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n952), .B2(new_n969), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n436), .A2(KEYINPUT35), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(G116), .A3(new_n217), .A4(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT36), .Z(new_n975));
  NAND3_X1  g0775(.A1(new_n215), .A2(G77), .A3(new_n600), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n246), .A2(G68), .ZN(new_n977));
  AOI211_X1 g0777(.A(new_n205), .B(G13), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n971), .A2(new_n975), .A3(new_n978), .ZN(G367));
  XOR2_X1   g0779(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n980));
  NOR2_X1   g0780(.A1(new_n730), .A2(new_n537), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n712), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n702), .B2(new_n982), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n980), .B1(new_n984), .B2(KEYINPUT105), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(KEYINPUT105), .B2(new_n984), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n729), .A2(new_n460), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n782), .A2(new_n785), .A3(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n691), .A2(new_n730), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n709), .B1(new_n994), .B2(new_n577), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n730), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n733), .A2(new_n745), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n989), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n987), .A2(KEYINPUT107), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n988), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n742), .A2(new_n994), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1001), .A2(new_n1002), .A3(new_n988), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n748), .B(KEYINPUT41), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n1011));
  NAND2_X1  g0811(.A1(new_n746), .A2(new_n743), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT109), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n1013), .A3(new_n994), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1013), .B1(new_n1012), .B2(new_n994), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1016), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1011), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1018), .A2(new_n1014), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n746), .A2(new_n743), .A3(new_n993), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT45), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1017), .A2(new_n1020), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n742), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1017), .A2(new_n1020), .A3(new_n742), .A4(new_n1023), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT110), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n731), .A2(KEYINPUT94), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n731), .A2(KEYINPUT94), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n735), .B1(new_n744), .B2(new_n729), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n746), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(new_n741), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n1033), .B2(new_n796), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1032), .A2(new_n741), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n740), .B1(new_n1031), .B2(new_n746), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1028), .B(new_n796), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1026), .A2(new_n1027), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1010), .B1(new_n1040), .B2(new_n796), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1009), .B1(new_n1041), .B2(new_n801), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n860), .B1(new_n209), .B2(new_n302), .C1(new_n236), .C2(new_n854), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n802), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n809), .A2(G77), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n253), .B2(new_n824), .C1(new_n334), .C2(new_n812), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n820), .A2(G150), .B1(new_n818), .B2(G50), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n282), .C1(new_n879), .C2(new_n814), .ZN(new_n1049));
  INV_X1    g0849(.A(G143), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1050), .A2(new_n830), .B1(new_n832), .B2(new_n597), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1047), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT112), .Z(new_n1053));
  AOI22_X1  g0853(.A1(G317), .A2(new_n838), .B1(new_n820), .B2(G303), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n824), .A2(new_n488), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1054), .B1(KEYINPUT46), .B2(new_n1055), .C1(new_n840), .C2(new_n819), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(KEYINPUT46), .B2(new_n1055), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n808), .A2(new_n430), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n523), .B1(new_n313), .B2(new_n812), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G311), .C2(new_n831), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(new_n550), .C2(new_n832), .ZN(new_n1061));
  AOI21_X1  g0861(.A(KEYINPUT47), .B1(new_n1053), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1062), .A2(new_n806), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1053), .A2(KEYINPUT47), .A3(new_n1061), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1045), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n864), .B2(new_n984), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1042), .A2(new_n1066), .ZN(G387));
  AOI21_X1  g0867(.A(new_n748), .B1(new_n1033), .B2(new_n796), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n796), .B2(new_n1033), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n849), .A2(new_n749), .B1(G107), .B2(new_n209), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n854), .B1(new_n233), .B2(G45), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n749), .B(new_n273), .C1(new_n334), .C2(new_n291), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n257), .A2(new_n246), .ZN(new_n1074));
  XOR2_X1   g0874(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1075));
  XNOR2_X1  g0875(.A(new_n1074), .B(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1072), .A2(KEYINPUT113), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1070), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n821), .A2(new_n246), .B1(new_n819), .B2(new_n334), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G150), .B2(new_n838), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n824), .A2(new_n291), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n812), .A2(new_n302), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1058), .A2(new_n1082), .A3(new_n1083), .A4(new_n523), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n257), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1081), .B(new_n1084), .C1(new_n1085), .C2(new_n832), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n830), .A2(new_n597), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT115), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n812), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n842), .A2(G294), .B1(new_n1090), .B2(G283), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n820), .A2(G317), .B1(new_n818), .B2(G303), .ZN(new_n1092));
  INV_X1    g0892(.A(G322), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1092), .B1(new_n872), .B2(new_n832), .C1(new_n1093), .C2(new_n830), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT116), .Z(new_n1095));
  OAI21_X1  g0895(.A(new_n1091), .B1(new_n1095), .B2(KEYINPUT48), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(KEYINPUT48), .B2(new_n1095), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(KEYINPUT49), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n463), .B1(G326), .B2(new_n838), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n488), .B2(new_n808), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n1097), .B2(KEYINPUT49), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1089), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n802), .B1(new_n861), .B2(new_n1079), .C1(new_n1102), .C2(new_n806), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT117), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n734), .A2(new_n735), .A3(new_n859), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1033), .A2(new_n801), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1069), .A2(new_n1106), .ZN(G393));
  AND2_X1   g0907(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1033), .A2(new_n796), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n798), .B(new_n1040), .C1(new_n1108), .C2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1026), .A2(new_n801), .A3(new_n1027), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n241), .A2(new_n854), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n860), .B1(new_n430), .B2(new_n209), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n802), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n831), .A2(G317), .B1(G311), .B2(new_n820), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT52), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n832), .A2(new_n874), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n290), .B1(new_n1093), .B2(new_n814), .C1(new_n819), .C2(new_n550), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n810), .B1(new_n488), .B2(new_n812), .C1(new_n840), .C2(new_n824), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(KEYINPUT118), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n250), .A2(new_n830), .B1(new_n821), .B2(new_n597), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT51), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n463), .B1(new_n1050), .B2(new_n814), .C1(new_n819), .C2(new_n1085), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n824), .A2(new_n334), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n812), .A2(new_n291), .ZN(new_n1127));
  NOR4_X1   g0927(.A1(new_n1125), .A2(new_n868), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1124), .B(new_n1128), .C1(new_n246), .C2(new_n832), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1121), .A2(new_n1122), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1114), .B1(new_n1130), .B2(new_n805), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n993), .B2(new_n864), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1111), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1110), .A2(new_n1134), .ZN(G390));
  INV_X1    g0935(.A(new_n945), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n781), .A2(new_n896), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n900), .A2(new_n946), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1136), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n930), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n929), .A2(new_n934), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n895), .A2(new_n331), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n709), .A2(new_n784), .A3(new_n710), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n784), .B1(new_n709), .B2(new_n710), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1143), .A2(new_n1144), .A3(new_n717), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n730), .B(new_n1142), .C1(new_n1145), .C2(new_n789), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n945), .B1(new_n1146), .B2(new_n946), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n927), .A2(new_n1140), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1137), .B1(new_n1141), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n924), .A2(new_n918), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n672), .A2(new_n925), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n932), .ZN(new_n1154));
  AOI21_X1  g0954(.A(KEYINPUT39), .B1(new_n1154), .B2(new_n922), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n955), .A2(new_n956), .A3(new_n928), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n1155), .A2(new_n1156), .B1(new_n930), .B2(new_n947), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n894), .B1(new_n791), .B2(new_n1142), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1140), .B(new_n927), .C1(new_n1158), .C2(new_n945), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n781), .A2(new_n896), .A3(new_n1136), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1150), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1136), .B1(new_n781), .B2(new_n896), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1138), .B1(new_n1137), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n898), .B1(new_n781), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n966), .A2(G330), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(KEYINPUT119), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1136), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1164), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n781), .A2(new_n686), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n685), .A2(new_n950), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(KEYINPUT120), .B1(new_n1162), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n896), .B1(new_n1167), .B2(KEYINPUT119), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n781), .A2(new_n1165), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n945), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1170), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1173), .B1(new_n1181), .B2(new_n1164), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT120), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1182), .A2(new_n1183), .A3(new_n1150), .A4(new_n1161), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1176), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n748), .B1(new_n1162), .B2(new_n1175), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1162), .A2(new_n800), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n857), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n892), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n802), .B1(new_n257), .B2(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1127), .B(new_n886), .C1(G87), .C2(new_n842), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G107), .A2(new_n833), .B1(new_n831), .B2(G283), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n282), .B1(new_n818), .B2(G97), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(G294), .A2(new_n838), .B1(new_n820), .B2(G116), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n824), .A2(new_n250), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT53), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT54), .B(G143), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n290), .B1(new_n1200), .B2(new_n818), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G125), .A2(new_n838), .B1(new_n820), .B2(G132), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n809), .A2(G50), .B1(new_n1090), .B2(G159), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1198), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(G128), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1205), .A2(new_n830), .B1(new_n832), .B2(new_n879), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1196), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1191), .B1(new_n1207), .B2(new_n805), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1188), .B1(new_n1189), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1187), .A2(new_n1209), .ZN(G378));
  NAND2_X1  g1010(.A1(new_n1185), .A2(new_n1174), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n935), .A2(new_n948), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n957), .A2(new_n958), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n682), .A2(new_n297), .A3(new_n683), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n271), .A2(new_n727), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1215), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n682), .A2(new_n297), .A3(new_n683), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1216), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n959), .A2(new_n927), .ZN(new_n1225));
  AND4_X1   g1025(.A1(G330), .A2(new_n1213), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1224), .B1(new_n960), .B2(G330), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1212), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1213), .A2(G330), .A3(new_n1225), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1224), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n960), .A2(G330), .A3(new_n1224), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1232), .A2(new_n949), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1228), .A2(new_n1229), .A3(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(KEYINPUT123), .B(new_n1212), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1211), .B2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1173), .B1(new_n1176), .B2(new_n1184), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1228), .A2(new_n1234), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT57), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n798), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1235), .A2(new_n801), .A3(new_n1236), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT124), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n891), .B1(new_n246), .B2(new_n892), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n523), .A2(new_n272), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n819), .A2(new_n302), .B1(new_n814), .B2(new_n840), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n1246), .B(new_n1247), .C1(G107), .C2(new_n820), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n812), .A2(new_n334), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1249), .B(new_n1082), .C1(G58), .C2(new_n809), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(G97), .A2(new_n833), .B1(new_n831), .B2(G116), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1248), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT58), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n1246), .B(new_n246), .C1(G33), .C2(G41), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n832), .A2(new_n884), .B1(new_n819), .B2(new_n879), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT121), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n842), .A2(new_n1200), .B1(new_n820), .B2(G128), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT122), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n831), .A2(G125), .B1(G150), .B2(new_n1090), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1259), .A2(new_n1261), .A3(new_n1262), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(KEYINPUT59), .ZN(new_n1264));
  AOI211_X1 g1064(.A(G33), .B(G41), .C1(new_n838), .C2(G124), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n597), .B2(new_n808), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1263), .B2(KEYINPUT59), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1254), .B(new_n1257), .C1(new_n1264), .C2(new_n1267), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1245), .B1(new_n806), .B2(new_n1268), .C1(new_n1224), .C2(new_n858), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1243), .A2(new_n1244), .A3(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1244), .B1(new_n1243), .B2(new_n1269), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1238), .A2(new_n1242), .B1(new_n1270), .B2(new_n1271), .ZN(G375));
  NAND3_X1  g1072(.A1(new_n1181), .A2(new_n1164), .A3(new_n1173), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1010), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1175), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1046), .B1(new_n430), .B2(new_n824), .C1(new_n302), .C2(new_n812), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n488), .A2(new_n832), .B1(new_n830), .B2(new_n550), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n290), .B1(new_n821), .B2(new_n840), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n819), .A2(new_n313), .B1(new_n814), .B2(new_n874), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1279), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n842), .A2(G159), .B1(new_n1090), .B2(G50), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1281), .B(new_n463), .C1(new_n253), .C2(new_n808), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n820), .A2(G137), .B1(new_n818), .B2(G150), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1205), .B2(new_n814), .ZN(new_n1284));
  OAI22_X1  g1084(.A1(new_n884), .A2(new_n830), .B1(new_n832), .B2(new_n1199), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1282), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n805), .B1(new_n1280), .B2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1287), .B(new_n802), .C1(G68), .C2(new_n1190), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(new_n945), .B2(new_n857), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1171), .B2(new_n801), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1275), .A2(new_n1290), .ZN(G381));
  NAND3_X1  g1091(.A1(new_n1069), .A2(new_n1106), .A3(new_n866), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1292), .A2(G384), .ZN(new_n1293));
  NOR4_X1   g1093(.A1(G390), .A2(G378), .A3(G381), .A4(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT57), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1239), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1241), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n748), .B1(new_n1211), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1243), .A2(new_n1269), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT124), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1243), .A2(new_n1244), .A3(new_n1269), .ZN(new_n1302));
  AOI22_X1  g1102(.A1(new_n1297), .A2(new_n1299), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1294), .A2(new_n1042), .A3(new_n1066), .A4(new_n1303), .ZN(G407));
  INV_X1    g1104(.A(G378), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n728), .A2(G213), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(G407), .A2(G213), .A3(new_n1308), .ZN(G409));
  NAND3_X1  g1109(.A1(new_n1211), .A2(new_n1274), .A3(new_n1237), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1240), .A2(new_n801), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1311), .A2(new_n1269), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1305), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(G375), .B2(new_n1305), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1273), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1316), .B1(KEYINPUT60), .B2(new_n1175), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1181), .A2(KEYINPUT60), .A3(new_n1164), .A4(new_n1173), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n798), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1290), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(G384), .B(new_n1290), .C1(new_n1317), .C2(new_n1319), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1315), .A2(new_n1306), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  OR2_X1    g1127(.A1(new_n1306), .A2(KEYINPUT125), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1322), .A2(new_n1323), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1307), .A2(G2897), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1329), .B(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G378), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1303), .B2(G378), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1331), .B1(new_n1333), .B2(new_n1307), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT62), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1315), .A2(new_n1335), .A3(new_n1306), .A4(new_n1324), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1326), .A2(new_n1327), .A3(new_n1334), .A4(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G393), .A2(G396), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1292), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1110), .A2(new_n1134), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1339), .B1(new_n1110), .B2(new_n1134), .ZN(new_n1341));
  OAI21_X1  g1141(.A(G387), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1339), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1040), .A2(new_n798), .ZN(new_n1344));
  AOI22_X1  g1144(.A1(new_n1026), .A2(new_n1027), .B1(new_n796), .B2(new_n1033), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1343), .B1(new_n1346), .B2(new_n1133), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1110), .A2(new_n1134), .A3(new_n1339), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1347), .A2(new_n1042), .A3(new_n1066), .A4(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT126), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1342), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1350), .B1(new_n1342), .B2(new_n1349), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1337), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1315), .A2(new_n1306), .ZN(new_n1355));
  AOI21_X1  g1155(.A(KEYINPUT61), .B1(new_n1355), .B2(new_n1331), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT63), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1325), .A2(new_n1357), .ZN(new_n1358));
  AND2_X1   g1158(.A1(new_n1342), .A2(new_n1349), .ZN(new_n1359));
  NAND4_X1  g1159(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1306), .A4(new_n1324), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1356), .A2(new_n1358), .A3(new_n1359), .A4(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1354), .A2(new_n1361), .ZN(G405));
  NAND2_X1  g1162(.A1(new_n1303), .A2(G378), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(G375), .A2(new_n1305), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1366));
  OR2_X1    g1166(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1365), .A2(new_n1366), .A3(new_n1367), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1363), .A2(KEYINPUT127), .A3(new_n1364), .A4(new_n1324), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1368), .A2(new_n1369), .ZN(new_n1370));
  XNOR2_X1  g1170(.A(new_n1370), .B(new_n1359), .ZN(G402));
endmodule


