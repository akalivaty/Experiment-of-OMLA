//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  XNOR2_X1  g002(.A(G127gat), .B(G134gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT74), .A2(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G113gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G120gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT72), .A2(G120gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n211), .B1(new_n214), .B2(G113gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n208), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT72), .B(G120gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n210), .B1(new_n218), .B2(new_n209), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT73), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n205), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n223), .B(new_n225), .C1(new_n226), .C2(KEYINPUT2), .ZN(new_n227));
  INV_X1    g026(.A(G148gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G141gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT81), .B(G148gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n229), .B1(new_n230), .B2(G141gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n224), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n233), .A2(new_n223), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n227), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT4), .B1(new_n222), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(KEYINPUT82), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n227), .B(new_n238), .C1(new_n231), .C2(new_n234), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n236), .B1(KEYINPUT4), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT5), .ZN(new_n242));
  NAND2_X1  g041(.A1(G225gat), .A2(G233gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n235), .B(KEYINPUT3), .Z(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n245), .B2(new_n222), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n221), .B(new_n235), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT5), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n240), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n251), .B1(new_n222), .B2(new_n235), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n252), .A2(new_n246), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n247), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G1gat), .B(G29gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT0), .ZN(new_n257));
  XOR2_X1   g056(.A(G57gat), .B(G85gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n255), .A2(KEYINPUT6), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n255), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(new_n260), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n255), .A2(new_n260), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT6), .B1(new_n255), .B2(new_n260), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n263), .A2(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  AOI21_X1  g067(.A(G190gat), .B1(new_n268), .B2(KEYINPUT27), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n269), .B(KEYINPUT28), .C1(KEYINPUT27), .C2(new_n268), .ZN(new_n270));
  AND2_X1   g069(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n271));
  NOR2_X1   g070(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n272));
  OAI21_X1  g071(.A(G183gat), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276));
  OAI211_X1 g075(.A(KEYINPUT69), .B(G183gat), .C1(new_n271), .C2(new_n272), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n269), .A4(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n269), .ZN(new_n281));
  OR2_X1    g080(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n268), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n281), .B1(new_n284), .B2(KEYINPUT69), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n276), .B1(new_n285), .B2(new_n275), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n270), .B1(new_n280), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G169gat), .ZN(new_n288));
  INV_X1    g087(.A(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT66), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT26), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT71), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n288), .A2(new_n289), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(KEYINPUT26), .B2(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n298), .A2(new_n302), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G190gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n268), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(KEYINPUT24), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(KEYINPUT67), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n306), .B(new_n307), .C1(new_n310), .C2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n290), .A2(new_n292), .A3(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT25), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(new_n301), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n313), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n319));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n320), .B1(KEYINPUT23), .B2(new_n299), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(KEYINPUT23), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT65), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n311), .ZN(new_n326));
  NAND4_X1  g125(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n325), .A2(new_n306), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n319), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n304), .A2(new_n334), .A3(new_n331), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n333), .A2(G226gat), .A3(G233gat), .A4(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT22), .ZN(new_n337));
  INV_X1    g136(.A(G211gat), .ZN(new_n338));
  INV_X1    g137(.A(G218gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G197gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT78), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G197gat), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n342), .A2(new_n344), .A3(G204gat), .ZN(new_n345));
  AOI21_X1  g144(.A(G204gat), .B1(new_n342), .B2(new_n344), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(G211gat), .B(G218gat), .Z(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n348), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n350), .B(new_n340), .C1(new_n345), .C2(new_n346), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n332), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n336), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AND4_X1   g159(.A1(G226gat), .A2(new_n304), .A3(G233gat), .A4(new_n331), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n333), .A2(new_n335), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n362), .B2(new_n358), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n360), .B1(new_n363), .B2(new_n357), .ZN(new_n364));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n360), .B(new_n367), .C1(new_n363), .C2(new_n357), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(KEYINPUT30), .A3(new_n370), .ZN(new_n371));
  OR3_X1    g170(.A1(new_n364), .A2(KEYINPUT30), .A3(new_n368), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n267), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n222), .B1(new_n304), .B2(new_n331), .ZN(new_n374));
  AOI211_X1 g173(.A(new_n221), .B(new_n330), .C1(new_n287), .C2(new_n303), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G227gat), .ZN(new_n377));
  INV_X1    g176(.A(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT34), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT34), .ZN(new_n381));
  OAI221_X1 g180(.A(new_n381), .B1(new_n377), .B2(new_n378), .C1(new_n374), .C2(new_n375), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT75), .B1(new_n376), .B2(new_n379), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n298), .A2(new_n302), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n308), .ZN(new_n387));
  INV_X1    g186(.A(new_n275), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n277), .A2(new_n269), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT70), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n279), .A3(new_n278), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n387), .B1(new_n391), .B2(new_n270), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n221), .B1(new_n392), .B2(new_n330), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n304), .A2(new_n222), .A3(new_n331), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n393), .A2(KEYINPUT75), .A3(new_n394), .A4(new_n379), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n384), .B1(new_n385), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT32), .B1(new_n385), .B2(new_n396), .ZN(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n397), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(KEYINPUT33), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT32), .B(new_n404), .C1(new_n385), .C2(new_n396), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n383), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n380), .A2(new_n382), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT32), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n379), .A3(new_n394), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n411), .B2(new_n395), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n407), .B1(new_n412), .B2(new_n404), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n406), .B1(new_n403), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n235), .A2(KEYINPUT3), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n354), .B(new_n355), .C1(KEYINPUT29), .C2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G228gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n378), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT29), .B1(new_n349), .B2(new_n351), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n235), .B1(new_n419), .B2(KEYINPUT3), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n237), .A2(new_n239), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(new_n419), .B2(KEYINPUT3), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT84), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n422), .B(new_n425), .C1(new_n419), .C2(KEYINPUT3), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n426), .A3(new_n416), .ZN(new_n427));
  INV_X1    g226(.A(new_n418), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n427), .A2(KEYINPUT85), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT85), .B1(new_n427), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n421), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(G22gat), .ZN(new_n432));
  INV_X1    g231(.A(G22gat), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n421), .C1(new_n429), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G78gat), .ZN(new_n436));
  INV_X1    g235(.A(G78gat), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n437), .A3(new_n434), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT31), .B(G50gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n439), .B(G106gat), .Z(new_n440));
  NAND3_X1  g239(.A1(new_n436), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n440), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n432), .A2(new_n437), .A3(new_n434), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n437), .B1(new_n432), .B2(new_n434), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n373), .A2(new_n414), .A3(new_n441), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT35), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n441), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT35), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n373), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT33), .B1(new_n411), .B2(new_n395), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n452), .A2(new_n412), .A3(new_n401), .ZN(new_n453));
  INV_X1    g252(.A(new_n405), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n407), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n405), .A2(new_n383), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT77), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n403), .A2(new_n413), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n447), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n363), .A2(new_n357), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n462), .A2(KEYINPUT88), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n357), .B1(new_n336), .B2(new_n359), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(KEYINPUT88), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n463), .B(KEYINPUT37), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n368), .B1(new_n364), .B2(KEYINPUT37), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(KEYINPUT38), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n364), .A2(KEYINPUT37), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT38), .B1(new_n470), .B2(new_n467), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(new_n267), .A3(new_n370), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n371), .A2(new_n372), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n255), .A2(new_n260), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n245), .A2(new_n222), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n243), .B1(new_n241), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT39), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n260), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT39), .B1(new_n248), .B2(new_n244), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(KEYINPUT87), .A2(KEYINPUT40), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n482), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n474), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n449), .A2(new_n472), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT36), .B1(new_n453), .B2(new_n456), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT76), .B1(new_n487), .B2(new_n406), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT36), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n403), .B2(new_n413), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT76), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n455), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n460), .A2(new_n489), .ZN(new_n494));
  INV_X1    g293(.A(new_n267), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n473), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n493), .A2(new_n494), .B1(new_n448), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n486), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n493), .A2(new_n494), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n448), .A2(new_n496), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n500), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n461), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT89), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g304(.A(KEYINPUT89), .B(new_n461), .C1(new_n499), .C2(new_n502), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n507), .A2(new_n508), .B1(G43gat), .B2(G50gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT95), .B(G50gat), .ZN(new_n510));
  OAI221_X1 g309(.A(new_n509), .B1(new_n507), .B2(new_n508), .C1(new_n510), .C2(G43gat), .ZN(new_n511));
  AND2_X1   g310(.A1(G43gat), .A2(G50gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(G43gat), .A2(G50gat), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT15), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G29gat), .A2(G36gat), .ZN(new_n515));
  OR3_X1    g314(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n511), .A2(new_n514), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT96), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(KEYINPUT93), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n517), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n516), .A2(KEYINPUT93), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n515), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n514), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT97), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT16), .ZN(new_n533));
  OR3_X1    g332(.A1(new_n533), .A2(KEYINPUT98), .A3(G1gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT98), .B1(new_n533), .B2(G1gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(KEYINPUT99), .ZN(new_n539));
  INV_X1    g338(.A(new_n538), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT99), .B1(new_n537), .B2(G1gat), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(G8gat), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT100), .B(G8gat), .Z(new_n543));
  OAI211_X1 g342(.A(new_n538), .B(new_n543), .C1(G1gat), .C2(new_n537), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT101), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n532), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT101), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n545), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n528), .A3(new_n531), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(KEYINPUT102), .A3(new_n550), .ZN(new_n551));
  OR3_X1    g350(.A1(new_n532), .A2(KEYINPUT102), .A3(new_n546), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n553), .B(KEYINPUT13), .Z(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n528), .A2(new_n556), .A3(new_n531), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n558));
  INV_X1    g357(.A(new_n545), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n553), .B(new_n550), .C1(new_n557), .C2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n559), .B(new_n558), .C1(new_n532), .C2(KEYINPUT17), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(KEYINPUT18), .A3(new_n553), .A4(new_n550), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n555), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT91), .ZN(new_n568));
  XOR2_X1   g367(.A(G113gat), .B(G141gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G169gat), .B(G197gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT92), .B(KEYINPUT12), .ZN(new_n573));
  XOR2_X1   g372(.A(new_n572), .B(new_n573), .Z(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n555), .A2(new_n563), .A3(new_n574), .A4(new_n565), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n505), .A2(new_n506), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT21), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581));
  INV_X1    g380(.A(G71gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n582), .B2(new_n437), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT103), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  XOR2_X1   g385(.A(G57gat), .B(G64gat), .Z(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G71gat), .B(G78gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n546), .B1(new_n580), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n590), .A2(KEYINPUT21), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT104), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n594), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n599), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT108), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(KEYINPUT108), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n613), .A2(KEYINPUT7), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  AOI22_X1  g415(.A1(KEYINPUT8), .A2(new_n616), .B1(new_n611), .B2(new_n612), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n615), .B(new_n617), .C1(KEYINPUT7), .C2(new_n613), .ZN(new_n618));
  XOR2_X1   g417(.A(G99gat), .B(G106gat), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT109), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n618), .A2(new_n619), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n532), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n625), .B(KEYINPUT107), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n558), .B(new_n623), .C1(new_n532), .C2(KEYINPUT17), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n632), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n629), .B2(new_n630), .ZN(new_n639));
  OR3_X1    g438(.A1(new_n633), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n637), .B1(new_n633), .B2(new_n639), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G120gat), .B(G148gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n644), .B(new_n645), .Z(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT110), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n623), .A2(new_n591), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n590), .A2(new_n622), .A3(new_n620), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n623), .A2(new_n651), .A3(new_n591), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n648), .B1(new_n650), .B2(new_n652), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n647), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n648), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n656), .A2(new_n647), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n609), .A2(new_n643), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n579), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n267), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g466(.A1(new_n579), .A2(new_n474), .A3(new_n663), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G8gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n664), .B2(new_n500), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n460), .A2(G15gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n664), .B2(new_n675), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n665), .A2(new_n448), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n642), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n505), .A2(new_n506), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n497), .A2(new_n486), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n461), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n643), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n680), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n608), .B(KEYINPUT113), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n578), .A2(KEYINPUT112), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n576), .A2(new_n690), .A3(new_n577), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n688), .A2(new_n662), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n682), .A2(new_n686), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G29gat), .B1(new_n694), .B2(new_n495), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n608), .A2(new_n642), .A3(new_n662), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n579), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n495), .A2(G29gat), .ZN(new_n698));
  OAI21_X1  g497(.A(KEYINPUT111), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT111), .ZN(new_n701));
  INV_X1    g500(.A(new_n698), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n579), .A2(new_n701), .A3(new_n696), .A4(new_n702), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n700), .B1(new_n699), .B2(new_n703), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n695), .B1(new_n704), .B2(new_n705), .ZN(G1328gat));
  OR2_X1    g505(.A1(new_n473), .A2(G36gat), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n697), .A2(KEYINPUT46), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G36gat), .B1(new_n694), .B2(new_n473), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT46), .B1(new_n697), .B2(new_n707), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(G1329gat));
  OAI21_X1  g510(.A(G43gat), .B1(new_n694), .B2(new_n500), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n460), .A2(G43gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n579), .A2(new_n696), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1330gat));
  OAI21_X1  g516(.A(new_n510), .B1(new_n694), .B2(new_n449), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n449), .A2(new_n510), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n579), .A2(new_n696), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT48), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1331gat));
  NAND4_X1  g522(.A1(new_n692), .A2(new_n608), .A3(new_n642), .A4(new_n662), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT114), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n684), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n267), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g528(.A1(new_n726), .A2(new_n473), .ZN(new_n730));
  NOR2_X1   g529(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n731));
  AND2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n730), .B2(new_n731), .ZN(G1333gat));
  OR3_X1    g533(.A1(new_n726), .A2(G71gat), .A3(new_n460), .ZN(new_n735));
  OAI21_X1  g534(.A(G71gat), .B1(new_n726), .B2(new_n500), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g537(.A1(new_n726), .A2(new_n449), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT115), .B(G78gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1335gat));
  INV_X1    g540(.A(new_n692), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n608), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n662), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n682), .A2(new_n686), .A3(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746), .B2(new_n495), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n684), .A2(new_n643), .A3(new_n743), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT51), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n267), .A2(new_n611), .A3(new_n662), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(G1336gat));
  NAND4_X1  g550(.A1(new_n682), .A2(new_n474), .A3(new_n686), .A4(new_n745), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G92gat), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n474), .A2(new_n612), .A3(new_n662), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n753), .B(new_n754), .C1(new_n749), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n748), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n748), .A2(new_n757), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n755), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(G92gat), .B2(new_n752), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n754), .B2(new_n761), .ZN(G1337gat));
  OAI21_X1  g561(.A(G99gat), .B1(new_n746), .B2(new_n500), .ZN(new_n763));
  INV_X1    g562(.A(new_n662), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n460), .A2(G99gat), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT117), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n763), .B1(new_n749), .B2(new_n766), .ZN(G1338gat));
  NAND4_X1  g566(.A1(new_n682), .A2(new_n448), .A3(new_n686), .A4(new_n745), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(G106gat), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770));
  OR3_X1    g569(.A1(new_n449), .A2(G106gat), .A3(new_n764), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n769), .B(new_n770), .C1(new_n749), .C2(new_n771), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n768), .A2(KEYINPUT118), .A3(G106gat), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT118), .B1(new_n768), .B2(G106gat), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n771), .B1(new_n758), .B2(new_n759), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n776), .B2(new_n770), .ZN(G1339gat));
  INV_X1    g576(.A(new_n649), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n659), .B(KEYINPUT54), .C1(new_n778), .C2(new_n658), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n646), .B1(new_n655), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(KEYINPUT119), .A3(new_n661), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT55), .B1(new_n779), .B2(new_n781), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT119), .B1(new_n782), .B2(new_n661), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n689), .A3(new_n691), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n554), .B1(new_n551), .B2(new_n552), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n553), .B1(new_n564), .B2(new_n550), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n572), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n577), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n662), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n643), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n643), .A2(new_n787), .A3(new_n792), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n687), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n663), .A2(new_n692), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n495), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n449), .A2(new_n414), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n473), .ZN(new_n802));
  AOI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n742), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n448), .B1(new_n797), .B2(new_n798), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n460), .A2(new_n474), .A3(new_n495), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n209), .B1(new_n576), .B2(new_n577), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(G1340gat));
  NAND3_X1  g608(.A1(new_n802), .A2(new_n214), .A3(new_n662), .ZN(new_n810));
  OAI21_X1  g609(.A(G120gat), .B1(new_n806), .B2(new_n764), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(G1341gat));
  INV_X1    g611(.A(G127gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n802), .A2(new_n813), .A3(new_n608), .ZN(new_n814));
  OAI21_X1  g613(.A(G127gat), .B1(new_n806), .B2(new_n687), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1342gat));
  INV_X1    g615(.A(G134gat), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n642), .A2(new_n474), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n819), .A2(KEYINPUT56), .ZN(new_n820));
  OAI21_X1  g619(.A(G134gat), .B1(new_n806), .B2(new_n642), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(KEYINPUT56), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(G1343gat));
  AOI21_X1  g622(.A(new_n449), .B1(new_n797), .B2(new_n798), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n782), .A2(new_n661), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n779), .A2(new_n781), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n578), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n643), .B1(new_n793), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n609), .B1(new_n796), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n798), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n448), .A2(KEYINPUT57), .ZN(new_n833));
  OAI22_X1  g632(.A1(new_n824), .A2(KEYINPUT57), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n500), .A2(new_n267), .A3(new_n473), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n578), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT121), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n834), .A2(new_n839), .A3(new_n578), .A4(new_n836), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n840), .A3(G141gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n799), .A2(new_n448), .A3(new_n500), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n474), .ZN(new_n843));
  AOI21_X1  g642(.A(G141gat), .B1(new_n576), .B2(new_n577), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT58), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n834), .A2(new_n836), .ZN(new_n847));
  OAI21_X1  g646(.A(G141gat), .B1(new_n847), .B2(new_n692), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n844), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT58), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n846), .A2(new_n851), .ZN(G1344gat));
  INV_X1    g651(.A(new_n663), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n831), .B1(new_n578), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT57), .B1(new_n854), .B2(new_n448), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n833), .B1(new_n797), .B2(new_n798), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n662), .A3(new_n836), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n859));
  INV_X1    g658(.A(new_n847), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n662), .ZN(new_n862));
  INV_X1    g661(.A(new_n230), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n861), .B1(new_n843), .B2(new_n662), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n859), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(G1345gat));
  AOI21_X1  g664(.A(G155gat), .B1(new_n843), .B2(new_n608), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n688), .A2(G155gat), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT122), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n860), .B2(new_n868), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n847), .B2(new_n642), .ZN(new_n870));
  INV_X1    g669(.A(G162gat), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n818), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n870), .B1(new_n842), .B2(new_n872), .ZN(G1347gat));
  NAND2_X1  g672(.A1(new_n797), .A2(new_n798), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n473), .A2(new_n267), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n800), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(G169gat), .B1(new_n878), .B2(new_n742), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n460), .A2(new_n267), .A3(new_n473), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n804), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n288), .B1(new_n576), .B2(new_n577), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(G1348gat));
  NOR3_X1   g682(.A1(new_n877), .A2(G176gat), .A3(new_n764), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n662), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(G176gat), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT123), .Z(G1349gat));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT60), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(KEYINPUT60), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n881), .A2(new_n688), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G183gat), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT27), .B(G183gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n608), .A3(new_n893), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n889), .B(new_n890), .C1(new_n892), .C2(new_n894), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n888), .A2(new_n892), .A3(KEYINPUT60), .A4(new_n894), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(G1350gat));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n305), .A3(new_n643), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n643), .ZN(new_n899));
  NOR2_X1   g698(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n305), .B1(KEYINPUT125), .B2(KEYINPUT61), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n898), .B1(new_n902), .B2(new_n903), .ZN(G1351gat));
  AND2_X1   g703(.A1(new_n500), .A2(new_n875), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n824), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(G197gat), .B1(new_n907), .B2(new_n742), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n857), .A2(new_n905), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n341), .B1(new_n576), .B2(new_n577), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1352gat));
  NOR2_X1   g711(.A1(new_n764), .A2(G204gat), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n874), .A2(new_n448), .A3(new_n905), .A4(new_n913), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT126), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(KEYINPUT126), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT127), .B1(new_n917), .B2(KEYINPUT62), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n915), .A2(new_n919), .A3(new_n920), .A4(new_n916), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n857), .A2(new_n662), .A3(new_n905), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n923), .A2(G204gat), .B1(new_n917), .B2(KEYINPUT62), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n338), .A3(new_n608), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n608), .B(new_n905), .C1(new_n855), .C2(new_n856), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n909), .B2(new_n642), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n907), .A2(new_n339), .A3(new_n643), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1355gat));
endmodule


