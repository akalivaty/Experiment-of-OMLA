//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT67), .B(G128), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(G143), .B2(new_n192), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n193), .A2(new_n195), .A3(new_n198), .A4(G128), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT65), .A2(G137), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT65), .A2(G137), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n207), .B2(G134), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n202), .B1(G131), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT11), .B1(new_n203), .B2(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n204), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT11), .A2(G134), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT66), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  NOR4_X1   g030(.A1(new_n205), .A2(new_n206), .A3(new_n213), .A4(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n210), .B(new_n212), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n209), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n212), .B1(new_n215), .B2(new_n217), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(new_n218), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n193), .A2(new_n195), .A3(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n193), .A2(new_n195), .ZN(new_n226));
  XOR2_X1   g040(.A(KEYINPUT0), .B(G128), .Z(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n220), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n228), .ZN(new_n230));
  AOI211_X1 g044(.A(KEYINPUT68), .B(new_n230), .C1(new_n222), .C2(new_n218), .ZN(new_n231));
  OAI211_X1 g045(.A(KEYINPUT30), .B(new_n219), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT30), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n228), .B(KEYINPUT64), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n219), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n232), .A2(new_n237), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n246), .B(new_n219), .C1(new_n229), .C2(new_n231), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n191), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n244), .B1(new_n235), .B2(new_n236), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n236), .A2(new_n244), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n223), .A2(new_n228), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT28), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  AOI211_X1 g069(.A(KEYINPUT29), .B(new_n248), .C1(new_n191), .C2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n219), .B1(new_n229), .B2(new_n231), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n244), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n249), .B1(new_n258), .B2(new_n247), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n254), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT29), .A3(new_n191), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(G472), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n247), .A2(new_n191), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n247), .A2(KEYINPUT69), .A3(new_n191), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n268), .A2(new_n269), .A3(new_n245), .A4(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT31), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n245), .A2(new_n270), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n274), .A2(new_n269), .A3(KEYINPUT31), .A4(new_n268), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n255), .A2(new_n191), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(G902), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G472), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n265), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n273), .B2(new_n275), .ZN(new_n282));
  NOR4_X1   g096(.A1(new_n282), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n264), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(G234), .B2(new_n262), .ZN(new_n286));
  INV_X1    g100(.A(G110), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G110), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n291), .B1(new_n288), .B2(new_n290), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G128), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n296), .A2(G119), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n197), .B2(G119), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT23), .B1(new_n296), .B2(G119), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n238), .B2(G128), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(KEYINPUT67), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G128), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT23), .A4(G119), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT74), .B(G110), .Z(new_n307));
  AOI22_X1  g121(.A1(new_n295), .A2(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT72), .A3(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(G125), .ZN(new_n311));
  INV_X1    g125(.A(G125), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(KEYINPUT16), .B(new_n310), .C1(new_n314), .C2(KEYINPUT72), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT16), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n192), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n314), .A2(G146), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n308), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n317), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n192), .A3(new_n317), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n301), .A2(new_n305), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n294), .A2(new_n298), .B1(new_n326), .B2(G110), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n321), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n315), .A2(new_n192), .A3(new_n317), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n327), .B(new_n321), .C1(new_n329), .C2(new_n318), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n320), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n308), .A2(new_n318), .A3(new_n319), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n327), .B1(new_n329), .B2(new_n318), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT73), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G137), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(G221), .A3(G234), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n340), .B(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n332), .A2(KEYINPUT75), .A3(new_n343), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT25), .B1(new_n346), .B2(new_n262), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n348));
  AOI211_X1 g162(.A(new_n348), .B(G902), .C1(new_n344), .C2(new_n345), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n286), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n286), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n343), .B1(new_n337), .B2(new_n338), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n332), .A2(KEYINPUT75), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n332), .A2(KEYINPUT75), .A3(new_n343), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n262), .B(new_n351), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT76), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n346), .A2(new_n358), .A3(new_n262), .A4(new_n351), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n350), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT3), .B1(new_n362), .B2(G107), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n364));
  INV_X1    g178(.A(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(G104), .ZN(new_n366));
  INV_X1    g180(.A(G101), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(G107), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n366), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n362), .A2(G107), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n365), .A2(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(G101), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n373), .A2(G128), .B1(new_n193), .B2(new_n195), .ZN(new_n374));
  INV_X1    g188(.A(new_n201), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n369), .B(new_n372), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n369), .A2(new_n372), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n200), .A3(new_n201), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n223), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT12), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(KEYINPUT80), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n222), .A2(new_n218), .B1(new_n376), .B2(new_n378), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(KEYINPUT12), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(KEYINPUT12), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(G110), .B(G140), .ZN(new_n388));
  INV_X1    g202(.A(G227), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G953), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n388), .B(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n363), .A2(new_n366), .A3(new_n368), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(G101), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n228), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(G101), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n369), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n369), .A2(KEYINPUT4), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT78), .A3(new_n396), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n395), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT10), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n376), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n377), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n200), .A2(new_n201), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT10), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n223), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n391), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n387), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n397), .A2(new_n398), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT78), .B1(new_n400), .B2(new_n396), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n228), .B(new_n394), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n410), .A3(new_n404), .A4(new_n407), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n223), .B1(new_n402), .B2(new_n408), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n391), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G469), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n387), .A2(new_n416), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n391), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n411), .A2(new_n417), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(G469), .A3(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n421), .A2(new_n262), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT9), .B(G234), .ZN(new_n430));
  OAI21_X1  g244(.A(G221), .B1(new_n430), .B2(G902), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT77), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT81), .Z(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT82), .ZN(new_n437));
  OAI21_X1  g251(.A(G210), .B1(G237), .B2(G902), .ZN(new_n438));
  XNOR2_X1  g252(.A(G116), .B(G119), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT5), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT84), .ZN(new_n441));
  INV_X1    g255(.A(G113), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n240), .A2(G119), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT5), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT84), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n439), .A2(new_n446), .A3(KEYINPUT5), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n441), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n242), .A2(new_n243), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n377), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n440), .A2(new_n445), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT83), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT83), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n440), .A2(new_n455), .A3(new_n445), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n454), .A2(new_n449), .A3(new_n377), .A4(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n458), .B(KEYINPUT8), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n451), .A2(new_n452), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n459), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT85), .B1(new_n461), .B2(new_n450), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G224), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(new_n464), .B2(G953), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(G125), .B(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT86), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n200), .A2(new_n312), .A3(new_n201), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n202), .A2(KEYINPUT86), .A3(new_n312), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n469), .A2(new_n467), .ZN(new_n473));
  OAI22_X1  g287(.A1(new_n472), .A2(KEYINPUT87), .B1(new_n473), .B2(new_n465), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n472), .A2(KEYINPUT87), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n463), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n244), .B(new_n394), .C1(new_n413), .C2(new_n414), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n454), .A2(new_n449), .A3(new_n456), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n477), .B(new_n458), .C1(new_n377), .C2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(G902), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n458), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n244), .A2(new_n394), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n399), .B2(new_n401), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n478), .A2(new_n377), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n479), .A2(new_n485), .A3(KEYINPUT6), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n487), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n464), .A2(G953), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n473), .B(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n438), .B1(new_n480), .B2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n460), .A2(new_n462), .ZN(new_n493));
  INV_X1    g307(.A(new_n475), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n473), .A2(new_n465), .ZN(new_n495));
  INV_X1    g309(.A(new_n472), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT87), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n493), .A2(new_n494), .A3(new_n479), .A4(new_n498), .ZN(new_n499));
  AND4_X1   g313(.A1(new_n262), .A2(new_n491), .A3(new_n499), .A4(new_n438), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n437), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G122), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT90), .B1(new_n502), .B2(G116), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n240), .A3(G122), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(G116), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n365), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n197), .A2(G143), .ZN(new_n509));
  INV_X1    g323(.A(G134), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n296), .A2(G143), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n510), .B1(new_n509), .B2(new_n512), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n508), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n506), .A2(KEYINPUT14), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n506), .A2(KEYINPUT14), .B1(G116), .B2(new_n502), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n365), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n508), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n365), .B1(new_n506), .B2(new_n507), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n513), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT13), .B1(new_n194), .B2(G128), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n197), .A2(G143), .B1(KEYINPUT13), .B2(new_n511), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n510), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI22_X1  g341(.A1(new_n516), .A2(new_n519), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n430), .A2(new_n285), .A3(G953), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT92), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n517), .A2(new_n518), .ZN(new_n532));
  OAI221_X1 g346(.A(new_n508), .B1(new_n514), .B2(new_n515), .C1(new_n532), .C2(new_n365), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n522), .A2(new_n527), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT92), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .A4(new_n529), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n528), .A2(new_n530), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G478), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n262), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n538), .B2(new_n262), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT88), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n548), .A2(new_n549), .A3(G131), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n187), .A2(G214), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n194), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n210), .B1(new_n552), .B2(new_n547), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n546), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT19), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n311), .A2(new_n313), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n310), .B1(new_n314), .B2(KEYINPUT72), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n192), .B(new_n556), .C1(new_n557), .C2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(G131), .B1(new_n548), .B2(new_n549), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n210), .A3(new_n547), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT88), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n554), .A2(new_n323), .A3(new_n558), .A4(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n552), .B(new_n547), .C1(new_n563), .C2(new_n210), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n557), .A2(new_n192), .ZN(new_n565));
  OAI221_X1 g379(.A(new_n564), .B1(new_n559), .B2(new_n563), .C1(new_n565), .C2(new_n319), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G113), .B(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n362), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n553), .A2(KEYINPUT17), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT17), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n559), .A2(new_n560), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n323), .A2(new_n324), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n566), .A3(new_n569), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT89), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT20), .ZN(new_n581));
  INV_X1    g395(.A(new_n578), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n571), .B2(new_n576), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n584));
  OAI21_X1  g398(.A(KEYINPUT89), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n575), .A2(new_n566), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n570), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n576), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n262), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G475), .ZN(new_n592));
  NAND2_X1  g406(.A1(G234), .A2(G237), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(G952), .A3(new_n341), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(G902), .A3(G953), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT21), .B(G898), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n545), .A2(new_n587), .A3(new_n592), .A4(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n434), .A2(new_n501), .A3(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n284), .A2(new_n361), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n279), .A2(new_n280), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n282), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n427), .B1(new_n420), .B2(new_n421), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n432), .B1(new_n609), .B2(new_n426), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n350), .A2(new_n360), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n533), .A2(new_n534), .A3(new_n529), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n537), .A3(KEYINPUT33), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n614), .A2(KEYINPUT93), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n538), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(KEYINPUT93), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n539), .A2(G902), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n615), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n538), .A2(new_n262), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n620), .B1(G478), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n587), .A2(new_n592), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n491), .A2(new_n499), .A3(new_n262), .ZN(new_n625));
  INV_X1    g439(.A(new_n438), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n491), .A2(new_n499), .A3(new_n262), .A4(new_n438), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n436), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n600), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n612), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT34), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  INV_X1    g447(.A(KEYINPUT95), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n545), .B1(G475), .B2(new_n591), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n581), .A2(new_n585), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT94), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n581), .A2(new_n585), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n586), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n634), .B1(new_n641), .B2(new_n630), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n635), .A2(new_n640), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n436), .B(new_n599), .C1(new_n627), .C2(new_n628), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(KEYINPUT95), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n612), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT96), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT97), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT36), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n343), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n337), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n262), .A3(new_n351), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n350), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n605), .A2(new_n602), .A3(new_n606), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT98), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT37), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  XNOR2_X1  g473(.A(KEYINPUT99), .B(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n595), .B1(new_n660), .B2(new_n597), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n641), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n655), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n284), .A2(new_n610), .A3(new_n629), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT100), .B(G128), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G30));
  NAND2_X1  g480(.A1(new_n274), .A2(new_n268), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n258), .A2(new_n247), .ZN(new_n668));
  INV_X1    g482(.A(new_n191), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n667), .A2(KEYINPUT101), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n262), .ZN(new_n672));
  AOI21_X1  g486(.A(KEYINPUT101), .B1(new_n667), .B2(new_n670), .ZN(new_n673));
  OAI21_X1  g487(.A(G472), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n281), .B2(new_n283), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n675), .B(KEYINPUT102), .Z(new_n676));
  XOR2_X1   g490(.A(new_n661), .B(KEYINPUT39), .Z(new_n677));
  NAND2_X1  g491(.A1(new_n610), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT40), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n627), .A2(new_n628), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT38), .Z(new_n681));
  INV_X1    g495(.A(new_n545), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n623), .ZN(new_n683));
  OR3_X1    g497(.A1(new_n655), .A2(new_n436), .A3(new_n683), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n676), .A2(new_n679), .A3(new_n681), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n194), .ZN(G45));
  INV_X1    g500(.A(new_n655), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n624), .A2(new_n661), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n284), .A2(new_n610), .A3(new_n629), .A4(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT103), .B(G146), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G48));
  NAND2_X1  g507(.A1(new_n284), .A2(new_n361), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n387), .A2(new_n411), .B1(new_n418), .B2(new_n391), .ZN(new_n696));
  OAI21_X1  g510(.A(G469), .B1(new_n696), .B2(G902), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n422), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n431), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n630), .A2(new_n699), .A3(new_n624), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  AOI21_X1  g517(.A(new_n699), .B1(new_n645), .B2(new_n642), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n695), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  NOR3_X1   g520(.A1(new_n687), .A2(new_n601), .A3(new_n699), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n284), .A2(new_n629), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  INV_X1    g523(.A(new_n436), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n680), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n422), .A2(new_n697), .A3(new_n431), .A4(new_n600), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n683), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n669), .B1(new_n259), .B2(new_n254), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n276), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(G472), .A2(G902), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n713), .A2(new_n361), .A3(new_n606), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NAND4_X1  g533(.A1(new_n606), .A2(new_n717), .A3(new_n655), .A4(new_n688), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n629), .A2(new_n698), .A3(new_n431), .ZN(new_n721));
  OR3_X1    g535(.A1(new_n720), .A2(KEYINPUT104), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT104), .B1(new_n720), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  OR3_X1    g539(.A1(new_n680), .A2(KEYINPUT106), .A3(new_n436), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n426), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n426), .A2(new_n727), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n609), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT106), .B1(new_n680), .B2(new_n436), .ZN(new_n731));
  AND4_X1   g545(.A1(new_n431), .A2(new_n726), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n284), .A2(new_n361), .A3(new_n688), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT107), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n733), .A2(new_n734), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n733), .A2(new_n734), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND4_X1  g557(.A1(new_n284), .A2(new_n361), .A3(new_n662), .A4(new_n732), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  AND2_X1   g559(.A1(new_n587), .A2(new_n592), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n622), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n747), .B1(new_n748), .B2(KEYINPUT43), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n748), .A2(KEYINPUT43), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n608), .A3(new_n687), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT44), .Z(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n424), .A2(new_n425), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT45), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n756), .A2(G469), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n754), .B1(new_n757), .B2(new_n427), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n757), .A2(new_n754), .A3(new_n427), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n422), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n431), .B(new_n677), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n726), .A2(new_n731), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n753), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  OAI21_X1  g581(.A(new_n431), .B1(new_n761), .B2(new_n762), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OR4_X1    g586(.A1(new_n284), .A2(new_n361), .A3(new_n689), .A4(new_n764), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  NOR3_X1   g590(.A1(new_n655), .A2(KEYINPUT112), .A3(new_n661), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n629), .A2(new_n623), .A3(new_n682), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n730), .A2(new_n431), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(KEYINPUT112), .B1(new_n655), .B2(new_n661), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n675), .A3(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n724), .A2(new_n782), .A3(new_n664), .A4(new_n691), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT113), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n788));
  INV_X1    g602(.A(new_n661), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n545), .A2(new_n592), .A3(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n640), .A3(KEYINPUT110), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT110), .B1(new_n790), .B2(new_n640), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n655), .A2(new_n610), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n606), .A2(new_n717), .A3(new_n655), .A4(new_n688), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n730), .A2(new_n431), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n284), .A2(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n744), .B1(new_n798), .B2(new_n764), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n284), .B(new_n361), .C1(new_n704), .C2(new_n700), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n437), .B(new_n600), .C1(new_n492), .C2(new_n500), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n746), .A2(new_n682), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n801), .B1(new_n624), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n605), .A2(new_n611), .A3(new_n803), .A4(new_n606), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n804), .A2(new_n656), .A3(new_n718), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n800), .A2(new_n805), .A3(new_n603), .A4(new_n708), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n799), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n737), .A3(new_n741), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n737), .A3(new_n741), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT111), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n787), .A2(new_n788), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n783), .B(new_n784), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(KEYINPUT53), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n815), .A3(KEYINPUT54), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n814), .A2(new_n788), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT53), .B1(new_n735), .B2(new_n736), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n806), .A3(new_n799), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n787), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n817), .A2(new_n820), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n751), .A2(new_n594), .ZN(new_n828));
  INV_X1    g642(.A(new_n431), .ZN(new_n829));
  INV_X1    g643(.A(new_n698), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n764), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n695), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n833), .B(KEYINPUT48), .Z(new_n834));
  NAND4_X1  g648(.A1(new_n676), .A2(new_n361), .A3(new_n595), .A4(new_n831), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n835), .A2(new_n624), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n606), .A2(new_n717), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n828), .A2(new_n361), .A3(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(G952), .B(new_n341), .C1(new_n838), .C2(new_n721), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n834), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(KEYINPUT116), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n770), .B(new_n771), .C1(new_n433), .C2(new_n830), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n838), .A2(new_n764), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n837), .A2(new_n655), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n842), .A2(new_n843), .B1(new_n844), .B2(new_n832), .ZN(new_n845));
  OR3_X1    g659(.A1(new_n835), .A2(new_n623), .A3(new_n622), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n681), .A2(new_n431), .A3(new_n436), .A4(new_n698), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT115), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT50), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT51), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n841), .A2(new_n851), .ZN(new_n852));
  OAI22_X1  g666(.A1(new_n827), .A2(new_n852), .B1(G952), .B2(G953), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n698), .B(KEYINPUT49), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n433), .A2(new_n854), .A3(new_n437), .A4(new_n747), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n676), .A2(new_n361), .A3(new_n681), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n856), .ZN(G75));
  NOR2_X1   g671(.A1(new_n341), .A2(G952), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n814), .A2(new_n788), .B1(new_n787), .B2(new_n824), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n262), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT56), .B1(new_n861), .B2(G210), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n486), .A2(new_n488), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(new_n490), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT55), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n859), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n862), .B2(new_n865), .ZN(G51));
  INV_X1    g681(.A(new_n696), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n860), .A2(KEYINPUT117), .A3(new_n822), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n821), .A2(new_n825), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n826), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n427), .B(KEYINPUT57), .Z(new_n875));
  OAI21_X1  g689(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n861), .A2(new_n757), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n858), .B1(new_n876), .B2(new_n877), .ZN(G54));
  NAND2_X1  g692(.A1(KEYINPUT58), .A2(G475), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT118), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n879), .A2(KEYINPUT118), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n861), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n577), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n858), .ZN(G60));
  AND3_X1   g700(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n887));
  NAND2_X1  g701(.A1(G478), .A2(G902), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT59), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n827), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n889), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n873), .A2(new_n871), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n870), .A2(new_n872), .A3(KEYINPUT54), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n891), .B1(new_n895), .B2(new_n858), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT119), .B(new_n859), .C1(new_n874), .C2(new_n892), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n890), .B1(new_n896), .B2(new_n897), .ZN(G63));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n901));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT60), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n821), .B2(new_n825), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT120), .B1(new_n905), .B2(new_n653), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n907));
  INV_X1    g721(.A(new_n653), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n860), .A2(new_n907), .A3(new_n908), .A4(new_n904), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n859), .B1(new_n905), .B2(new_n346), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n900), .B(new_n901), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n870), .A2(new_n903), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n907), .B1(new_n913), .B2(new_n908), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n905), .A2(KEYINPUT120), .A3(new_n653), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n911), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(KEYINPUT121), .A3(new_n899), .A4(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n912), .A2(new_n918), .ZN(G66));
  NAND2_X1  g733(.A1(new_n806), .A2(new_n341), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(KEYINPUT122), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n598), .B2(new_n464), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n863), .B1(G898), .B2(new_n341), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(G69));
  AOI21_X1  g740(.A(new_n341), .B1(G227), .B2(G900), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT125), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n232), .A2(new_n237), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n556), .B1(new_n557), .B2(new_n555), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n802), .A2(new_n624), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OR4_X1    g751(.A1(new_n694), .A2(new_n678), .A3(new_n764), .A4(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n775), .A2(new_n766), .A3(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n940));
  AND2_X1   g754(.A1(new_n664), .A2(new_n691), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n724), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n685), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n685), .A2(new_n942), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n944), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n939), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n935), .B1(new_n946), .B2(G953), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT124), .B(new_n935), .C1(new_n946), .C2(G953), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR3_X1    g765(.A1(new_n763), .A2(new_n694), .A3(new_n778), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n775), .A2(new_n766), .A3(new_n744), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n942), .ZN(new_n954));
  AOI21_X1  g768(.A(G953), .B1(new_n954), .B2(new_n742), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n341), .A2(G900), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n934), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n930), .B(new_n931), .C1(new_n951), .C2(new_n957), .ZN(new_n958));
  AND4_X1   g772(.A1(KEYINPUT126), .A2(new_n951), .A3(new_n957), .A4(new_n929), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(G72));
  NAND2_X1  g774(.A1(new_n245), .A2(new_n247), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n191), .ZN(new_n962));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT63), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n858), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n954), .A2(new_n742), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n191), .A3(new_n961), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n946), .A2(new_n191), .A3(new_n961), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n969), .B2(new_n806), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n248), .B(KEYINPUT127), .Z(new_n971));
  AOI21_X1  g785(.A(new_n964), .B1(new_n971), .B2(new_n667), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n816), .B2(new_n972), .ZN(G57));
endmodule


