

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(KEYINPUT31), .ZN(n740) );
  XOR2_X1 U554 ( .A(KEYINPUT100), .B(n701), .Z(n774) );
  XNOR2_X1 U555 ( .A(G2104), .B(KEYINPUT65), .ZN(n523) );
  XOR2_X1 U556 ( .A(KEYINPUT32), .B(n751), .Z(n521) );
  OR2_X1 U557 ( .A1(n755), .A2(n734), .ZN(n735) );
  INV_X1 U558 ( .A(n703), .ZN(n717) );
  INV_X1 U559 ( .A(n717), .ZN(n744) );
  XNOR2_X1 U560 ( .A(n741), .B(n740), .ZN(n742) );
  AND2_X1 U561 ( .A1(n774), .A2(n732), .ZN(n755) );
  INV_X1 U562 ( .A(n784), .ZN(n700) );
  NAND2_X1 U563 ( .A1(n783), .A2(n700), .ZN(n703) );
  NAND2_X1 U564 ( .A1(n703), .A2(G8), .ZN(n701) );
  NOR2_X1 U565 ( .A1(G164), .A2(G1384), .ZN(n699) );
  NOR2_X1 U566 ( .A1(n648), .A2(G651), .ZN(n659) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  NOR2_X1 U568 ( .A1(n529), .A2(n528), .ZN(G164) );
  XOR2_X2 U569 ( .A(KEYINPUT17), .B(n522), .Z(n893) );
  AND2_X1 U570 ( .A1(G138), .A2(n893), .ZN(n529) );
  AND2_X1 U571 ( .A1(n523), .A2(G2105), .ZN(n898) );
  NAND2_X1 U572 ( .A1(G126), .A2(n898), .ZN(n527) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n896) );
  NAND2_X1 U574 ( .A1(G114), .A2(n896), .ZN(n525) );
  NOR2_X2 U575 ( .A1(G2105), .A2(n523), .ZN(n545) );
  NAND2_X1 U576 ( .A1(G102), .A2(n545), .ZN(n524) );
  AND2_X1 U577 ( .A1(n525), .A2(n524), .ZN(n526) );
  NAND2_X1 U578 ( .A1(n527), .A2(n526), .ZN(n528) );
  INV_X1 U579 ( .A(G651), .ZN(n536) );
  NOR2_X1 U580 ( .A1(G543), .A2(n536), .ZN(n530) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n530), .Z(n663) );
  NAND2_X1 U582 ( .A1(G63), .A2(n663), .ZN(n533) );
  XNOR2_X1 U583 ( .A(G543), .B(KEYINPUT0), .ZN(n531) );
  XNOR2_X1 U584 ( .A(n531), .B(KEYINPUT67), .ZN(n648) );
  NAND2_X1 U585 ( .A1(G51), .A2(n659), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U587 ( .A(KEYINPUT6), .B(n534), .ZN(n542) );
  NOR2_X1 U588 ( .A1(G543), .A2(G651), .ZN(n655) );
  NAND2_X1 U589 ( .A1(n655), .A2(G89), .ZN(n535) );
  XNOR2_X1 U590 ( .A(n535), .B(KEYINPUT4), .ZN(n538) );
  NOR2_X1 U591 ( .A1(n648), .A2(n536), .ZN(n654) );
  NAND2_X1 U592 ( .A1(G76), .A2(n654), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U594 ( .A(KEYINPUT74), .B(n539), .Z(n540) );
  XNOR2_X1 U595 ( .A(KEYINPUT5), .B(n540), .ZN(n541) );
  NOR2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U597 ( .A(KEYINPUT7), .B(n543), .Z(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U599 ( .A1(G125), .A2(n898), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n544), .B(KEYINPUT66), .ZN(n548) );
  NAND2_X1 U601 ( .A1(G101), .A2(n545), .ZN(n546) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(n546), .Z(n547) );
  NAND2_X1 U603 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n896), .A2(G113), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n893), .A2(G137), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n552), .A2(n551), .ZN(G160) );
  XOR2_X1 U608 ( .A(G2438), .B(G2454), .Z(n554) );
  XNOR2_X1 U609 ( .A(G2435), .B(G2430), .ZN(n553) );
  XNOR2_X1 U610 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U611 ( .A(n555), .B(KEYINPUT108), .Z(n557) );
  XNOR2_X1 U612 ( .A(G1341), .B(G1348), .ZN(n556) );
  XNOR2_X1 U613 ( .A(n557), .B(n556), .ZN(n561) );
  XOR2_X1 U614 ( .A(G2427), .B(G2443), .Z(n559) );
  XNOR2_X1 U615 ( .A(G2451), .B(G2446), .ZN(n558) );
  XNOR2_X1 U616 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U617 ( .A(n561), .B(n560), .Z(n562) );
  AND2_X1 U618 ( .A1(G14), .A2(n562), .ZN(G401) );
  NAND2_X1 U619 ( .A1(G64), .A2(n663), .ZN(n564) );
  NAND2_X1 U620 ( .A1(G52), .A2(n659), .ZN(n563) );
  NAND2_X1 U621 ( .A1(n564), .A2(n563), .ZN(n569) );
  NAND2_X1 U622 ( .A1(G77), .A2(n654), .ZN(n566) );
  NAND2_X1 U623 ( .A1(G90), .A2(n655), .ZN(n565) );
  NAND2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n567), .Z(n568) );
  NOR2_X1 U626 ( .A1(n569), .A2(n568), .ZN(G171) );
  AND2_X1 U627 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U628 ( .A(G132), .ZN(G219) );
  INV_X1 U629 ( .A(G82), .ZN(G220) );
  INV_X1 U630 ( .A(G57), .ZN(G237) );
  INV_X1 U631 ( .A(G120), .ZN(G236) );
  NAND2_X1 U632 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U633 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U634 ( .A(G223), .B(KEYINPUT70), .Z(n834) );
  NAND2_X1 U635 ( .A1(n834), .A2(G567), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT71), .ZN(n572) );
  XNOR2_X1 U637 ( .A(KEYINPUT11), .B(n572), .ZN(G234) );
  NAND2_X1 U638 ( .A1(G56), .A2(n663), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n573), .Z(n579) );
  NAND2_X1 U640 ( .A1(n655), .A2(G81), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G68), .A2(n654), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT13), .B(n577), .Z(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n659), .A2(G43), .ZN(n580) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n998) );
  INV_X1 U648 ( .A(G860), .ZN(n603) );
  OR2_X1 U649 ( .A1(n998), .A2(n603), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U652 ( .A1(G54), .A2(n659), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G79), .A2(n654), .ZN(n583) );
  NAND2_X1 U654 ( .A1(G66), .A2(n663), .ZN(n582) );
  NAND2_X1 U655 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n655), .A2(G92), .ZN(n584) );
  XOR2_X1 U657 ( .A(KEYINPUT72), .B(n584), .Z(n585) );
  NOR2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT15), .ZN(n590) );
  XNOR2_X1 U661 ( .A(KEYINPUT73), .B(n590), .ZN(n1004) );
  INV_X1 U662 ( .A(G868), .ZN(n676) );
  NAND2_X1 U663 ( .A1(n1004), .A2(n676), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(G284) );
  NOR2_X1 U665 ( .A1(G286), .A2(n676), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT75), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G65), .A2(n663), .ZN(n595) );
  NAND2_X1 U668 ( .A1(G53), .A2(n659), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U670 ( .A1(G78), .A2(n654), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G91), .A2(n655), .ZN(n596) );
  NAND2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U673 ( .A1(n599), .A2(n598), .ZN(n917) );
  NAND2_X1 U674 ( .A1(n917), .A2(n676), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT76), .B(n602), .Z(G297) );
  NAND2_X1 U677 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U678 ( .A(n1004), .ZN(n841) );
  NAND2_X1 U679 ( .A1(n604), .A2(n841), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT16), .ZN(n606) );
  XOR2_X1 U681 ( .A(KEYINPUT77), .B(n606), .Z(G148) );
  NAND2_X1 U682 ( .A1(n841), .A2(G868), .ZN(n607) );
  NOR2_X1 U683 ( .A1(G559), .A2(n607), .ZN(n608) );
  XOR2_X1 U684 ( .A(KEYINPUT79), .B(n608), .Z(n611) );
  NOR2_X1 U685 ( .A1(G868), .A2(n998), .ZN(n609) );
  XNOR2_X1 U686 ( .A(KEYINPUT78), .B(n609), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U688 ( .A1(n898), .A2(G123), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G111), .A2(n896), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U692 ( .A1(G135), .A2(n893), .ZN(n616) );
  NAND2_X1 U693 ( .A1(G99), .A2(n545), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n979) );
  XOR2_X1 U696 ( .A(G2096), .B(n979), .Z(n619) );
  NOR2_X1 U697 ( .A1(G2100), .A2(n619), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT80), .B(n620), .Z(G156) );
  NAND2_X1 U699 ( .A1(G80), .A2(n654), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G93), .A2(n655), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n663), .A2(G67), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n623), .B(KEYINPUT82), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G55), .A2(n659), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n675) );
  NAND2_X1 U707 ( .A1(G559), .A2(n841), .ZN(n628) );
  XOR2_X1 U708 ( .A(n998), .B(n628), .Z(n672) );
  XNOR2_X1 U709 ( .A(KEYINPUT81), .B(n672), .ZN(n629) );
  NOR2_X1 U710 ( .A1(G860), .A2(n629), .ZN(n630) );
  XOR2_X1 U711 ( .A(n675), .B(n630), .Z(G145) );
  NAND2_X1 U712 ( .A1(G75), .A2(n654), .ZN(n631) );
  XNOR2_X1 U713 ( .A(n631), .B(KEYINPUT86), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G62), .A2(n663), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G50), .A2(n659), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n634) );
  XOR2_X1 U717 ( .A(KEYINPUT84), .B(n634), .Z(n635) );
  NAND2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G88), .A2(n655), .ZN(n637) );
  XNOR2_X1 U720 ( .A(KEYINPUT85), .B(n637), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n639), .A2(n638), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G73), .A2(n654), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n640), .B(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n663), .A2(G61), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U726 ( .A1(G86), .A2(n655), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G48), .A2(n659), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U730 ( .A(KEYINPUT83), .B(n647), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G49), .A2(n659), .ZN(n650) );
  NAND2_X1 U732 ( .A1(G87), .A2(n648), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U734 ( .A1(n663), .A2(n651), .ZN(n653) );
  NAND2_X1 U735 ( .A1(G651), .A2(G74), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n653), .A2(n652), .ZN(G288) );
  NAND2_X1 U737 ( .A1(G72), .A2(n654), .ZN(n657) );
  NAND2_X1 U738 ( .A1(G85), .A2(n655), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U740 ( .A(KEYINPUT68), .B(n658), .ZN(n662) );
  NAND2_X1 U741 ( .A1(G47), .A2(n659), .ZN(n660) );
  XNOR2_X1 U742 ( .A(KEYINPUT69), .B(n660), .ZN(n661) );
  NOR2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n665) );
  NAND2_X1 U744 ( .A1(n663), .A2(G60), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n665), .A2(n664), .ZN(G290) );
  XNOR2_X1 U746 ( .A(G166), .B(G305), .ZN(n671) );
  XNOR2_X1 U747 ( .A(KEYINPUT19), .B(KEYINPUT87), .ZN(n667) );
  XNOR2_X1 U748 ( .A(G288), .B(n917), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U750 ( .A(n675), .B(n668), .Z(n669) );
  XNOR2_X1 U751 ( .A(n669), .B(G290), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n671), .B(n670), .ZN(n840) );
  XNOR2_X1 U753 ( .A(n840), .B(n672), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n673), .A2(G868), .ZN(n674) );
  XNOR2_X1 U755 ( .A(n674), .B(KEYINPUT88), .ZN(n678) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U762 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XOR2_X1 U763 ( .A(KEYINPUT89), .B(G44), .Z(n683) );
  XNOR2_X1 U764 ( .A(KEYINPUT3), .B(n683), .ZN(G218) );
  NOR2_X1 U765 ( .A1(G236), .A2(G237), .ZN(n684) );
  NAND2_X1 U766 ( .A1(G69), .A2(n684), .ZN(n685) );
  XNOR2_X1 U767 ( .A(KEYINPUT91), .B(n685), .ZN(n686) );
  NAND2_X1 U768 ( .A1(n686), .A2(G108), .ZN(n838) );
  NAND2_X1 U769 ( .A1(n838), .A2(G567), .ZN(n692) );
  NOR2_X1 U770 ( .A1(G220), .A2(G219), .ZN(n687) );
  XOR2_X1 U771 ( .A(KEYINPUT22), .B(n687), .Z(n688) );
  NOR2_X1 U772 ( .A1(G218), .A2(n688), .ZN(n689) );
  XNOR2_X1 U773 ( .A(KEYINPUT90), .B(n689), .ZN(n690) );
  NAND2_X1 U774 ( .A1(n690), .A2(G96), .ZN(n839) );
  NAND2_X1 U775 ( .A1(n839), .A2(G2106), .ZN(n691) );
  NAND2_X1 U776 ( .A1(n692), .A2(n691), .ZN(n916) );
  NAND2_X1 U777 ( .A1(G661), .A2(G483), .ZN(n693) );
  XNOR2_X1 U778 ( .A(KEYINPUT92), .B(n693), .ZN(n694) );
  NOR2_X1 U779 ( .A1(n916), .A2(n694), .ZN(n837) );
  NAND2_X1 U780 ( .A1(G36), .A2(n837), .ZN(n695) );
  XOR2_X1 U781 ( .A(KEYINPUT93), .B(n695), .Z(G176) );
  XOR2_X1 U782 ( .A(KEYINPUT94), .B(G166), .Z(G303) );
  NOR2_X1 U783 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U784 ( .A(KEYINPUT24), .B(KEYINPUT102), .Z(n696) );
  XNOR2_X1 U785 ( .A(KEYINPUT101), .B(n696), .ZN(n697) );
  XNOR2_X1 U786 ( .A(n698), .B(n697), .ZN(n702) );
  XNOR2_X1 U787 ( .A(n699), .B(KEYINPUT64), .ZN(n783) );
  NAND2_X1 U788 ( .A1(G160), .A2(G40), .ZN(n784) );
  AND2_X1 U789 ( .A1(n702), .A2(n774), .ZN(n766) );
  INV_X1 U790 ( .A(KEYINPUT106), .ZN(n764) );
  NOR2_X1 U791 ( .A1(n717), .A2(G1961), .ZN(n704) );
  XNOR2_X1 U792 ( .A(n704), .B(KEYINPUT103), .ZN(n706) );
  XNOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .ZN(n921) );
  NAND2_X1 U794 ( .A1(n717), .A2(n921), .ZN(n705) );
  NAND2_X1 U795 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U796 ( .A(KEYINPUT104), .B(n707), .ZN(n737) );
  NAND2_X1 U797 ( .A1(G171), .A2(n737), .ZN(n731) );
  NAND2_X1 U798 ( .A1(n717), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U799 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  INV_X1 U800 ( .A(G1956), .ZN(n946) );
  NOR2_X1 U801 ( .A1(n946), .A2(n717), .ZN(n709) );
  NOR2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n712) );
  NOR2_X1 U803 ( .A1(n917), .A2(n712), .ZN(n711) );
  XOR2_X1 U804 ( .A(n711), .B(KEYINPUT28), .Z(n728) );
  NAND2_X1 U805 ( .A1(n917), .A2(n712), .ZN(n726) );
  AND2_X1 U806 ( .A1(n717), .A2(G1996), .ZN(n713) );
  XOR2_X1 U807 ( .A(n713), .B(KEYINPUT26), .Z(n715) );
  NAND2_X1 U808 ( .A1(n744), .A2(G1341), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U810 ( .A1(n998), .A2(n716), .ZN(n721) );
  NAND2_X1 U811 ( .A1(G1348), .A2(n744), .ZN(n719) );
  NAND2_X1 U812 ( .A1(G2067), .A2(n717), .ZN(n718) );
  NAND2_X1 U813 ( .A1(n719), .A2(n718), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n1004), .A2(n722), .ZN(n720) );
  OR2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n1004), .A2(n722), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U820 ( .A(KEYINPUT29), .B(n729), .Z(n730) );
  NAND2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n743) );
  INV_X1 U822 ( .A(G1966), .ZN(n732) );
  INV_X1 U823 ( .A(G8), .ZN(n733) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n744), .ZN(n752) );
  OR2_X1 U825 ( .A1(n733), .A2(n752), .ZN(n734) );
  XNOR2_X1 U826 ( .A(KEYINPUT30), .B(n735), .ZN(n736) );
  NOR2_X1 U827 ( .A1(G168), .A2(n736), .ZN(n739) );
  NOR2_X1 U828 ( .A1(G171), .A2(n737), .ZN(n738) );
  NOR2_X1 U829 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n743), .A2(n742), .ZN(n754) );
  NAND2_X1 U831 ( .A1(n754), .A2(G286), .ZN(n749) );
  INV_X1 U832 ( .A(n774), .ZN(n761) );
  NOR2_X1 U833 ( .A1(n761), .A2(G1971), .ZN(n746) );
  NOR2_X1 U834 ( .A1(G2090), .A2(n744), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n747), .A2(G303), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n750), .A2(G8), .ZN(n751) );
  NAND2_X1 U839 ( .A1(G8), .A2(n752), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U842 ( .A1(n521), .A2(n757), .ZN(n768) );
  INV_X1 U843 ( .A(n768), .ZN(n760) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U845 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U848 ( .A(n764), .B(n763), .ZN(n765) );
  NOR2_X1 U849 ( .A1(n766), .A2(n765), .ZN(n782) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n1001) );
  AND2_X1 U851 ( .A1(n1001), .A2(KEYINPUT33), .ZN(n767) );
  NAND2_X1 U852 ( .A1(n767), .A2(n774), .ZN(n780) );
  XNOR2_X1 U853 ( .A(G1981), .B(G305), .ZN(n1016) );
  NOR2_X1 U854 ( .A1(n768), .A2(n1001), .ZN(n773) );
  NOR2_X1 U855 ( .A1(G303), .A2(G1971), .ZN(n769) );
  XNOR2_X1 U856 ( .A(n769), .B(KEYINPUT105), .ZN(n771) );
  INV_X1 U857 ( .A(KEYINPUT33), .ZN(n770) );
  AND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U859 ( .A1(n773), .A2(n772), .ZN(n777) );
  NAND2_X1 U860 ( .A1(G1976), .A2(G288), .ZN(n1002) );
  AND2_X1 U861 ( .A1(n774), .A2(n1002), .ZN(n775) );
  OR2_X1 U862 ( .A1(KEYINPUT33), .A2(n775), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U864 ( .A1(n1016), .A2(n778), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U866 ( .A1(n782), .A2(n781), .ZN(n816) );
  NOR2_X1 U867 ( .A1(n784), .A2(n783), .ZN(n829) );
  NAND2_X1 U868 ( .A1(n545), .A2(G105), .ZN(n785) );
  XNOR2_X1 U869 ( .A(n785), .B(KEYINPUT38), .ZN(n792) );
  NAND2_X1 U870 ( .A1(G129), .A2(n898), .ZN(n787) );
  NAND2_X1 U871 ( .A1(G141), .A2(n893), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G117), .A2(n896), .ZN(n788) );
  XNOR2_X1 U874 ( .A(KEYINPUT97), .B(n788), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U876 ( .A1(n792), .A2(n791), .ZN(n888) );
  NAND2_X1 U877 ( .A1(n888), .A2(G1996), .ZN(n801) );
  NAND2_X1 U878 ( .A1(G119), .A2(n898), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G107), .A2(n896), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U881 ( .A(KEYINPUT96), .B(n795), .Z(n799) );
  NAND2_X1 U882 ( .A1(G131), .A2(n893), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G95), .A2(n545), .ZN(n796) );
  AND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n904) );
  NAND2_X1 U886 ( .A1(G1991), .A2(n904), .ZN(n800) );
  NAND2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U888 ( .A(n802), .B(KEYINPUT98), .ZN(n985) );
  NAND2_X1 U889 ( .A1(n829), .A2(n985), .ZN(n803) );
  XNOR2_X1 U890 ( .A(n803), .B(KEYINPUT99), .ZN(n821) );
  INV_X1 U891 ( .A(n821), .ZN(n814) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NAND2_X1 U893 ( .A1(n893), .A2(G140), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT95), .B(n804), .Z(n806) );
  NAND2_X1 U895 ( .A1(n545), .A2(G104), .ZN(n805) );
  NAND2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n807), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G128), .A2(n898), .ZN(n809) );
  NAND2_X1 U899 ( .A1(G116), .A2(n896), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U901 ( .A(KEYINPUT35), .B(n810), .Z(n811) );
  NOR2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n813), .ZN(n907) );
  NOR2_X1 U904 ( .A1(n826), .A2(n907), .ZN(n982) );
  NAND2_X1 U905 ( .A1(n829), .A2(n982), .ZN(n824) );
  NAND2_X1 U906 ( .A1(n814), .A2(n824), .ZN(n815) );
  NOR2_X1 U907 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n1008) );
  NAND2_X1 U909 ( .A1(n1008), .A2(n829), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n832) );
  NOR2_X1 U911 ( .A1(G1996), .A2(n888), .ZN(n975) );
  NOR2_X1 U912 ( .A1(G1986), .A2(G290), .ZN(n819) );
  NOR2_X1 U913 ( .A1(G1991), .A2(n904), .ZN(n980) );
  NOR2_X1 U914 ( .A1(n819), .A2(n980), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U916 ( .A1(n975), .A2(n822), .ZN(n823) );
  XNOR2_X1 U917 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n826), .A2(n907), .ZN(n989) );
  NAND2_X1 U920 ( .A1(n827), .A2(n989), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U922 ( .A(KEYINPUT107), .B(n830), .Z(n831) );
  NAND2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U924 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U927 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U931 ( .A(G108), .ZN(G238) );
  INV_X1 U932 ( .A(G96), .ZN(G221) );
  NOR2_X1 U933 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(G286), .B(n840), .ZN(n843) );
  XNOR2_X1 U936 ( .A(n998), .B(n841), .ZN(n842) );
  XNOR2_X1 U937 ( .A(n843), .B(n842), .ZN(n844) );
  XNOR2_X1 U938 ( .A(G171), .B(n844), .ZN(n845) );
  NOR2_X1 U939 ( .A1(G37), .A2(n845), .ZN(G397) );
  XOR2_X1 U940 ( .A(KEYINPUT112), .B(G1956), .Z(n847) );
  XNOR2_X1 U941 ( .A(G1981), .B(G1966), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U943 ( .A(n848), .B(KEYINPUT41), .Z(n850) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U946 ( .A(G1986), .B(G1971), .Z(n852) );
  XNOR2_X1 U947 ( .A(G1976), .B(G1961), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U949 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U950 ( .A(KEYINPUT111), .B(G2474), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U952 ( .A(KEYINPUT109), .B(G2678), .Z(n858) );
  XNOR2_X1 U953 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U955 ( .A(KEYINPUT110), .B(G2090), .Z(n860) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U958 ( .A(n862), .B(n861), .Z(n864) );
  XNOR2_X1 U959 ( .A(G2096), .B(G2100), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n866) );
  XOR2_X1 U961 ( .A(G2078), .B(G2084), .Z(n865) );
  XNOR2_X1 U962 ( .A(n866), .B(n865), .ZN(G227) );
  NAND2_X1 U963 ( .A1(G124), .A2(n898), .ZN(n867) );
  XOR2_X1 U964 ( .A(KEYINPUT113), .B(n867), .Z(n868) );
  XNOR2_X1 U965 ( .A(n868), .B(KEYINPUT44), .ZN(n870) );
  NAND2_X1 U966 ( .A1(G112), .A2(n896), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n870), .A2(n869), .ZN(n874) );
  NAND2_X1 U968 ( .A1(G136), .A2(n893), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G100), .A2(n545), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  NOR2_X1 U971 ( .A1(n874), .A2(n873), .ZN(G162) );
  NAND2_X1 U972 ( .A1(G130), .A2(n898), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G118), .A2(n896), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U975 ( .A1(G142), .A2(n893), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G106), .A2(n545), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  XNOR2_X1 U979 ( .A(KEYINPUT114), .B(n880), .ZN(n881) );
  NOR2_X1 U980 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U981 ( .A(G164), .B(n883), .ZN(n887) );
  XOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n885) );
  XNOR2_X1 U983 ( .A(KEYINPUT117), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n892) );
  XNOR2_X1 U986 ( .A(n979), .B(G162), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n888), .B(G160), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n906) );
  NAND2_X1 U990 ( .A1(G139), .A2(n893), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G103), .A2(n545), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n903) );
  NAND2_X1 U993 ( .A1(n896), .A2(G115), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n897), .B(KEYINPUT116), .ZN(n900) );
  NAND2_X1 U995 ( .A1(G127), .A2(n898), .ZN(n899) );
  NAND2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U998 ( .A1(n903), .A2(n902), .ZN(n969) );
  XNOR2_X1 U999 ( .A(n904), .B(n969), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1001 ( .A(n908), .B(n907), .Z(n909) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n916), .ZN(n913) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n911), .ZN(n912) );
  NAND2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(n914), .A2(G395), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1010 ( .A(G308), .ZN(G225) );
  INV_X1 U1011 ( .A(n916), .ZN(G319) );
  INV_X1 U1012 ( .A(G69), .ZN(G235) );
  INV_X1 U1013 ( .A(n917), .ZN(G299) );
  XNOR2_X1 U1014 ( .A(KEYINPUT121), .B(G2090), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(n918), .B(G35), .ZN(n936) );
  XNOR2_X1 U1016 ( .A(G1996), .B(G32), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(G26), .B(G2067), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n925) );
  XOR2_X1 U1019 ( .A(n921), .B(G27), .Z(n923) );
  XNOR2_X1 U1020 ( .A(G2072), .B(G33), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n929) );
  XOR2_X1 U1023 ( .A(G1991), .B(G25), .Z(n926) );
  NAND2_X1 U1024 ( .A1(n926), .A2(G28), .ZN(n927) );
  XNOR2_X1 U1025 ( .A(KEYINPUT122), .B(n927), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(n930), .B(KEYINPUT123), .Z(n931) );
  XNOR2_X1 U1028 ( .A(KEYINPUT53), .B(n931), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G34), .B(G2084), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(KEYINPUT54), .B(n932), .ZN(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(G29), .A2(KEYINPUT55), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n937), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(G11), .A2(n938), .ZN(n968) );
  INV_X1 U1036 ( .A(KEYINPUT55), .ZN(n993) );
  OR2_X1 U1037 ( .A1(n993), .A2(n939), .ZN(n966) );
  XOR2_X1 U1038 ( .A(G1986), .B(G24), .Z(n943) );
  XNOR2_X1 U1039 ( .A(G1976), .B(G23), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G22), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(n945), .B(n944), .ZN(n961) );
  XOR2_X1 U1045 ( .A(G1961), .B(G5), .Z(n956) );
  XNOR2_X1 U1046 ( .A(G20), .B(n946), .ZN(n950) );
  XNOR2_X1 U1047 ( .A(G1981), .B(G6), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(G1341), .B(G19), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n953) );
  XOR2_X1 U1051 ( .A(KEYINPUT59), .B(G1348), .Z(n951) );
  XNOR2_X1 U1052 ( .A(G4), .B(n951), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT60), .B(n954), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(G21), .B(G1966), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(KEYINPUT126), .B(n957), .ZN(n958) );
  NOR2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1060 ( .A(KEYINPUT61), .B(n962), .Z(n964) );
  INV_X1 U1061 ( .A(G16), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n997) );
  XOR2_X1 U1065 ( .A(G164), .B(G2078), .Z(n972) );
  XOR2_X1 U1066 ( .A(n969), .B(KEYINPUT120), .Z(n970) );
  XNOR2_X1 U1067 ( .A(G2072), .B(n970), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1069 ( .A(KEYINPUT50), .B(n973), .ZN(n978) );
  XOR2_X1 U1070 ( .A(G2090), .B(G162), .Z(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1072 ( .A(KEYINPUT51), .B(n976), .Z(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n991) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n984) );
  XOR2_X1 U1075 ( .A(G160), .B(G2084), .Z(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1079 ( .A(KEYINPUT119), .B(n987), .Z(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT52), .B(n992), .ZN(n994) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n995), .A2(G29), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1025) );
  XOR2_X1 U1086 ( .A(G16), .B(KEYINPUT56), .Z(n1023) );
  XNOR2_X1 U1087 ( .A(G301), .B(G1961), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(n998), .B(G1341), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1014) );
  INV_X1 U1090 ( .A(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1348), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G299), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(G1971), .B(G303), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1020) );
  XOR2_X1 U1100 ( .A(G1966), .B(G168), .Z(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT124), .B(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT57), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT125), .B(n1021), .Z(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1107 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1108 ( .A(n1026), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

