//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT81), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G143), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n189), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n193), .A2(KEYINPUT65), .A3(new_n195), .A4(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n189), .A2(G143), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT64), .B(G146), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n196), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n201), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n193), .A2(new_n195), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n193), .A2(KEYINPUT68), .A3(new_n195), .A4(new_n211), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G128), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n214), .A2(new_n215), .B1(new_n217), .B2(new_n204), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n188), .B1(new_n209), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n199), .A2(new_n200), .B1(new_n204), .B2(new_n206), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(new_n219), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT81), .ZN(new_n224));
  OAI211_X1 g038(.A(G224), .B(new_n187), .C1(new_n221), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n224), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n187), .A2(G224), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n214), .A2(new_n215), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(new_n203), .B2(G143), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n204), .B1(new_n230), .B2(new_n210), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n228), .A2(new_n219), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT81), .B1(new_n223), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n226), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G107), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G104), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(new_n236), .A3(G104), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n239), .B2(KEYINPUT3), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n238), .A2(new_n241), .A3(new_n236), .A4(G104), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(G101), .ZN(new_n245));
  XOR2_X1   g059(.A(G116), .B(G119), .Z(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G101), .ZN(new_n251));
  AOI211_X1 g065(.A(KEYINPUT75), .B(new_n251), .C1(new_n240), .C2(new_n242), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g067(.A(G104), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G107), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n251), .A3(new_n242), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT4), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n243), .A2(G101), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT75), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT76), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT75), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n254), .A2(KEYINPUT74), .A3(G107), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n255), .B1(new_n263), .B2(new_n241), .ZN(new_n264));
  INV_X1    g078(.A(new_n242), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n262), .B(G101), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n256), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT76), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n262), .B1(new_n243), .B2(G101), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n250), .B1(new_n261), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n272));
  INV_X1    g086(.A(G119), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(G116), .ZN(new_n274));
  OAI211_X1 g088(.A(G113), .B(new_n274), .C1(new_n246), .C2(new_n272), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n246), .B2(new_n247), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n254), .A2(G107), .ZN(new_n277));
  OAI21_X1  g091(.A(G101), .B1(new_n277), .B2(new_n237), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n256), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G110), .B(G122), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n271), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n282), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n285));
  INV_X1    g099(.A(new_n257), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n260), .A2(KEYINPUT76), .A3(new_n286), .A4(new_n266), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n249), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n288), .B2(new_n280), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n289), .A3(KEYINPUT6), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n271), .A2(new_n281), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n282), .A2(KEYINPUT6), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n291), .B(new_n293), .C1(new_n288), .C2(new_n280), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n235), .B(new_n290), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n298));
  AOI22_X1  g112(.A1(KEYINPUT82), .A2(new_n298), .B1(new_n187), .B2(G224), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(KEYINPUT82), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n223), .B2(new_n232), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n282), .B(KEYINPUT8), .ZN(new_n302));
  AND2_X1   g116(.A1(new_n276), .A2(new_n279), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n303), .B2(new_n280), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n288), .A2(new_n280), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(new_n282), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n226), .A2(KEYINPUT7), .A3(new_n233), .A4(new_n227), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n297), .A2(new_n309), .A3(new_n311), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(KEYINPUT83), .A3(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT83), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n317), .A3(new_n312), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT16), .ZN(new_n321));
  INV_X1    g135(.A(G140), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G125), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n321), .B1(KEYINPUT16), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n189), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n321), .B(G146), .C1(KEYINPUT16), .C2(new_n323), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n273), .A2(G128), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n273), .A2(G128), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(KEYINPUT23), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G110), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n334), .B(new_n335), .C1(new_n273), .C2(G128), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n327), .B(new_n332), .C1(new_n333), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n333), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(G110), .B2(new_n331), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n203), .A2(new_n320), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n326), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G137), .ZN(new_n343));
  INV_X1    g157(.A(G221), .ZN(new_n344));
  INV_X1    g158(.A(G234), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n344), .A2(new_n345), .A3(G953), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n343), .B(new_n346), .Z(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G902), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n337), .A2(new_n341), .A3(new_n347), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT25), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G217), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(G234), .B2(new_n350), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n349), .A2(new_n351), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(G902), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n354), .A2(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G472), .ZN(new_n361));
  INV_X1    g175(.A(G134), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT66), .B1(new_n362), .B2(G137), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT11), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT11), .ZN(new_n365));
  OAI211_X1 g179(.A(KEYINPUT66), .B(new_n365), .C1(new_n362), .C2(G137), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n362), .A2(G137), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G131), .ZN(new_n369));
  INV_X1    g183(.A(G131), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n364), .A2(new_n370), .A3(new_n366), .A4(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n372), .A2(new_n201), .A3(new_n207), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n362), .A2(KEYINPUT67), .A3(G137), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n362), .A2(G137), .ZN(new_n377));
  OAI211_X1 g191(.A(G131), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n228), .B2(new_n231), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n373), .A2(new_n380), .A3(KEYINPUT30), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n228), .A2(new_n231), .ZN(new_n383));
  INV_X1    g197(.A(new_n379), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n222), .A2(new_n372), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n248), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT31), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n390));
  NOR2_X1   g204(.A1(G237), .A2(G953), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G210), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n390), .B(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT26), .B(G101), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n248), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n385), .A2(new_n397), .A3(new_n386), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n388), .A2(new_n389), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT28), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n248), .B1(new_n373), .B2(new_n380), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(new_n398), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n373), .A2(new_n380), .A3(new_n248), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT28), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n395), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT30), .B1(new_n373), .B2(new_n380), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n385), .A2(new_n382), .A3(new_n386), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n403), .B1(new_n409), .B2(new_n248), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n389), .B1(new_n410), .B2(new_n396), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n361), .B(new_n350), .C1(new_n406), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT32), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n388), .A2(new_n396), .A3(new_n398), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT31), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(new_n405), .A3(new_n399), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT32), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n416), .A2(new_n417), .A3(new_n361), .A4(new_n350), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  OR3_X1    g233(.A1(new_n410), .A2(KEYINPUT70), .A3(new_n396), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT70), .B1(new_n410), .B2(new_n396), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n402), .A2(new_n404), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT29), .B1(new_n422), .B2(new_n396), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n402), .ZN(new_n425));
  INV_X1    g239(.A(new_n404), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT29), .A4(new_n396), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT71), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT71), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n422), .A2(new_n429), .A3(KEYINPUT29), .A4(new_n396), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n430), .A3(new_n350), .ZN(new_n431));
  OAI21_X1  g245(.A(G472), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n360), .B1(new_n419), .B2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT9), .B(G234), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n344), .B1(new_n435), .B2(new_n350), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT79), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n187), .A2(G227), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT73), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT78), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT10), .ZN(new_n444));
  INV_X1    g258(.A(new_n279), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(new_n383), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n193), .A2(new_n195), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G128), .ZN(new_n449));
  AOI22_X1  g263(.A1(new_n214), .A2(new_n215), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(KEYINPUT10), .A3(new_n279), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n222), .A2(new_n245), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n285), .B2(new_n287), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n452), .A2(new_n454), .A3(new_n372), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT77), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n372), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n194), .B1(new_n203), .B2(G143), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT68), .B1(new_n459), .B2(new_n211), .ZN(new_n460));
  INV_X1    g274(.A(new_n215), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n231), .B(new_n279), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n447), .A2(new_n449), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n279), .B1(new_n228), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n458), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT12), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n462), .B1(new_n279), .B2(new_n450), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT12), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n458), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n443), .B1(new_n455), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n464), .B1(new_n460), .B2(new_n461), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n445), .ZN(new_n474));
  AOI211_X1 g288(.A(KEYINPUT12), .B(new_n457), .C1(new_n474), .C2(new_n462), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n469), .B1(new_n468), .B2(new_n458), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n453), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n261), .B2(new_n270), .ZN(new_n479));
  INV_X1    g293(.A(new_n372), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT10), .B1(new_n218), .B2(new_n279), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(KEYINPUT10), .B2(new_n474), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(KEYINPUT78), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n442), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n455), .A2(new_n441), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n372), .B1(new_n452), .B2(new_n454), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n437), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n477), .A2(KEYINPUT78), .A3(new_n483), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT78), .B1(new_n477), .B2(new_n483), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n441), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n486), .A2(new_n487), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(KEYINPUT79), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n494), .A3(G469), .ZN(new_n495));
  INV_X1    g309(.A(G469), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(new_n350), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n487), .A2(new_n483), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n441), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n477), .A2(new_n442), .A3(new_n483), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n497), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n436), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G475), .A2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n391), .A2(G143), .A3(G214), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(G143), .B1(new_n391), .B2(G214), .ZN(new_n508));
  OAI21_X1  g322(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n508), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n370), .A3(new_n506), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n203), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n219), .A2(G140), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n323), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT19), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n512), .B(new_n326), .C1(new_n513), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(new_n506), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT18), .A3(G131), .ZN(new_n519));
  NAND2_X1  g333(.A1(KEYINPUT18), .A2(G131), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n510), .A2(new_n506), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n515), .A2(G146), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT84), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n340), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n340), .B2(new_n522), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n519), .B(new_n521), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(new_n254), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n529), .B(KEYINPUT85), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n509), .A2(new_n511), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n518), .A2(KEYINPUT17), .A3(G131), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n534), .A2(new_n325), .A3(new_n535), .A4(new_n326), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n536), .A3(new_n526), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n505), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT86), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n537), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n529), .B1(new_n536), .B2(new_n526), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n350), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G475), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT20), .B1(new_n538), .B2(KEYINPUT86), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n540), .B(new_n505), .C1(new_n531), .C2(new_n537), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n542), .B(new_n546), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G143), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n210), .A2(G143), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(G134), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(G116), .B(G122), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n236), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n556), .A2(new_n236), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n210), .A2(G143), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(KEYINPUT13), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(KEYINPUT13), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n561), .A2(new_n562), .A3(new_n552), .ZN(new_n563));
  OAI221_X1 g377(.A(new_n555), .B1(new_n558), .B2(new_n559), .C1(new_n563), .C2(new_n362), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n362), .B1(new_n551), .B2(new_n552), .ZN(new_n565));
  OR3_X1    g379(.A1(new_n554), .A2(KEYINPUT87), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT87), .B1(new_n554), .B2(new_n565), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n557), .ZN(new_n568));
  INV_X1    g382(.A(G116), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G122), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n569), .A2(G122), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(KEYINPUT14), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT88), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(new_n570), .C1(new_n571), .C2(KEYINPUT14), .ZN(new_n575));
  OR3_X1    g389(.A1(new_n570), .A2(KEYINPUT89), .A3(KEYINPUT14), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT89), .B1(new_n570), .B2(KEYINPUT14), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n573), .A2(new_n575), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  AND2_X1   g392(.A1(new_n578), .A2(G107), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n564), .B1(new_n568), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n434), .A2(new_n355), .A3(G953), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n564), .B(new_n581), .C1(new_n568), .C2(new_n579), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n350), .ZN(new_n586));
  INV_X1    g400(.A(G478), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n586), .B(new_n588), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n549), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n187), .A2(G952), .ZN(new_n591));
  INV_X1    g405(.A(G237), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n345), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI211_X1 g408(.A(new_n350), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT21), .B(G898), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n319), .A2(new_n433), .A3(new_n503), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n495), .A2(new_n502), .ZN(new_n601));
  INV_X1    g415(.A(new_n436), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n350), .B1(new_n406), .B2(new_n411), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G472), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n604), .A2(new_n412), .A3(new_n359), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n549), .ZN(new_n608));
  NOR2_X1   g422(.A1(KEYINPUT91), .A2(G478), .ZN(new_n609));
  AND2_X1   g423(.A1(KEYINPUT91), .A2(G478), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n586), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n587), .A2(G902), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n583), .A2(new_n613), .A3(new_n584), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n583), .B2(new_n584), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n597), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n297), .A2(KEYINPUT90), .A3(new_n309), .A4(new_n311), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n316), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT90), .B1(new_n310), .B2(new_n312), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n314), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n607), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT92), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND2_X1  g444(.A1(new_n608), .A2(new_n589), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n597), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n607), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  AND2_X1   g450(.A1(new_n352), .A2(new_n353), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n352), .A2(new_n353), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n356), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n348), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n342), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n358), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n604), .A2(new_n412), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  AND4_X1   g459(.A1(new_n319), .A2(new_n503), .A3(new_n598), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT37), .B(G110), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  INV_X1    g462(.A(KEYINPUT94), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n419), .A2(new_n432), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n625), .A3(new_n643), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n593), .B(KEYINPUT93), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n654), .B2(new_n595), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n608), .A2(new_n589), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n601), .A2(new_n602), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n649), .B1(new_n651), .B2(new_n659), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n436), .B(new_n657), .C1(new_n495), .C2(new_n502), .ZN(new_n661));
  INV_X1    g475(.A(new_n643), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n419), .B2(new_n432), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n661), .A2(KEYINPUT94), .A3(new_n625), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  NAND2_X1  g480(.A1(new_n315), .A2(new_n318), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT38), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n410), .A2(new_n395), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n401), .A2(new_n398), .A3(new_n395), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n350), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n419), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n549), .A2(new_n589), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n662), .A2(new_n316), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n669), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT95), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n655), .B(KEYINPUT39), .Z(new_n681));
  AND2_X1   g495(.A1(new_n503), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT96), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT96), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n680), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n550), .ZN(G45));
  NAND3_X1  g503(.A1(new_n549), .A2(new_n617), .A3(new_n656), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT97), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT97), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n549), .A2(new_n617), .A3(new_n692), .A4(new_n656), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n663), .A2(new_n503), .A3(new_n625), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  NAND2_X1  g511(.A1(new_n650), .A2(new_n359), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n486), .A2(new_n477), .B1(new_n498), .B2(new_n441), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n501), .A2(new_n496), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n699), .B1(new_n703), .B2(new_n436), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT98), .A4(new_n602), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n698), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n626), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n633), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G116), .ZN(G18));
  INV_X1    g526(.A(new_n651), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n704), .A2(new_n598), .A3(new_n705), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G119), .ZN(G21));
  INV_X1    g530(.A(new_n597), .ZN(new_n717));
  AND4_X1   g531(.A1(new_n717), .A2(new_n704), .A3(new_n605), .A4(new_n705), .ZN(new_n718));
  INV_X1    g532(.A(new_n625), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n676), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR2_X1   g536(.A1(new_n694), .A2(new_n644), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n723), .A2(new_n625), .A3(new_n704), .A4(new_n705), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G125), .ZN(G27));
  INV_X1    g539(.A(new_n316), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n315), .B2(new_n318), .ZN(new_n727));
  XOR2_X1   g541(.A(new_n497), .B(KEYINPUT99), .Z(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n501), .B2(new_n496), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n492), .A2(G469), .A3(new_n493), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n436), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n433), .A2(new_n727), .A3(new_n695), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  NAND2_X1  g552(.A1(new_n314), .A2(KEYINPUT83), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n311), .B1(new_n297), .B2(new_n309), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n318), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n732), .B(new_n316), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(KEYINPUT100), .A3(new_n433), .A4(new_n658), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n433), .A2(new_n727), .A3(new_n658), .A4(new_n732), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT100), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  AOI21_X1  g564(.A(KEYINPUT45), .B1(new_n489), .B2(new_n494), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n492), .A2(KEYINPUT45), .A3(new_n493), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(G469), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT46), .A3(new_n728), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n728), .B1(new_n751), .B2(new_n753), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n702), .A3(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n759), .A2(new_n602), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT101), .A3(new_n681), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT101), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n602), .ZN(new_n763));
  INV_X1    g577(.A(new_n681), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n662), .B1(new_n412), .B2(new_n604), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT103), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT102), .B1(new_n608), .B2(new_n617), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT43), .Z(new_n769));
  AND3_X1   g583(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT44), .B1(new_n767), .B2(new_n769), .ZN(new_n771));
  INV_X1    g585(.A(new_n727), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n761), .A2(new_n765), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  OR3_X1    g590(.A1(new_n760), .A2(KEYINPUT105), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT105), .B1(new_n760), .B2(new_n776), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT104), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n763), .B2(KEYINPUT47), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n760), .A2(KEYINPUT104), .A3(new_n776), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n777), .A2(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n772), .A2(new_n650), .A3(new_n359), .A4(new_n694), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NAND4_X1  g599(.A1(new_n632), .A2(new_n315), .A3(new_n316), .A4(new_n318), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n606), .B1(KEYINPUT108), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n646), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n319), .A2(new_n503), .A3(new_n605), .A4(new_n621), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n599), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT107), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n599), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n789), .A2(new_n792), .A3(KEYINPUT109), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n626), .A2(new_n707), .B1(new_n718), .B2(new_n720), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n707), .A2(new_n633), .B1(new_n713), .B2(new_n714), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n800), .B(new_n801), .C1(new_n735), .C2(new_n736), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n663), .A2(new_n727), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n590), .A2(new_n655), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n503), .A2(new_n804), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n803), .A2(new_n805), .B1(new_n744), .B2(new_n723), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n749), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT110), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n749), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n802), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n696), .A2(new_n724), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n643), .A2(new_n655), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT112), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n720), .A2(new_n674), .A3(new_n732), .A4(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n665), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n665), .A2(new_n812), .A3(KEYINPUT52), .A4(new_n815), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n799), .A2(new_n811), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n696), .A2(new_n724), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n660), .B2(new_n664), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n825), .B2(new_n815), .ZN(new_n826));
  AND4_X1   g640(.A1(KEYINPUT52), .A2(new_n665), .A3(new_n812), .A4(new_n815), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT113), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n818), .A2(new_n829), .A3(new_n819), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n799), .A2(new_n811), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n823), .A2(new_n833), .A3(KEYINPUT54), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n821), .A2(new_n822), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n832), .A2(KEYINPUT111), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n818), .A2(new_n829), .A3(new_n819), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n829), .B1(new_n818), .B2(new_n819), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(KEYINPUT111), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n836), .B1(new_n842), .B2(new_n822), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n835), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n769), .A2(new_n605), .A3(new_n653), .ZN(new_n847));
  OR3_X1    g661(.A1(new_n847), .A2(new_n316), .A3(new_n706), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT50), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n848), .A2(new_n849), .A3(new_n669), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n848), .B2(new_n669), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n772), .A2(new_n706), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n359), .A2(new_n853), .A3(new_n594), .A4(new_n675), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n549), .A2(new_n617), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n853), .A2(new_n653), .A3(new_n769), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(new_n645), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n846), .B1(new_n859), .B2(KEYINPUT115), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n847), .A2(new_n772), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n703), .A2(new_n602), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n861), .B1(new_n782), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n860), .B(new_n863), .C1(KEYINPUT115), .C2(new_n859), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n704), .A2(new_n625), .A3(new_n705), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n591), .B1(new_n847), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n433), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT48), .Z(new_n868));
  AOI211_X1 g682(.A(new_n866), .B(new_n868), .C1(new_n619), .C2(new_n854), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n858), .A2(KEYINPUT114), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n858), .A2(KEYINPUT114), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n870), .A2(new_n863), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n864), .B(new_n869), .C1(new_n872), .C2(KEYINPUT51), .ZN(new_n873));
  OAI22_X1  g687(.A1(new_n845), .A2(new_n873), .B1(G952), .B2(G953), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n703), .A2(KEYINPUT49), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT106), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n703), .A2(KEYINPUT49), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n359), .A2(new_n316), .A3(new_n602), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n878), .A2(new_n549), .A3(new_n618), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n675), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  OR3_X1    g694(.A1(new_n669), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n874), .A2(new_n881), .ZN(G75));
  NOR2_X1   g696(.A1(new_n187), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n799), .A2(new_n811), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n840), .A3(KEYINPUT53), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n821), .A2(new_n822), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n350), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n290), .B1(new_n294), .B2(new_n296), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(new_n235), .Z(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT55), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n884), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(G210), .B(G902), .C1(new_n823), .C2(new_n833), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n892), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT116), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n883), .B1(new_n897), .B2(new_n892), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n889), .A2(new_n893), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(G51));
  XOR2_X1   g718(.A(new_n728), .B(KEYINPUT57), .Z(new_n905));
  AOI21_X1  g719(.A(new_n844), .B1(new_n886), .B2(new_n887), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(new_n834), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT117), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n700), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT117), .B(new_n905), .C1(new_n834), .C2(new_n906), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n823), .A2(new_n833), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n913), .A2(new_n350), .A3(new_n754), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n883), .B1(new_n912), .B2(new_n914), .ZN(G54));
  NAND2_X1  g729(.A1(new_n531), .A2(new_n537), .ZN(new_n916));
  AND2_X1   g730(.A1(KEYINPUT58), .A2(G475), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n888), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n888), .B2(new_n917), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n920), .A2(new_n921), .A3(new_n883), .A4(new_n922), .ZN(G60));
  OR2_X1    g737(.A1(new_n614), .A2(new_n615), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n925));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n845), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n924), .B(new_n927), .C1(new_n834), .C2(new_n906), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n884), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT60), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n641), .B(new_n934), .C1(new_n823), .C2(new_n833), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n913), .A2(new_n933), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n884), .B(new_n935), .C1(new_n936), .C2(new_n357), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G66));
  INV_X1    g753(.A(G224), .ZN(new_n940));
  OAI21_X1  g754(.A(G953), .B1(new_n596), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n890), .B1(G898), .B2(new_n187), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT120), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  INV_X1    g760(.A(G227), .ZN(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n947), .B2(new_n654), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n516), .B(KEYINPUT121), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n409), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(G953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n620), .A2(new_n631), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n682), .A2(new_n433), .A3(new_n727), .A4(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n774), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n784), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT62), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n685), .A2(new_n960), .A3(new_n687), .A4(new_n825), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT122), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n959), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n685), .A2(new_n687), .A3(new_n825), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(KEYINPUT62), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n967), .A2(new_n966), .A3(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n955), .B1(new_n965), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n654), .A2(G953), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n953), .A2(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n782), .A2(new_n783), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n698), .A2(new_n719), .A3(new_n676), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n761), .B(new_n765), .C1(new_n773), .C2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n737), .A3(new_n749), .A4(new_n825), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n974), .B1(new_n980), .B2(new_n187), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n950), .B(new_n951), .C1(new_n972), .C2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n959), .ZN(new_n983));
  INV_X1    g797(.A(new_n964), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n961), .A2(new_n962), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n970), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n968), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n954), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n973), .B(new_n953), .C1(new_n979), .C2(G953), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(new_n949), .A3(new_n948), .A4(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n982), .A2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(new_n420), .A2(new_n421), .ZN(new_n993));
  AOI22_X1  g807(.A1(new_n993), .A2(KEYINPUT127), .B1(new_n396), .B2(new_n410), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(KEYINPUT127), .B2(new_n993), .ZN(new_n995));
  XNOR2_X1  g809(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n843), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n998), .B(KEYINPUT126), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n979), .B2(new_n942), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n410), .A2(new_n395), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n884), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n965), .A2(new_n971), .A3(new_n942), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n1001), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n1000), .B(new_n1005), .C1(new_n1007), .C2(new_n670), .ZN(G57));
endmodule


