//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(new_n202), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n210), .A2(G20), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n214), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n213), .B(new_n217), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XOR2_X1   g0026(.A(G250), .B(G257), .Z(new_n227));
  XNOR2_X1  g0027(.A(G264), .B(G270), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n227), .B(new_n228), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n230), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G351));
  NOR2_X1   g0042(.A1(G20), .A2(G33), .ZN(new_n243));
  AOI22_X1  g0043(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G58), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n245), .A2(KEYINPUT8), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT70), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(KEYINPUT8), .ZN(new_n249));
  OR2_X1    g0049(.A1(new_n249), .A2(KEYINPUT69), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G20), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n244), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n211), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n260), .A3(new_n211), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G50), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n256), .A2(new_n263), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n266), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n265), .A2(G20), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G50), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1698), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G222), .ZN(new_n277));
  INV_X1    g0077(.A(G77), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n274), .A2(new_n275), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(G1698), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n277), .B1(new_n278), .B2(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G45), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n265), .A2(G274), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n295), .B1(G226), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n284), .A2(new_n285), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n284), .A2(new_n298), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n273), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n273), .B(KEYINPUT9), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(G200), .B2(new_n300), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n305), .B1(new_n304), .B2(new_n308), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT17), .ZN(new_n313));
  XNOR2_X1  g0113(.A(new_n246), .B(KEYINPUT70), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n314), .A2(new_n251), .A3(new_n250), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n315), .A2(new_n271), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n270), .B1(new_n267), .B2(new_n253), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n245), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n319), .B2(new_n202), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n243), .A2(G159), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NOR2_X1   g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT7), .B1(new_n325), .B2(new_n254), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NOR4_X1   g0127(.A1(new_n323), .A2(new_n324), .A3(new_n327), .A4(G20), .ZN(new_n328));
  OAI21_X1  g0128(.A(G68), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT78), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n322), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n274), .A2(new_n254), .A3(new_n275), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n327), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(KEYINPUT7), .A3(new_n254), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n318), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT78), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT16), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n322), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n329), .A2(KEYINPUT16), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n263), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n317), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n293), .A2(G232), .A3(new_n296), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT80), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT80), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n346), .A3(new_n343), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n306), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(G223), .A2(G1698), .ZN(new_n350));
  INV_X1    g0150(.A(G226), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n351), .B2(G1698), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n279), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G87), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n355), .A2(KEYINPUT79), .A3(new_n283), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT79), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n352), .A2(new_n279), .B1(G33), .B2(G87), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n358), .B2(new_n293), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n355), .A2(new_n283), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n345), .A2(new_n347), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G200), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n349), .A2(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n313), .B1(new_n341), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n315), .A2(new_n271), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n367), .A2(new_n269), .B1(new_n266), .B2(new_n315), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n338), .B1(new_n335), .B2(KEYINPUT78), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n329), .A2(new_n330), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n335), .A2(new_n322), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n262), .B1(new_n373), .B2(KEYINPUT16), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n368), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n345), .A2(new_n347), .A3(new_n362), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n345), .A2(new_n285), .A3(new_n347), .ZN(new_n377));
  OAI22_X1  g0177(.A1(new_n376), .A2(G169), .B1(new_n377), .B2(new_n360), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT18), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT18), .ZN(new_n380));
  INV_X1    g0180(.A(new_n377), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n361), .B1(new_n363), .B2(new_n301), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n341), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n376), .A2(G200), .B1(new_n348), .B2(new_n360), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n375), .A2(KEYINPUT17), .A3(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n366), .A2(new_n379), .A3(new_n383), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G97), .ZN(new_n389));
  INV_X1    g0189(.A(new_n276), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n388), .B(new_n389), .C1(new_n390), .C2(new_n351), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n283), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n295), .B1(G238), .B2(new_n297), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT13), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n392), .B2(new_n393), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G190), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n318), .A2(G20), .ZN(new_n399));
  INV_X1    g0199(.A(new_n243), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n399), .B1(new_n255), .B2(new_n278), .C1(new_n400), .C2(new_n264), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n263), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT11), .ZN(new_n403));
  INV_X1    g0203(.A(G13), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n404), .A2(G1), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT72), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(G20), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n266), .A2(KEYINPUT72), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n262), .A2(new_n409), .A3(G68), .A4(new_n271), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT12), .B1(new_n409), .B2(G68), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT12), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n411), .B1(new_n399), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n403), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G200), .B1(new_n395), .B2(new_n396), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n398), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(KEYINPUT76), .B(KEYINPUT14), .C1(new_n397), .C2(new_n301), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n421));
  OAI211_X1 g0221(.A(G169), .B(new_n421), .C1(new_n395), .C2(new_n396), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT77), .B1(new_n397), .B2(G179), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT77), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n395), .A2(new_n396), .A3(new_n424), .A4(new_n285), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n420), .B(new_n422), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n419), .B1(new_n426), .B2(new_n415), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n262), .A2(new_n409), .A3(G77), .A4(new_n271), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT73), .ZN(new_n429));
  INV_X1    g0229(.A(new_n409), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n278), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT71), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT8), .B(G58), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n433), .A2(new_n400), .B1(new_n254), .B2(new_n278), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT15), .B(G87), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(new_n255), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n432), .B1(new_n437), .B2(new_n262), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n263), .B(KEYINPUT71), .C1(new_n434), .C2(new_n436), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n429), .A2(new_n431), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT74), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n429), .A2(new_n440), .A3(KEYINPUT74), .A4(new_n431), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n297), .A2(G244), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n342), .ZN(new_n447));
  INV_X1    g0247(.A(G1698), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n279), .A2(G232), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n325), .A2(G107), .ZN(new_n450));
  INV_X1    g0250(.A(G238), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n449), .B(new_n450), .C1(new_n281), .C2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n447), .B1(new_n283), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G169), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT75), .B1(new_n453), .B2(new_n285), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(KEYINPUT75), .A3(new_n285), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n445), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n453), .A2(new_n364), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(G190), .B2(new_n453), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n443), .A2(new_n461), .A3(new_n444), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n312), .A2(new_n387), .A3(new_n427), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G116), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n257), .A2(new_n211), .B1(G20), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n254), .C1(G33), .C2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT20), .B1(new_n466), .B2(new_n469), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n470), .A2(new_n471), .B1(G116), .B2(new_n409), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n465), .B1(new_n265), .B2(G33), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n262), .A2(new_n409), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G264), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n476));
  OAI211_X1 g0276(.A(G257), .B(new_n448), .C1(new_n323), .C2(new_n324), .ZN(new_n477));
  INV_X1    g0277(.A(G303), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n279), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n283), .ZN(new_n480));
  XNOR2_X1  g0280(.A(KEYINPUT5), .B(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n286), .A2(G1), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n481), .A2(new_n482), .B1(new_n212), .B2(new_n292), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n265), .A2(G45), .A3(G274), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n212), .B2(new_n292), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n483), .A2(G270), .B1(new_n485), .B2(new_n481), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n486), .A3(G179), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT86), .B1(new_n475), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n481), .ZN(new_n489));
  AND2_X1   g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n265), .A2(G45), .ZN(new_n493));
  OAI211_X1 g0293(.A(G270), .B(new_n293), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n495), .B1(new_n283), .B2(new_n479), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n466), .A2(new_n469), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n466), .A2(KEYINPUT20), .A3(new_n469), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n430), .A2(new_n465), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n262), .A2(new_n409), .A3(new_n473), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT86), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n496), .A2(new_n504), .A3(new_n505), .A4(G179), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n480), .A2(new_n486), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT21), .A4(G169), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n488), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT87), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT87), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n488), .A2(new_n506), .A3(new_n511), .A4(new_n508), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n504), .A2(new_n507), .A3(G169), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(KEYINPUT21), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n504), .B1(G200), .B2(new_n507), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n306), .B2(new_n507), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n510), .A2(new_n512), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G244), .B(new_n448), .C1(new_n323), .C2(new_n324), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g0321(.A1(KEYINPUT4), .A2(G244), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n279), .A2(new_n448), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n521), .A2(new_n467), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT81), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n279), .A2(KEYINPUT81), .A3(G250), .A4(G1698), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n293), .B1(new_n524), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G257), .B(new_n293), .C1(new_n492), .C2(new_n493), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n489), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(KEYINPUT82), .B(G200), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT82), .ZN(new_n534));
  INV_X1    g0334(.A(new_n467), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n276), .B2(new_n522), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n521), .A3(new_n527), .A4(new_n528), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n532), .B1(new_n537), .B2(new_n283), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n534), .B1(new_n538), .B2(new_n364), .ZN(new_n539));
  OAI21_X1  g0339(.A(G107), .B1(new_n326), .B2(new_n328), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  AND2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(new_n205), .ZN(new_n543));
  INV_X1    g0343(.A(G107), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n544), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(G20), .B1(G77), .B2(new_n243), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n262), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n265), .A2(G33), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n262), .A2(new_n266), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(new_n468), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n266), .A2(G97), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n548), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n538), .A2(G190), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n533), .A2(new_n539), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n254), .B(G87), .C1(new_n323), .C2(new_n324), .ZN(new_n556));
  AND2_X1   g0356(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n557));
  NOR2_X1   g0357(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n279), .A2(new_n254), .A3(G87), .A4(new_n557), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT89), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n562), .B(KEYINPUT23), .C1(new_n254), .C2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n254), .A2(G33), .A3(G116), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT23), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n544), .A3(G20), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT23), .B1(new_n254), .B2(G107), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT89), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n560), .A2(new_n561), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT24), .ZN(new_n571));
  AND4_X1   g0371(.A1(new_n569), .A2(new_n563), .A3(new_n564), .A4(new_n566), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT24), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(new_n561), .A4(new_n560), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n262), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n266), .A2(G107), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n576), .B(KEYINPUT25), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n550), .B2(new_n544), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G257), .B(G1698), .C1(new_n323), .C2(new_n324), .ZN(new_n580));
  OAI211_X1 g0380(.A(G250), .B(new_n448), .C1(new_n323), .C2(new_n324), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G294), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n283), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT90), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(KEYINPUT90), .A3(new_n283), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n483), .A2(G264), .B1(new_n485), .B2(new_n481), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n586), .A2(new_n306), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n483), .A2(G264), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n584), .A2(new_n489), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n364), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n579), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n537), .A2(new_n283), .ZN(new_n595));
  INV_X1    g0395(.A(new_n532), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n301), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n540), .A2(new_n547), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n263), .ZN(new_n600));
  INV_X1    g0400(.A(new_n551), .ZN(new_n601));
  INV_X1    g0401(.A(new_n552), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n538), .A2(new_n285), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n598), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n555), .A2(new_n594), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n279), .A2(new_n254), .A3(G68), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n254), .B1(new_n389), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G87), .B2(new_n206), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n608), .B1(new_n255), .B2(new_n468), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n263), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n430), .A2(new_n435), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n270), .A2(KEYINPUT85), .A3(G87), .A4(new_n549), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  INV_X1    g0417(.A(G87), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n550), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n615), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n279), .A2(G244), .A3(G1698), .ZN(new_n621));
  NAND2_X1  g0421(.A1(G33), .A2(G116), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n390), .C2(new_n451), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT83), .B1(new_n283), .B2(new_n484), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT83), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n293), .A2(new_n625), .A3(G274), .A4(new_n482), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n293), .A2(G250), .A3(new_n493), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n624), .A2(KEYINPUT84), .A3(new_n627), .A4(new_n626), .ZN(new_n631));
  AOI221_X4 g0431(.A(G190), .B1(new_n623), .B2(new_n283), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(new_n283), .ZN(new_n634));
  AOI21_X1  g0434(.A(G200), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n620), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n587), .A2(new_n588), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n301), .B1(new_n637), .B2(new_n586), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n591), .A2(new_n285), .ZN(new_n639));
  OAI22_X1  g0439(.A1(new_n638), .A2(new_n639), .B1(new_n575), .B2(new_n578), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n613), .A2(new_n614), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n550), .A2(new_n435), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n633), .A2(new_n285), .A3(new_n634), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n630), .A2(new_n631), .B1(new_n283), .B2(new_n623), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n643), .B(new_n644), .C1(G169), .C2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n636), .A2(new_n640), .A3(new_n646), .ZN(new_n647));
  NOR4_X1   g0447(.A1(new_n464), .A2(new_n518), .A3(new_n606), .A4(new_n647), .ZN(G372));
  INV_X1    g0448(.A(new_n464), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n645), .A2(new_n285), .B1(new_n641), .B2(new_n642), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n633), .A2(new_n634), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT91), .B1(new_n651), .B2(new_n301), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT91), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n645), .A2(new_n653), .A3(G169), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n650), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n636), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n606), .ZN(new_n658));
  INV_X1    g0458(.A(new_n640), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n659), .A2(new_n509), .A3(new_n514), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n656), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n598), .A2(new_n603), .A3(new_n604), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n655), .A2(new_n662), .A3(new_n636), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT26), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n645), .A2(new_n306), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(G200), .B2(new_n645), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n651), .A2(new_n301), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n667), .A2(new_n620), .B1(new_n650), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(KEYINPUT92), .A3(KEYINPUT26), .A4(new_n662), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n662), .A2(new_n636), .A3(KEYINPUT26), .A4(new_n646), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT92), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n665), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n661), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n649), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n303), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n379), .A2(new_n383), .ZN(new_n678));
  INV_X1    g0478(.A(new_n457), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n679), .A2(new_n455), .B1(G169), .B2(new_n453), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n443), .B2(new_n444), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n426), .A2(new_n415), .B1(new_n681), .B2(new_n418), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n366), .A2(new_n385), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n678), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n309), .A2(new_n310), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n677), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n676), .A2(new_n687), .ZN(G369));
  NAND2_X1  g0488(.A1(new_n405), .A2(new_n254), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n691), .A3(G213), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n475), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n509), .B2(new_n514), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n518), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g0498(.A(KEYINPUT93), .B(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n694), .B1(new_n575), .B2(new_n578), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n594), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n640), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n640), .A2(new_n694), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n702), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n514), .B1(new_n509), .B2(KEYINPUT87), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n694), .B1(new_n711), .B2(new_n512), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n706), .B1(new_n712), .B2(new_n705), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n215), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n209), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n510), .A2(new_n512), .A3(new_n515), .A4(new_n640), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n555), .A2(new_n594), .A3(new_n605), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n651), .A2(KEYINPUT91), .A3(new_n301), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n653), .B1(new_n645), .B2(G169), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n727), .A2(new_n650), .B1(new_n667), .B2(new_n620), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n723), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n662), .A2(new_n636), .A3(new_n664), .A4(new_n646), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n729), .A2(new_n730), .A3(new_n655), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n722), .B1(new_n732), .B2(new_n695), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR4_X1   g0534(.A1(new_n518), .A2(new_n606), .A3(new_n647), .A4(new_n694), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n480), .A2(new_n486), .A3(G179), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n584), .A2(new_n590), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n645), .A2(new_n736), .A3(new_n738), .A4(new_n538), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n487), .A2(new_n737), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT30), .A3(new_n538), .A4(new_n645), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n496), .A2(G179), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n651), .A3(new_n591), .A4(new_n597), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n694), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT31), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n700), .B1(new_n735), .B2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT94), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n675), .A2(new_n722), .A3(new_n695), .ZN(new_n755));
  AND3_X1   g0555(.A1(new_n636), .A2(new_n640), .A3(new_n646), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n724), .A2(new_n756), .A3(new_n695), .ZN(new_n757));
  OAI211_X1 g0557(.A(new_n749), .B(new_n750), .C1(new_n757), .C2(new_n518), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(KEYINPUT94), .A3(new_n700), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n734), .A2(new_n754), .A3(new_n755), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n721), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n404), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n265), .B1(new_n763), .B2(G45), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n717), .A2(KEYINPUT95), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT95), .ZN(new_n766));
  INV_X1    g0566(.A(new_n764), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n716), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G355), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n279), .A2(new_n215), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n771), .A2(new_n772), .B1(G116), .B2(new_n215), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n238), .A2(G45), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n715), .A2(new_n279), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AND2_X1   g0576(.A1(new_n287), .A2(new_n289), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n210), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n773), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n211), .B1(G20), .B2(new_n301), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT96), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n770), .B1(new_n779), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n254), .A2(new_n285), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(G190), .A3(new_n364), .ZN(new_n789));
  INV_X1    g0589(.A(G322), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G190), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G311), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n325), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n254), .A2(G179), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n792), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n791), .B(new_n795), .C1(G329), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n788), .A2(G200), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n306), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G326), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(G190), .ZN(new_n803));
  XNOR2_X1  g0603(.A(KEYINPUT33), .B(G317), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n796), .A2(G190), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n803), .A2(new_n804), .B1(new_n806), .B2(G303), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n796), .A2(new_n306), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n285), .A2(new_n364), .A3(G190), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G20), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n809), .A2(G283), .B1(new_n811), .B2(G294), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n799), .A2(new_n802), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n805), .A2(new_n618), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n798), .A2(G159), .ZN(new_n816));
  INV_X1    g0616(.A(new_n803), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n816), .B2(KEYINPUT32), .C1(new_n817), .C2(new_n318), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n816), .A2(KEYINPUT32), .B1(G107), .B2(new_n809), .ZN(new_n819));
  INV_X1    g0619(.A(new_n801), .ZN(new_n820));
  INV_X1    g0620(.A(new_n811), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n819), .B1(new_n264), .B2(new_n820), .C1(new_n468), .C2(new_n821), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n279), .B1(new_n793), .B2(new_n278), .C1(new_n245), .C2(new_n789), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n813), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n787), .B1(new_n825), .B2(new_n781), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n784), .B(KEYINPUT97), .Z(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n698), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n701), .A2(new_n769), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n698), .A2(new_n700), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT98), .ZN(G396));
  AOI21_X1  g0632(.A(new_n694), .B1(new_n661), .B2(new_n674), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n445), .A2(new_n694), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n459), .A2(new_n834), .A3(new_n462), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT100), .B1(new_n681), .B2(new_n694), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n445), .A2(new_n458), .A3(new_n694), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT100), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n833), .B(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n518), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n842), .A2(new_n724), .A3(new_n756), .A4(new_n695), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT31), .B1(new_n746), .B2(new_n694), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n753), .B(new_n699), .C1(new_n843), .C2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(KEYINPUT94), .B1(new_n758), .B2(new_n700), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n770), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n849), .B2(new_n841), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n781), .A2(new_n782), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(G77), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n325), .B1(new_n805), .B2(new_n544), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT99), .Z(new_n856));
  OAI22_X1  g0656(.A1(new_n793), .A2(new_n465), .B1(new_n797), .B2(new_n794), .ZN(new_n857));
  INV_X1    g0657(.A(new_n789), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(G294), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n803), .A2(G283), .B1(G97), .B2(new_n811), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n801), .A2(G303), .B1(new_n809), .B2(G87), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n856), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n279), .B1(new_n797), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n809), .A2(G68), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n264), .B2(new_n805), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n864), .B(new_n866), .C1(G58), .C2(new_n811), .ZN(new_n867));
  INV_X1    g0667(.A(new_n793), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n858), .A2(G143), .B1(new_n868), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(G150), .ZN(new_n870));
  INV_X1    g0670(.A(G137), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n869), .B1(new_n817), .B2(new_n870), .C1(new_n871), .C2(new_n820), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT34), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n862), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n769), .B(new_n854), .C1(new_n877), .C2(new_n781), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n878), .B1(new_n840), .B2(new_n783), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n851), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n763), .A2(new_n265), .ZN(new_n882));
  XNOR2_X1  g0682(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n341), .A2(new_n382), .ZN(new_n884));
  INV_X1    g0684(.A(new_n692), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n341), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n375), .A2(new_n384), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n884), .A2(new_n886), .A3(new_n887), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n386), .A2(new_n341), .A3(new_n885), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n883), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n369), .B1(new_n335), .B2(new_n322), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n339), .A3(new_n263), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n692), .B1(new_n317), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n386), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n341), .A2(new_n365), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n378), .A2(new_n692), .B1(new_n317), .B2(new_n896), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n891), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n386), .A2(new_n897), .B1(new_n901), .B2(new_n891), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(KEYINPUT104), .A3(KEYINPUT38), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n894), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n426), .A2(new_n415), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n415), .A2(new_n694), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n418), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n415), .B(new_n694), .C1(new_n426), .C2(new_n419), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n758), .A3(new_n840), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT40), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n898), .B2(new_n902), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT40), .B1(new_n917), .B2(new_n903), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n918), .A2(new_n758), .A3(new_n840), .A4(new_n913), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT105), .Z(new_n921));
  INV_X1    g0721(.A(new_n758), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n464), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n699), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n923), .B2(new_n921), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n902), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT39), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n926), .A2(new_n916), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n892), .A2(new_n893), .ZN(new_n929));
  INV_X1    g0729(.A(new_n883), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT104), .B1(new_n906), .B2(KEYINPUT38), .ZN(new_n932));
  AND4_X1   g0732(.A1(KEYINPUT104), .A2(new_n898), .A3(KEYINPUT38), .A4(new_n902), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n928), .B1(new_n934), .B2(new_n927), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n909), .A2(new_n694), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n675), .A2(new_n840), .A3(new_n695), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n681), .A2(new_n695), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n940), .B(new_n913), .C1(new_n926), .C2(new_n916), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n678), .A2(new_n885), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n733), .B1(new_n722), .B2(new_n833), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(new_n464), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n687), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n943), .B(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n882), .B1(new_n925), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n925), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n211), .A2(new_n254), .A3(new_n465), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n546), .B(KEYINPUT101), .Z(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT35), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  XNOR2_X1  g0755(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n201), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n318), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n209), .A2(new_n278), .A3(new_n319), .ZN(new_n960));
  OAI211_X1 g0760(.A(G1), .B(new_n404), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n949), .A2(new_n957), .A3(new_n961), .ZN(G367));
  INV_X1    g0762(.A(new_n435), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n786), .B1(new_n715), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n229), .A2(new_n775), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n769), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(G317), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n325), .B1(new_n797), .B2(new_n967), .C1(new_n789), .C2(new_n478), .ZN(new_n968));
  INV_X1    g0768(.A(G294), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n817), .A2(new_n969), .B1(new_n468), .B2(new_n808), .ZN(new_n970));
  AOI211_X1 g0770(.A(new_n968), .B(new_n970), .C1(G311), .C2(new_n801), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n868), .A2(G283), .B1(G107), .B2(new_n811), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT111), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n806), .A2(G116), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(KEYINPUT111), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n971), .A2(new_n973), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT112), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n809), .A2(G77), .ZN(new_n980));
  INV_X1    g0780(.A(G159), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n980), .B1(new_n245), .B2(new_n805), .C1(new_n817), .C2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(G143), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n820), .A2(new_n983), .B1(new_n318), .B2(new_n821), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n279), .B1(new_n793), .B2(new_n201), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n789), .A2(new_n870), .B1(new_n797), .B2(new_n871), .ZN(new_n986));
  OR4_X1    g0786(.A1(new_n982), .A2(new_n984), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n977), .A2(new_n978), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n979), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT47), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n781), .B1(new_n989), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n966), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n827), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n620), .A2(new_n695), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n655), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n728), .B2(new_n995), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT106), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n993), .B1(new_n994), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT108), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n712), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n708), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n510), .A2(new_n512), .A3(new_n515), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n594), .A2(new_n703), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1004), .A2(new_n640), .A3(new_n695), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n702), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n701), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1001), .B1(new_n760), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n944), .A2(new_n849), .A3(KEYINPUT108), .A4(new_n1010), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT44), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n555), .B(new_n605), .C1(new_n553), .C2(new_n695), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT107), .B1(new_n662), .B2(new_n694), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT107), .ZN(new_n1017));
  NOR3_X1   g0817(.A1(new_n605), .A2(new_n1017), .A3(new_n695), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1014), .B1(new_n713), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1006), .A2(new_n707), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1019), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(KEYINPUT44), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1006), .A2(new_n1019), .A3(new_n707), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n713), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AND3_X1   g0829(.A1(new_n1024), .A2(new_n1029), .A3(new_n710), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n710), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1012), .A2(new_n1013), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT109), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1012), .A2(new_n1032), .A3(KEYINPUT109), .A4(new_n1013), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n761), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n716), .B(KEYINPUT41), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(KEYINPUT110), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT110), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n760), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1042), .B1(new_n1043), .B2(new_n1039), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n767), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n709), .A2(new_n712), .A3(new_n1019), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT42), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n662), .B1(new_n1019), .B2(new_n659), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n1048), .B2(new_n694), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1046), .A2(KEYINPUT42), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT43), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1049), .A2(new_n1050), .B1(new_n1051), .B2(new_n998), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n998), .A2(new_n1051), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n710), .A2(new_n1022), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1000), .B1(new_n1045), .B2(new_n1056), .ZN(G387));
  NAND2_X1  g0857(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n716), .C1(new_n761), .C2(new_n1010), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n772), .A2(new_n718), .B1(G107), .B2(new_n215), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n718), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n286), .B1(new_n318), .B2(new_n278), .C1(new_n1061), .C2(KEYINPUT113), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(KEYINPUT113), .B2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n433), .A2(G50), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n777), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n776), .B1(new_n234), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1060), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n770), .B1(new_n1069), .B2(new_n786), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n963), .A2(new_n811), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n264), .B2(new_n789), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT114), .Z(new_n1073));
  OAI221_X1 g0873(.A(new_n279), .B1(new_n797), .B2(new_n870), .C1(new_n318), .C2(new_n793), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n315), .B2(new_n803), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n808), .A2(new_n468), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n805), .A2(new_n278), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(G159), .C2(new_n801), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1073), .A2(new_n1075), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(G283), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n821), .A2(new_n1080), .B1(new_n805), .B2(new_n969), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n858), .A2(G317), .B1(new_n868), .B2(G303), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n817), .B2(new_n794), .C1(new_n790), .C2(new_n820), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT48), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT49), .ZN(new_n1087));
  AND2_X1   g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n279), .B1(new_n798), .B2(G326), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n465), .B2(new_n808), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT115), .Z(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1079), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1070), .B1(new_n1093), .B2(new_n781), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n709), .B2(new_n827), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT116), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1059), .B(new_n1096), .C1(new_n764), .C2(new_n1011), .ZN(G393));
  INV_X1    g0897(.A(new_n1032), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n717), .B1(new_n1058), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1037), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1022), .A2(new_n784), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n785), .B1(new_n468), .B2(new_n215), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n241), .A2(new_n776), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n770), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n817), .A2(new_n478), .B1(new_n465), .B2(new_n821), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n325), .B1(new_n797), .B2(new_n790), .C1(new_n969), .C2(new_n793), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n544), .A2(new_n808), .B1(new_n805), .B2(new_n1080), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G317), .A2(new_n801), .B1(new_n858), .B2(G311), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT52), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G150), .A2(new_n801), .B1(new_n858), .B2(G159), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT51), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n821), .A2(new_n278), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(G68), .B2(new_n806), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n279), .B1(new_n797), .B2(new_n983), .C1(new_n433), .C2(new_n793), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n803), .A2(new_n958), .B1(new_n809), .B2(G87), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1108), .A2(new_n1110), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1104), .B1(new_n1119), .B2(new_n781), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1032), .A2(new_n767), .B1(new_n1101), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1100), .A2(new_n1121), .ZN(G390));
  INV_X1    g0922(.A(new_n936), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n939), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n833), .B2(new_n840), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n913), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n917), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n908), .B2(KEYINPUT39), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n732), .A2(new_n695), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n681), .A2(KEYINPUT100), .A3(new_n694), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n837), .A2(new_n838), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n463), .A2(new_n834), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n939), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n913), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n905), .A2(new_n907), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n936), .B1(new_n1136), .B2(new_n931), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1127), .A2(new_n1129), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n840), .B(new_n913), .C1(new_n847), .C2(new_n848), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(KEYINPUT117), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n754), .A2(new_n759), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT117), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n840), .A4(new_n913), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT118), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1138), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n731), .A2(new_n655), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(KEYINPUT26), .B2(new_n663), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n694), .B1(new_n1148), .B2(new_n729), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1124), .B1(new_n1149), .B2(new_n840), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n934), .B(new_n1123), .C1(new_n1150), .C2(new_n1126), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n936), .B1(new_n940), .B2(new_n913), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n935), .ZN(new_n1153));
  AND4_X1   g0953(.A1(G330), .A2(new_n913), .A3(new_n758), .A4(new_n840), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1146), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1145), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n767), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n770), .B1(new_n853), .B2(new_n315), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n806), .A2(G150), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT53), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n279), .B1(new_n797), .B2(new_n1163), .C1(new_n793), .C2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n817), .A2(new_n871), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n821), .A2(new_n981), .B1(new_n808), .B2(new_n201), .ZN(new_n1167));
  OR4_X1    g0967(.A1(new_n1162), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G128), .A2(new_n801), .B1(new_n858), .B2(G132), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT121), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1113), .B1(G283), .B2(new_n801), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n544), .B2(new_n817), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n789), .A2(new_n465), .B1(new_n797), .B2(new_n969), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n279), .B(new_n1173), .C1(G97), .C2(new_n868), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n815), .A3(new_n865), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1168), .A2(new_n1170), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1160), .B1(new_n1176), .B2(new_n781), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n935), .B2(new_n783), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1159), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n758), .A2(G330), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n649), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n945), .A2(new_n1182), .A3(new_n687), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT119), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n840), .B1(new_n847), .B2(new_n848), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1154), .B1(new_n1185), .B2(new_n1126), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1186), .B2(new_n1125), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1181), .A2(new_n840), .A3(new_n913), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1133), .B1(new_n754), .B2(new_n759), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1189), .B2(new_n913), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1190), .A2(KEYINPUT119), .A3(new_n940), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1181), .A2(new_n840), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1134), .B1(new_n1193), .B2(new_n1126), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1144), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1183), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(KEYINPUT118), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1146), .A2(new_n1155), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1187), .A2(new_n1191), .B1(new_n1144), .B2(new_n1194), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n1157), .A2(new_n1156), .B1(new_n1201), .B2(new_n1183), .ZN(new_n1202));
  AND4_X1   g1002(.A1(KEYINPUT120), .A2(new_n1200), .A3(new_n716), .A4(new_n1202), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1186), .A2(new_n1184), .A3(new_n1125), .ZN(new_n1204));
  AOI21_X1  g1004(.A(KEYINPUT119), .B1(new_n1190), .B2(new_n940), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1195), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1183), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1198), .A2(new_n1155), .A3(new_n1146), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n717), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT120), .B1(new_n1210), .B2(new_n1200), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1180), .B1(new_n1203), .B2(new_n1211), .ZN(G378));
  NAND3_X1  g1012(.A1(new_n311), .A2(new_n273), .A3(new_n885), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n273), .A2(new_n885), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n303), .B(new_n1214), .C1(new_n309), .C2(new_n310), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1213), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1213), .B2(new_n1215), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n920), .A2(new_n1219), .A3(G330), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1219), .B1(new_n920), .B2(G330), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n943), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n920), .A2(G330), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1219), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n937), .A2(new_n941), .A3(new_n942), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1227), .A3(new_n1220), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1223), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(new_n782), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n770), .B1(new_n853), .B2(new_n958), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G33), .A2(G41), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G50), .B(new_n1232), .C1(new_n325), .C2(new_n290), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n817), .A2(new_n468), .B1(new_n245), .B2(new_n808), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G116), .B2(new_n801), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G41), .B(new_n279), .C1(new_n798), .C2(G283), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n858), .A2(G107), .B1(new_n868), .B2(new_n963), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1077), .B1(G68), .B2(new_n811), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1164), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n806), .A2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT122), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n801), .A2(G125), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n858), .A2(G128), .B1(new_n868), .B2(G137), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n803), .A2(G132), .B1(G150), .B2(new_n811), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT59), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n809), .A2(G159), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT123), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1251), .A2(G124), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(G124), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n798), .A2(new_n1252), .A3(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1249), .A2(new_n1250), .A3(new_n1254), .A4(new_n1232), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1248), .A2(KEYINPUT59), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1241), .B1(new_n1240), .B2(new_n1239), .C1(new_n1255), .C2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1231), .B1(new_n1257), .B2(new_n781), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1229), .A2(new_n767), .B1(new_n1230), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1183), .B1(new_n1158), .B2(new_n1196), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n1221), .A2(new_n1222), .A3(new_n943), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1227), .B1(new_n1226), .B2(new_n1220), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT57), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n716), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1207), .B1(new_n1209), .B2(new_n1201), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT57), .B1(new_n1265), .B2(new_n1229), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1259), .B1(new_n1264), .B2(new_n1266), .ZN(G375));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n1201), .B2(new_n764), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1206), .A2(KEYINPUT124), .A3(new_n767), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n770), .B1(new_n853), .B2(G68), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n817), .A2(new_n465), .B1(new_n820), .B2(new_n969), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G97), .B2(new_n806), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n789), .A2(new_n1080), .B1(new_n793), .B2(new_n544), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n279), .B(new_n1274), .C1(G303), .C2(new_n798), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1273), .A2(new_n980), .A3(new_n1071), .A4(new_n1275), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n821), .A2(new_n264), .B1(new_n805), .B2(new_n981), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G132), .B2(new_n801), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n325), .B1(new_n798), .B2(G128), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n858), .A2(G137), .B1(new_n868), .B2(G150), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n803), .A2(new_n1242), .B1(new_n809), .B2(G58), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1278), .A2(new_n1279), .A3(new_n1280), .A4(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1276), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1271), .B1(new_n1283), .B2(new_n781), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n913), .B2(new_n783), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1269), .A2(new_n1270), .A3(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1192), .A2(new_n1183), .A3(new_n1195), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1208), .A2(new_n1040), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(G381));
  NOR2_X1   g1089(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1202), .A2(new_n716), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1180), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G390), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1286), .A2(new_n1293), .A3(new_n1294), .A4(new_n1288), .ZN(new_n1295));
  OR4_X1    g1095(.A1(G387), .A2(G375), .A3(new_n1292), .A4(new_n1295), .ZN(G407));
  NAND2_X1  g1096(.A1(new_n1230), .A2(new_n1258), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1229), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1298), .B2(new_n764), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT57), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1260), .B2(new_n1298), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1300), .B1(new_n1223), .B2(new_n1228), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n717), .B1(new_n1265), .B2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1299), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1179), .B1(new_n1200), .B2(new_n1210), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1304), .A2(new_n693), .A3(new_n1305), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(G407), .A2(G213), .A3(new_n1306), .ZN(G409));
  NAND3_X1  g1107(.A1(new_n1265), .A2(new_n1040), .A3(new_n1229), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1259), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT120), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1291), .B2(new_n1290), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1210), .A2(KEYINPUT120), .A3(new_n1200), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1179), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1310), .B1(new_n1314), .B2(G375), .ZN(new_n1315));
  INV_X1    g1115(.A(G213), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1316), .A2(G343), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT125), .B1(new_n1287), .B2(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1196), .A2(new_n717), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT125), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1201), .A2(new_n1322), .A3(KEYINPUT60), .A4(new_n1183), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1287), .A2(new_n1319), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(new_n1321), .A3(new_n1323), .A4(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1325), .A2(G384), .A3(new_n1286), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(G384), .B1(new_n1325), .B2(new_n1286), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1315), .A2(new_n1318), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT61), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1315), .A2(new_n1333), .A3(new_n1318), .A4(new_n1329), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1325), .A2(new_n1286), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n880), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1317), .A2(G2897), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1336), .A2(new_n1326), .A3(new_n1337), .ZN(new_n1338));
  OAI211_X1 g1138(.A(G2897), .B(new_n1317), .C1(new_n1327), .C2(new_n1328), .ZN(new_n1339));
  AOI22_X1  g1139(.A1(G378), .A2(new_n1304), .B1(new_n1305), .B2(new_n1309), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1338), .B(new_n1339), .C1(new_n1340), .C2(new_n1317), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1331), .A2(new_n1332), .A3(new_n1334), .A4(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G387), .A2(new_n1293), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT126), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1000), .B(G390), .C1(new_n1045), .C2(new_n1056), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(G393), .B(G396), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1343), .A2(new_n1344), .A3(new_n1345), .A4(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1345), .A2(KEYINPUT126), .ZN(new_n1349));
  AOI22_X1  g1149(.A1(new_n1349), .A2(new_n1346), .B1(new_n1343), .B2(new_n1345), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1348), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1342), .A2(new_n1351), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1339), .A2(new_n1338), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1315), .A2(new_n1318), .ZN(new_n1354));
  AOI21_X1  g1154(.A(KEYINPUT61), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1349), .A2(new_n1346), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1347), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT63), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1330), .A2(new_n1360), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1318), .A4(new_n1329), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1355), .A2(new_n1359), .A3(new_n1361), .A4(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1352), .A2(new_n1363), .ZN(G405));
  NAND2_X1  g1164(.A1(G378), .A2(new_n1304), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(G375), .A2(new_n1305), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1336), .A2(new_n1326), .ZN(new_n1367));
  AND3_X1   g1167(.A1(new_n1365), .A2(new_n1366), .A3(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(new_n1367), .B1(new_n1365), .B2(new_n1366), .ZN(new_n1369));
  OAI22_X1  g1169(.A1(new_n1348), .A2(new_n1350), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1314), .A2(G375), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1304), .A2(new_n1292), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1329), .B1(new_n1371), .B2(new_n1372), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1365), .A2(new_n1366), .A3(new_n1367), .ZN(new_n1374));
  NAND4_X1  g1174(.A1(new_n1358), .A2(new_n1373), .A3(new_n1347), .A4(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT127), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1370), .B1(new_n1375), .B2(new_n1376), .ZN(new_n1377));
  NOR2_X1   g1177(.A1(new_n1368), .A2(new_n1369), .ZN(new_n1378));
  AOI21_X1  g1178(.A(KEYINPUT127), .B1(new_n1351), .B2(new_n1378), .ZN(new_n1379));
  NOR2_X1   g1179(.A1(new_n1377), .A2(new_n1379), .ZN(G402));
endmodule


