//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT78), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  OAI21_X1  g003(.A(G221), .B1(new_n189), .B2(G902), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G469), .ZN(new_n192));
  INV_X1    g006(.A(G902), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .A4(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OR2_X1    g019(.A1(KEYINPUT80), .A2(G104), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT80), .A2(G104), .ZN(new_n207));
  AOI21_X1  g021(.A(G107), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(G101), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n209), .A3(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n208), .B2(new_n212), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(G107), .A3(new_n207), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n205), .B(new_n211), .C1(new_n214), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT69), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n199), .B2(new_n204), .ZN(new_n220));
  AOI21_X1  g034(.A(G128), .B1(new_n200), .B2(new_n201), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n202), .A2(new_n197), .A3(G143), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(KEYINPUT69), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n203), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n213), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT80), .A2(G104), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT80), .A2(G104), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n209), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n215), .A2(new_n216), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n228), .B1(G104), .B2(new_n209), .ZN(new_n231));
  AOI22_X1  g045(.A1(new_n229), .A2(new_n230), .B1(new_n231), .B2(G101), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n218), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  INV_X1    g048(.A(G134), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G137), .ZN(new_n236));
  AOI21_X1  g050(.A(G131), .B1(new_n235), .B2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT66), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(new_n237), .A3(new_n242), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n236), .B(new_n239), .C1(G134), .C2(new_n238), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n233), .A2(KEYINPUT12), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT12), .B1(new_n233), .B2(new_n247), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n200), .A2(new_n201), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR3_X1   g066(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(G143), .B(G146), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT0), .A3(G128), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n215), .B(new_n213), .C1(new_n208), .C2(new_n212), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n262));
  OR2_X1    g076(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(KEYINPUT4), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n216), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n214), .B2(new_n217), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n216), .B1(new_n229), .B2(new_n215), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n260), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n224), .A2(KEYINPUT10), .A3(new_n232), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n241), .A2(new_n243), .B1(G131), .B2(new_n245), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT10), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n218), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n269), .A2(new_n270), .A3(new_n271), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(G953), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G227), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT79), .ZN(new_n277));
  XNOR2_X1  g091(.A(G110), .B(G140), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n250), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n269), .A2(new_n270), .A3(new_n273), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n247), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n279), .B1(new_n283), .B2(new_n274), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n192), .B(new_n193), .C1(new_n281), .C2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT82), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n279), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT69), .B1(new_n221), .B2(new_n222), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n204), .B(new_n219), .C1(new_n257), .C2(G128), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n272), .B1(new_n291), .B2(new_n203), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n292), .A2(new_n232), .B1(new_n272), .B2(new_n218), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n271), .B1(new_n293), .B2(new_n269), .ZN(new_n294));
  AND4_X1   g108(.A1(new_n271), .A2(new_n269), .A3(new_n270), .A4(new_n273), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n274), .B(new_n279), .C1(new_n248), .C2(new_n249), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT82), .A3(new_n192), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n280), .A2(new_n294), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n274), .B1(new_n248), .B2(new_n249), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n288), .ZN(new_n303));
  OAI21_X1  g117(.A(G469), .B1(new_n303), .B2(G902), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n191), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n275), .A2(G952), .ZN(new_n307));
  NAND2_X1  g121(.A1(G234), .A2(G237), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(G902), .A3(G953), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT21), .B(G898), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G125), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n291), .A2(new_n316), .A3(new_n203), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n259), .A2(G125), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n317), .B2(new_n319), .ZN(new_n321));
  INV_X1    g135(.A(G224), .ZN(new_n322));
  OAI22_X1  g136(.A1(new_n320), .A2(new_n321), .B1(new_n322), .B2(G953), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT84), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n322), .A2(G953), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n230), .A2(new_n229), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT70), .ZN(new_n331));
  INV_X1    g145(.A(G119), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G116), .ZN(new_n333));
  INV_X1    g147(.A(G116), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G119), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT2), .B(G113), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G113), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT2), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT2), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G113), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G116), .B(G119), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT70), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n338), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT83), .B1(new_n333), .B2(KEYINPUT5), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n333), .A2(new_n335), .A3(KEYINPUT5), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n332), .A4(G116), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n348), .A3(G113), .A4(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n330), .A2(new_n346), .A3(new_n211), .A4(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n267), .A2(new_n268), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n336), .A2(new_n337), .ZN(new_n355));
  NOR3_X1   g169(.A1(new_n336), .A2(new_n337), .A3(new_n331), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT70), .B1(new_n343), .B2(new_n344), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n266), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n353), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(G110), .B(G122), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n361), .B(new_n353), .C1(new_n354), .C2(new_n359), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(KEYINPUT6), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n366), .A3(new_n362), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n329), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n361), .B(KEYINPUT8), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n211), .B1(new_n214), .B2(new_n217), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n330), .A2(new_n211), .B1(new_n346), .B2(new_n352), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n369), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT7), .B1(new_n322), .B2(G953), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n317), .A2(new_n319), .A3(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n364), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT85), .B1(new_n324), .B2(new_n375), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n380));
  AOI211_X1 g194(.A(new_n380), .B(new_n376), .C1(new_n317), .C2(new_n319), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G210), .B1(G237), .B2(G902), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n368), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n384), .B1(new_n368), .B2(new_n383), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n306), .B(new_n315), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G125), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n316), .A2(G140), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT16), .ZN(new_n391));
  OR3_X1    g205(.A1(new_n316), .A2(KEYINPUT16), .A3(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n197), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n392), .A3(G146), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(KEYINPUT74), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT74), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n397), .A3(new_n197), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(G237), .A2(G953), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(G143), .A3(G214), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(G143), .B1(new_n400), .B2(G214), .ZN(new_n403));
  OAI211_X1 g217(.A(KEYINPUT17), .B(G131), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT88), .ZN(new_n405));
  INV_X1    g219(.A(G131), .ZN(new_n406));
  INV_X1    g220(.A(G237), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(new_n275), .A3(G214), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n195), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n409), .B2(new_n401), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n410), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT17), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n406), .A3(new_n401), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n399), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  XOR2_X1   g232(.A(G113), .B(G122), .Z(new_n419));
  XOR2_X1   g233(.A(KEYINPUT87), .B(G104), .Z(new_n420));
  XOR2_X1   g234(.A(new_n419), .B(new_n420), .Z(new_n421));
  NAND2_X1  g235(.A1(new_n409), .A2(new_n401), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT18), .A2(G131), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n389), .A2(new_n390), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT86), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n389), .A2(new_n390), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(G146), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n389), .A2(new_n390), .A3(new_n197), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n418), .A2(new_n421), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n414), .A2(new_n416), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n426), .A2(KEYINPUT19), .A3(new_n428), .ZN(new_n435));
  OR2_X1    g249(.A1(new_n425), .A2(KEYINPUT19), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n197), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n437), .A3(new_n395), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n432), .ZN(new_n439));
  INV_X1    g253(.A(new_n421), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT20), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n433), .A2(new_n441), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(new_n443), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n418), .A2(new_n421), .A3(new_n432), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n421), .B1(new_n418), .B2(new_n432), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n193), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n445), .A2(new_n448), .B1(G475), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n334), .A2(G122), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT90), .B1(new_n453), .B2(KEYINPUT14), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT90), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT14), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n334), .A4(G122), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G116), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(KEYINPUT14), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n454), .A2(new_n457), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G107), .ZN(new_n462));
  XNOR2_X1  g276(.A(G128), .B(G143), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n235), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n453), .A2(new_n459), .A3(new_n209), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n463), .A2(KEYINPUT13), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n195), .A2(G128), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n467), .B(G134), .C1(KEYINPUT13), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n453), .A2(new_n459), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G107), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  INV_X1    g286(.A(new_n463), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT89), .B1(new_n473), .B2(G134), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n463), .A2(new_n475), .A3(new_n235), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n469), .A2(new_n472), .A3(new_n474), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n275), .A2(G217), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n189), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n466), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n466), .B2(new_n477), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n193), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G478), .ZN(new_n483));
  NOR2_X1   g297(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n482), .B(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n452), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n387), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n238), .A2(G134), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n235), .A2(G137), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT68), .B(G131), .C1(new_n492), .C2(new_n493), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n496), .A2(new_n497), .B1(new_n241), .B2(new_n243), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n224), .A2(new_n498), .B1(new_n247), .B2(new_n260), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT28), .ZN(new_n500));
  INV_X1    g314(.A(new_n358), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n497), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n244), .ZN(new_n504));
  INV_X1    g318(.A(new_n203), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(new_n289), .B2(new_n290), .ZN(new_n506));
  OAI22_X1  g320(.A1(new_n504), .A2(new_n506), .B1(new_n271), .B2(new_n259), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT28), .B1(new_n507), .B2(new_n358), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n358), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n400), .A2(G210), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(KEYINPUT27), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(G101), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n514), .A2(KEYINPUT29), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n509), .A2(KEYINPUT71), .A3(new_n510), .A4(new_n515), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n193), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n507), .A2(KEYINPUT28), .A3(new_n358), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n247), .A2(new_n523), .A3(new_n260), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT67), .B1(new_n271), .B2(new_n259), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n524), .A2(new_n525), .B1(new_n224), .B2(new_n498), .ZN(new_n526));
  OAI22_X1  g340(.A1(new_n521), .A2(new_n522), .B1(new_n501), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n514), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n514), .B1(new_n499), .B2(new_n501), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n524), .A2(new_n525), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n224), .A2(new_n498), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n358), .B1(new_n507), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n529), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT29), .B1(new_n528), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(G472), .B1(new_n520), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n514), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n527), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n499), .B2(new_n501), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n533), .B2(new_n535), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT31), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT31), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n541), .C1(new_n533), .C2(new_n535), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n540), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT32), .ZN(new_n547));
  NOR2_X1   g361(.A1(G472), .A2(G902), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n538), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n275), .A2(G221), .A3(G234), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT76), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n332), .A2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n194), .A2(G119), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT24), .B(G110), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT73), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n332), .B2(G128), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT23), .A3(new_n556), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT23), .B1(new_n194), .B2(G119), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT73), .B1(new_n194), .B2(G119), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n561), .A2(new_n563), .B1(new_n570), .B2(G110), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n396), .A3(new_n398), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n571), .A2(new_n396), .A3(KEYINPUT75), .A4(new_n398), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n395), .A2(new_n430), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n570), .A2(G110), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n562), .B1(new_n559), .B2(new_n560), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n555), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n555), .ZN(new_n583));
  AOI211_X1 g397(.A(new_n580), .B(new_n583), .C1(new_n574), .C2(new_n575), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G217), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(G234), .B2(new_n193), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n587), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n193), .B1(new_n582), .B2(new_n584), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT25), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(KEYINPUT77), .A3(KEYINPUT25), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n590), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n305), .A2(new_n491), .A3(new_n551), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NAND2_X1  g413(.A1(new_n546), .A2(new_n193), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(G472), .B1(new_n548), .B2(new_n546), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n305), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n368), .A2(new_n383), .ZN(new_n604));
  INV_X1    g418(.A(new_n384), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n368), .A2(new_n383), .A3(new_n384), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n603), .B1(new_n608), .B2(new_n306), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n603), .B(new_n306), .C1(new_n385), .C2(new_n386), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n445), .A2(new_n448), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n451), .A2(G475), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT93), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT33), .B1(new_n480), .B2(new_n481), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n466), .A2(new_n477), .ZN(new_n617));
  INV_X1    g431(.A(new_n479), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n466), .A2(new_n477), .A3(new_n479), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n616), .A2(new_n622), .A3(G478), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n483), .B(new_n193), .C1(new_n480), .C2(new_n481), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n483), .A2(new_n193), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n615), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n616), .A2(new_n622), .A3(G478), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n624), .A3(KEYINPUT93), .A4(new_n626), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n613), .A2(new_n614), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n315), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n602), .A2(new_n612), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT34), .B(G104), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  AOI21_X1  g449(.A(new_n447), .B1(new_n446), .B2(new_n443), .ZN(new_n636));
  AOI211_X1 g450(.A(KEYINPUT20), .B(new_n444), .C1(new_n433), .C2(new_n441), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n614), .B(new_n488), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT94), .B1(new_n638), .B2(new_n314), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n452), .A2(new_n640), .A3(new_n315), .A4(new_n488), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n602), .A2(new_n612), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT95), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NAND2_X1  g460(.A1(new_n593), .A2(new_n594), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n596), .A3(new_n587), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n576), .A2(new_n581), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n555), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n589), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n601), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT96), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n654), .A2(new_n601), .A3(KEYINPUT96), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n657), .A2(new_n305), .A3(new_n491), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT37), .B(G110), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT97), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n659), .B(new_n661), .ZN(G12));
  OAI21_X1  g476(.A(new_n306), .B1(new_n385), .B2(new_n386), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT92), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n610), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n275), .A2(G900), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(G902), .A3(new_n308), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT98), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT98), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n309), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n452), .A2(new_n488), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n648), .B2(new_n653), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n665), .A2(new_n551), .A3(new_n305), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XOR2_X1   g488(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n670), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n305), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT40), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT40), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n677), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT101), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n608), .B(KEYINPUT38), .Z(new_n684));
  NOR2_X1   g498(.A1(new_n452), .A2(new_n489), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n306), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n684), .A2(new_n654), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n533), .A2(new_n535), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n499), .A2(new_n501), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n539), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n529), .B2(new_n510), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n549), .B2(new_n550), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT99), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n687), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n680), .A2(new_n683), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT102), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n680), .A2(new_n683), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n195), .ZN(G45));
  NAND2_X1  g516(.A1(new_n628), .A2(new_n630), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n614), .B1(new_n636), .B2(new_n637), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n704), .A3(new_n670), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n648), .B2(new_n653), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n665), .A2(new_n551), .A3(new_n305), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  INV_X1    g522(.A(new_n590), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n648), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n546), .A2(new_n548), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT32), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n710), .B1(new_n714), .B2(new_n538), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n632), .B1(new_n664), .B2(new_n610), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n296), .A2(new_n297), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n192), .B1(new_n717), .B2(new_n193), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n191), .B(new_n718), .C1(new_n287), .C2(new_n299), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n715), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  AOI21_X1  g536(.A(new_n642), .B1(new_n664), .B2(new_n610), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n715), .A3(new_n719), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  AOI21_X1  g539(.A(new_n490), .B1(new_n648), .B2(new_n653), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n551), .A3(new_n315), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n719), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT103), .B1(new_n665), .B2(new_n719), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  INV_X1    g546(.A(new_n685), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n664), .B2(new_n610), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT104), .B(G472), .Z(new_n735));
  AND2_X1   g549(.A1(new_n509), .A2(new_n510), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n543), .B(new_n545), .C1(new_n736), .C2(new_n514), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n600), .A2(new_n735), .B1(new_n548), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(new_n597), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n734), .A2(new_n739), .A3(new_n315), .A4(new_n719), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT105), .B(G122), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G24));
  INV_X1    g556(.A(new_n705), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n654), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n729), .B2(new_n730), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  AND4_X1   g561(.A1(KEYINPUT82), .A2(new_n717), .A3(new_n192), .A4(new_n193), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT82), .B1(new_n298), .B2(new_n192), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n304), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT106), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n300), .A2(new_n752), .A3(new_n304), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n606), .A2(new_n306), .A3(new_n607), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n191), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n751), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(new_n715), .A3(new_n743), .A4(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n751), .A2(new_n753), .A3(new_n755), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n551), .A2(new_n597), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(new_n705), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n761), .B1(new_n764), .B2(new_n757), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n406), .ZN(G33));
  INV_X1    g580(.A(new_n671), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n756), .A2(new_n715), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  NAND2_X1  g583(.A1(G469), .A2(G902), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n303), .A2(KEYINPUT45), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n303), .B2(KEYINPUT45), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI22_X1  g589(.A1(new_n773), .A2(new_n774), .B1(new_n287), .B2(new_n299), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n191), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n676), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n703), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(KEYINPUT43), .A3(new_n704), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n703), .B2(new_n452), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n601), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n785), .A3(new_n654), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT44), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n754), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n779), .B(new_n788), .C1(new_n787), .C2(new_n786), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  NOR4_X1   g604(.A1(new_n551), .A2(new_n597), .A3(new_n705), .A4(new_n754), .ZN(new_n791));
  XOR2_X1   g605(.A(new_n791), .B(KEYINPUT108), .Z(new_n792));
  XNOR2_X1  g606(.A(new_n777), .B(KEYINPUT47), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G140), .ZN(G42));
  INV_X1    g609(.A(new_n754), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n719), .A2(new_n310), .A3(new_n796), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n695), .A2(new_n710), .A3(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n798), .A2(new_n452), .A3(new_n780), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n784), .A2(new_n310), .A3(new_n719), .A4(new_n796), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n763), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT48), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n729), .A2(new_n730), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n739), .A2(new_n784), .A3(new_n310), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n307), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n799), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n804), .ZN(new_n807));
  INV_X1    g621(.A(new_n306), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n684), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n809), .A3(new_n719), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT115), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n810), .B(new_n812), .Z(new_n813));
  OAI21_X1  g627(.A(new_n300), .B1(new_n192), .B2(new_n298), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n190), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n796), .B(new_n807), .C1(new_n793), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n780), .A2(new_n452), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n798), .A2(KEYINPUT116), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n800), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n654), .A3(new_n738), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT116), .B1(new_n798), .B2(new_n818), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n817), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n826), .A3(KEYINPUT51), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n828));
  OAI221_X1 g642(.A(new_n806), .B1(new_n824), .B2(KEYINPUT51), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n719), .B1(new_n609), .B2(new_n611), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT103), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n665), .A2(KEYINPUT103), .A3(new_n719), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n744), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n190), .A2(new_n670), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n652), .B(new_n835), .C1(new_n595), .C2(new_n596), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n665), .A2(new_n694), .A3(new_n685), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n751), .A2(new_n753), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n673), .B(new_n707), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT109), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n673), .A2(new_n707), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n836), .A2(new_n694), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n734), .A3(new_n751), .A4(new_n753), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n746), .A2(new_n841), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n746), .A2(new_n841), .A3(KEYINPUT52), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n760), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n762), .A2(new_n763), .A3(new_n705), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n756), .A2(new_n715), .A3(new_n743), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n758), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n724), .A2(new_n740), .A3(new_n720), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n727), .B1(new_n832), .B2(new_n833), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n856), .A3(KEYINPUT112), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n715), .B(new_n719), .C1(new_n723), .C2(new_n716), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n731), .A2(new_n740), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n858), .B1(new_n860), .B2(new_n765), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n756), .A2(new_n745), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n551), .A2(new_n670), .A3(new_n796), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n305), .A2(new_n726), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n768), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n638), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n631), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n387), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n597), .A3(new_n305), .A4(new_n601), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n659), .A2(new_n598), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT111), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n658), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n305), .A2(new_n491), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT96), .B1(new_n654), .B2(new_n601), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n598), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT111), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n745), .A2(new_n756), .B1(new_n865), .B2(new_n866), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n881), .A3(new_n768), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n863), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n849), .A2(new_n862), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT113), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n849), .A2(new_n862), .A3(new_n884), .A4(KEYINPUT113), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n840), .A2(new_n845), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n724), .A2(new_n740), .A3(new_n720), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n852), .A2(new_n758), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n731), .A4(new_n761), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n880), .A2(new_n768), .A3(new_n882), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n840), .A2(new_n845), .A3(KEYINPUT52), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n892), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n863), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n887), .A2(new_n888), .A3(new_n889), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(KEYINPUT53), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n849), .A2(new_n863), .A3(new_n897), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(KEYINPUT54), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI22_X1  g719(.A1(new_n829), .A2(new_n905), .B1(G952), .B2(G953), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n695), .A2(new_n710), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n814), .A2(KEYINPUT49), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n814), .A2(KEYINPUT49), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n780), .A2(new_n191), .A3(new_n704), .A4(new_n808), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n684), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n906), .A2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n275), .A2(G952), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n887), .A2(new_n889), .A3(new_n900), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(G902), .ZN(new_n917));
  INV_X1    g731(.A(G210), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n365), .A2(new_n367), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n329), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT55), .Z(new_n922));
  AOI21_X1  g736(.A(new_n914), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n922), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n915), .B(new_n924), .C1(new_n917), .C2(new_n918), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(G51));
  INV_X1    g740(.A(new_n901), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n885), .A2(new_n886), .B1(new_n899), .B2(new_n863), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n888), .B1(new_n928), .B2(new_n889), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g744(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(new_n770), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n717), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  OR3_X1    g747(.A1(new_n917), .A2(new_n771), .A3(new_n772), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n914), .B1(new_n933), .B2(new_n934), .ZN(G54));
  AOI21_X1  g749(.A(new_n193), .B1(new_n928), .B2(new_n889), .ZN(new_n936));
  NAND2_X1  g750(.A1(KEYINPUT58), .A2(G475), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT119), .Z(new_n938));
  AND3_X1   g752(.A1(new_n936), .A2(new_n446), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n446), .B1(new_n936), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n914), .ZN(G60));
  NAND2_X1  g755(.A1(new_n616), .A2(new_n622), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n625), .B(KEYINPUT59), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n888), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n916), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(new_n901), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT120), .B1(new_n949), .B2(new_n914), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n945), .B1(new_n927), .B2(new_n929), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT120), .ZN(new_n952));
  INV_X1    g766(.A(new_n914), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n944), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n905), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n957), .A3(new_n943), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n944), .B1(new_n901), .B2(new_n904), .ZN(new_n959));
  OAI21_X1  g773(.A(KEYINPUT121), .B1(new_n959), .B2(new_n942), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n950), .A2(new_n954), .B1(new_n958), .B2(new_n960), .ZN(G63));
  INV_X1    g775(.A(KEYINPUT61), .ZN(new_n962));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT60), .Z(new_n964));
  NAND2_X1  g778(.A1(new_n916), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n585), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n953), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n965), .A2(new_n651), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n962), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n914), .B1(new_n965), .B2(new_n585), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n970), .B(KEYINPUT61), .C1(new_n651), .C2(new_n965), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(G66));
  OAI21_X1  g786(.A(G953), .B1(new_n313), .B2(new_n322), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n860), .A2(new_n873), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n920), .B1(G898), .B2(new_n275), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  AOI21_X1  g791(.A(new_n275), .B1(G227), .B2(G900), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n978), .B(KEYINPUT124), .Z(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n746), .A2(new_n841), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n698), .A2(new_n700), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n698), .A2(new_n984), .A3(new_n700), .A4(new_n981), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n794), .A2(new_n789), .ZN(new_n986));
  NOR4_X1   g800(.A1(new_n677), .A2(new_n763), .A3(new_n754), .A4(new_n870), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n275), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n533), .B1(KEYINPUT30), .B2(new_n499), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT122), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n435), .A2(new_n436), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n715), .A2(new_n734), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n981), .B(new_n768), .C1(new_n778), .C2(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(new_n765), .ZN(new_n1000));
  INV_X1    g814(.A(new_n986), .ZN(new_n1001));
  AOI21_X1  g815(.A(G953), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n997), .B1(new_n1002), .B2(new_n666), .ZN(new_n1003));
  INV_X1    g817(.A(new_n666), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n986), .A2(new_n999), .A3(new_n765), .ZN(new_n1005));
  OAI211_X1 g819(.A(KEYINPUT125), .B(new_n1004), .C1(new_n1005), .C2(G953), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n995), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n996), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g823(.A(KEYINPUT126), .B(new_n995), .C1(new_n1003), .C2(new_n1006), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n980), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1007), .A2(new_n980), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n990), .A2(KEYINPUT123), .A3(new_n995), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT123), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n996), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1011), .A2(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  INV_X1    g833(.A(new_n974), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1019), .B1(new_n989), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n690), .ZN(new_n1022));
  INV_X1    g836(.A(new_n536), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1019), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n690), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n902), .A2(new_n903), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1005), .A2(new_n974), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(new_n1019), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n914), .B1(new_n1028), .B2(new_n1023), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1022), .A2(new_n1026), .A3(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(KEYINPUT127), .ZN(G57));
endmodule


