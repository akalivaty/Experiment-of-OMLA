//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  OR2_X1    g003(.A1(G57gat), .A2(G64gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G57gat), .A2(G64gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT93), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(new_n202), .ZN(new_n210));
  AND2_X1   g009(.A1(G71gat), .A2(G78gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT93), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n211), .A2(new_n212), .ZN(new_n215));
  AND2_X1   g014(.A1(G57gat), .A2(G64gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G57gat), .A2(G64gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n215), .A2(new_n218), .A3(new_n209), .A4(new_n204), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(KEYINPUT21), .ZN(new_n221));
  NAND2_X1  g020(.A1(G231gat), .A2(G233gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n223), .A2(G127gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(G127gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G22gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G15gat), .ZN(new_n228));
  INV_X1    g027(.A(G15gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G22gat), .ZN(new_n230));
  INV_X1    g029(.A(G1gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT16), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(G1gat), .B1(new_n228), .B2(new_n230), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT89), .B(G8gat), .ZN(new_n236));
  NOR3_X1   g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G15gat), .B(G22gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT87), .B1(new_n239), .B2(G1gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n228), .A2(new_n230), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT87), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n231), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n243), .A3(new_n233), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n244), .A2(KEYINPUT88), .A3(G8gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT88), .B1(new_n244), .B2(G8gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n238), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(KEYINPUT21), .B2(new_n220), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n226), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n250));
  INV_X1    g049(.A(G155gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G183gat), .B(G211gat), .Z(new_n253));
  XNOR2_X1  g052(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n249), .B(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G43gat), .A2(G50gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G43gat), .A2(G50gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT15), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT84), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n261), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT14), .ZN(new_n264));
  INV_X1    g063(.A(G29gat), .ZN(new_n265));
  INV_X1    g064(.A(G36gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR3_X1   g068(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT85), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n263), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G29gat), .A2(G36gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n258), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n270), .B1(new_n260), .B2(new_n262), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT15), .ZN(new_n276));
  INV_X1    g075(.A(G43gat), .ZN(new_n277));
  INV_X1    g076(.A(G50gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT86), .B(G43gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n258), .A2(new_n273), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n275), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n274), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G99gat), .A2(G106gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT8), .ZN(new_n287));
  NAND2_X1  g086(.A1(G85gat), .A2(G92gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT7), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G85gat), .ZN(new_n291));
  INV_X1    g090(.A(G92gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n287), .A2(new_n290), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G99gat), .B(G106gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI22_X1  g100(.A1(KEYINPUT8), .A2(new_n286), .B1(new_n291), .B2(new_n292), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n296), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G232gat), .A2(G233gat), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n285), .A2(new_n304), .B1(KEYINPUT41), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT17), .B1(new_n274), .B2(new_n283), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT17), .ZN(new_n308));
  INV_X1    g107(.A(new_n279), .ZN(new_n309));
  XOR2_X1   g108(.A(KEYINPUT86), .B(G43gat), .Z(new_n310));
  OAI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(G50gat), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n258), .A2(new_n273), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n263), .A2(new_n267), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n273), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n267), .A2(new_n268), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT85), .B1(new_n317), .B2(new_n266), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n315), .B1(new_n319), .B2(new_n263), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n308), .B(new_n314), .C1(new_n320), .C2(new_n258), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n307), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n304), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n322), .A2(KEYINPUT94), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT94), .B1(new_n322), .B2(new_n323), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n306), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G190gat), .B(G218gat), .Z(new_n327));
  OR2_X1    g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n305), .A2(KEYINPUT41), .ZN(new_n329));
  XNOR2_X1  g128(.A(G134gat), .B(G162gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n326), .A2(new_n327), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n328), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n255), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n303), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n301), .A2(new_n296), .A3(new_n302), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n220), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n219), .B(new_n214), .C1(new_n298), .C2(new_n303), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(G230gat), .A3(G233gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G120gat), .B(G148gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G176gat), .B(G204gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT10), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT95), .ZN(new_n351));
  NAND2_X1  g150(.A1(G230gat), .A2(G233gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT95), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n353), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n351), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT96), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n351), .A2(new_n357), .A3(new_n352), .A4(new_n354), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n346), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n352), .B(KEYINPUT97), .Z(new_n360));
  AND3_X1   g159(.A1(new_n350), .A2(KEYINPUT98), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT98), .B1(new_n350), .B2(new_n360), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n345), .B1(new_n363), .B2(new_n342), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n336), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT92), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(G228gat), .A2(G233gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G141gat), .B(G148gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n373), .ZN(new_n376));
  INV_X1    g175(.A(G162gat), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT2), .B1(new_n251), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G197gat), .B(G204gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT22), .ZN(new_n386));
  INV_X1    g185(.A(G211gat), .ZN(new_n387));
  INV_X1    g186(.A(G218gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G211gat), .B(G218gat), .Z(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT70), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n390), .B(new_n391), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(KEYINPUT70), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n384), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT3), .B1(new_n396), .B2(new_n383), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n370), .B(new_n395), .C1(new_n397), .C2(new_n380), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n375), .A2(new_n379), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n393), .A2(new_n383), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n370), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT80), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(KEYINPUT80), .B(new_n370), .C1(new_n395), .C2(new_n401), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n398), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G22gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(new_n278), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n227), .B(new_n398), .C1(new_n404), .C2(new_n405), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n407), .B2(new_n411), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n369), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n407), .A2(new_n411), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n409), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n368), .A3(new_n412), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G169gat), .ZN(new_n420));
  INV_X1    g219(.A(G176gat), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT23), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n422), .B1(G169gat), .B2(G176gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT23), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(KEYINPUT25), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(G183gat), .A2(G190gat), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n426), .A2(KEYINPUT24), .ZN(new_n427));
  XNOR2_X1  g226(.A(G183gat), .B(G190gat), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT24), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT25), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT64), .B(G169gat), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT23), .A3(new_n421), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n423), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n435), .B2(new_n430), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n426), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT27), .B(G183gat), .ZN(new_n439));
  INV_X1    g238(.A(G190gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(KEYINPUT65), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(G169gat), .A2(G176gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT26), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n447), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  XOR2_X1   g248(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n450));
  OAI211_X1 g249(.A(new_n444), .B(new_n449), .C1(new_n441), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n437), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT71), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n437), .A2(KEYINPUT71), .A3(new_n451), .ZN(new_n455));
  AND2_X1   g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(KEYINPUT29), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n437), .A2(new_n456), .A3(new_n451), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n394), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n454), .A2(new_n455), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n461), .A2(new_n456), .B1(new_n452), .B2(new_n457), .ZN(new_n462));
  OAI211_X1 g261(.A(KEYINPUT72), .B(new_n460), .C1(new_n462), .C2(new_n394), .ZN(new_n463));
  OR2_X1    g262(.A1(new_n460), .A2(KEYINPUT72), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G8gat), .B(G36gat), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT73), .ZN(new_n467));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT30), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n472));
  XNOR2_X1  g271(.A(G1gat), .B(G29gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(KEYINPUT0), .ZN(new_n474));
  XNOR2_X1  g273(.A(G57gat), .B(G85gat), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n474), .B(new_n475), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G127gat), .B(G134gat), .Z(new_n478));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT66), .ZN(new_n481));
  XNOR2_X1  g280(.A(G113gat), .B(G120gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(KEYINPUT1), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(KEYINPUT66), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT1), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n479), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n478), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n399), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n484), .A2(new_n489), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n380), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G225gat), .A2(G233gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(KEYINPUT5), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n399), .A2(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n490), .A2(new_n498), .A3(new_n382), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT76), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT76), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n490), .A2(new_n501), .A3(new_n498), .A4(new_n382), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n493), .B(KEYINPUT4), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n495), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT5), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(KEYINPUT77), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n505), .A2(new_n507), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n477), .B(new_n497), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n472), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n497), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n505), .A2(new_n507), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n505), .A2(new_n507), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n516), .A2(KEYINPUT78), .A3(KEYINPUT6), .A4(new_n477), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n497), .B1(new_n508), .B2(new_n509), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n476), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(new_n511), .A3(new_n510), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n471), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n465), .A2(KEYINPUT30), .A3(new_n470), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n463), .A2(new_n464), .A3(new_n469), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n419), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G227gat), .ZN(new_n530));
  INV_X1    g329(.A(G233gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n452), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n437), .A2(KEYINPUT68), .A3(new_n451), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n490), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n452), .A2(new_n533), .A3(new_n492), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT34), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n532), .A3(new_n537), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT32), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT33), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G15gat), .B(G43gat), .Z(new_n544));
  XNOR2_X1  g343(.A(G71gat), .B(G99gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n541), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n546), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n540), .B(KEYINPUT32), .C1(new_n542), .C2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n539), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n539), .B1(new_n547), .B2(new_n549), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n551), .A2(new_n552), .A3(KEYINPUT36), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n539), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n547), .A2(new_n549), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n550), .B1(new_n557), .B2(KEYINPUT69), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT69), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n552), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n554), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n529), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n503), .A2(new_n504), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n496), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT39), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n494), .A2(new_n496), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT81), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n566), .B(new_n570), .C1(new_n569), .C2(new_n568), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n571), .B(new_n476), .C1(KEYINPUT39), .C2(new_n566), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT40), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n572), .A2(new_n573), .B1(new_n477), .B2(new_n516), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n523), .A2(new_n525), .ZN(new_n575));
  OAI221_X1 g374(.A(new_n574), .B1(new_n573), .B2(new_n572), .C1(new_n471), .C2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n470), .B1(new_n465), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n458), .A2(new_n396), .A3(new_n459), .ZN(new_n579));
  OAI211_X1 g378(.A(KEYINPUT37), .B(new_n579), .C1(new_n462), .C2(new_n396), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT38), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582));
  INV_X1    g381(.A(new_n465), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n582), .B1(new_n583), .B2(KEYINPUT37), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n581), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n518), .B(new_n521), .C1(new_n469), .C2(new_n583), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n576), .B(new_n419), .C1(new_n585), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n522), .A2(new_n528), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n561), .A2(new_n419), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT35), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n575), .A2(new_n471), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT82), .B(KEYINPUT35), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n419), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n518), .A2(new_n521), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n551), .A2(new_n552), .ZN(new_n595));
  AND2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n564), .A2(new_n587), .B1(new_n590), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n233), .B1(new_n235), .B2(new_n242), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n239), .A2(KEYINPUT87), .A3(G1gat), .ZN(new_n600));
  OAI21_X1  g399(.A(G8gat), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT88), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n244), .A2(KEYINPUT88), .A3(G8gat), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n237), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n322), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n247), .A2(new_n285), .ZN(new_n607));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT18), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT18), .A4(new_n608), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n284), .B(new_n238), .C1(new_n245), .C2(new_n246), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n608), .B(KEYINPUT13), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT90), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT90), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G113gat), .B(G141gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G169gat), .B(G197gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n630));
  INV_X1    g429(.A(new_n616), .ZN(new_n631));
  AOI211_X1 g430(.A(KEYINPUT90), .B(new_n631), .C1(new_n607), .C2(new_n614), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n611), .A2(new_n612), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n629), .A2(new_n635), .A3(KEYINPUT91), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT91), .B1(new_n629), .B2(new_n635), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n367), .B1(new_n598), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n590), .A2(new_n597), .ZN(new_n640));
  INV_X1    g439(.A(new_n419), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n588), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n558), .ZN(new_n643));
  INV_X1    g442(.A(new_n560), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n553), .B1(new_n645), .B2(KEYINPUT36), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n587), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n638), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(KEYINPUT92), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n366), .B1(new_n639), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n594), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  INV_X1    g453(.A(new_n591), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  AND3_X1   g455(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(G8gat), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n651), .B2(new_n655), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT42), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(KEYINPUT42), .B2(new_n657), .ZN(G1325gat));
  INV_X1    g460(.A(new_n651), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n662), .B2(new_n646), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n651), .A2(new_n229), .A3(new_n595), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(G1326gat));
  NAND2_X1  g464(.A1(new_n651), .A2(new_n641), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  INV_X1    g467(.A(new_n255), .ZN(new_n669));
  INV_X1    g468(.A(new_n365), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n335), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n672), .B1(new_n639), .B2(new_n650), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n265), .A3(new_n652), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  INV_X1    g477(.A(new_n335), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n598), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n648), .A2(KEYINPUT44), .A3(new_n335), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n629), .A2(new_n635), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n671), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT99), .Z(new_n686));
  AND3_X1   g485(.A1(new_n683), .A2(new_n652), .A3(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n676), .B(new_n677), .C1(new_n265), .C2(new_n687), .ZN(G1328gat));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n266), .A3(new_n655), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT46), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(KEYINPUT46), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n683), .A2(new_n655), .A3(new_n686), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n690), .B(new_n691), .C1(new_n266), .C2(new_n692), .ZN(G1329gat));
  INV_X1    g492(.A(new_n672), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n551), .A2(new_n552), .A3(new_n310), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT92), .B1(new_n648), .B2(new_n649), .ZN(new_n696));
  AOI211_X1 g495(.A(new_n367), .B(new_n638), .C1(new_n640), .C2(new_n647), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n694), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n673), .A2(KEYINPUT100), .A3(new_n695), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT47), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n680), .A2(new_n681), .A3(new_n563), .A4(new_n686), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT101), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n707), .A3(new_n280), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n700), .A2(new_n701), .B1(new_n310), .B2(new_n704), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n703), .A2(new_n708), .B1(new_n709), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g509(.A1(new_n673), .A2(new_n641), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n278), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n683), .A2(G50gat), .A3(new_n641), .A4(new_n686), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT102), .B(KEYINPUT48), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n684), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n336), .A2(new_n718), .A3(new_n670), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n598), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n652), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g521(.A1(new_n598), .A2(new_n591), .A3(new_n719), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(G1333gat));
  AND3_X1   g526(.A1(new_n720), .A2(G71gat), .A3(new_n563), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n720), .A2(new_n595), .ZN(new_n729));
  AOI21_X1  g528(.A(G71gat), .B1(new_n729), .B2(KEYINPUT103), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT103), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n720), .A2(new_n731), .A3(new_n595), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT104), .B(KEYINPUT50), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n733), .B(new_n735), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n641), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g537(.A(new_n679), .B1(new_n640), .B2(new_n647), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n669), .A2(new_n684), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n739), .A2(KEYINPUT51), .A3(new_n740), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n740), .ZN(new_n747));
  NOR4_X1   g546(.A1(new_n598), .A2(new_n742), .A3(new_n679), .A4(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n652), .A2(new_n291), .A3(new_n670), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT106), .ZN(new_n752));
  NOR4_X1   g551(.A1(new_n682), .A2(new_n594), .A3(new_n365), .A4(new_n747), .ZN(new_n753));
  OAI22_X1  g552(.A1(new_n750), .A2(new_n752), .B1(new_n753), .B2(new_n291), .ZN(G1336gat));
  NOR3_X1   g553(.A1(new_n591), .A2(G92gat), .A3(new_n365), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(new_n746), .B2(new_n749), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n747), .A2(new_n365), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n680), .A2(new_n681), .A3(new_n655), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G92gat), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n739), .B2(new_n740), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n755), .B1(new_n748), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT107), .B1(new_n764), .B2(KEYINPUT52), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n766), .B(new_n757), .C1(new_n760), .C2(new_n763), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n761), .B1(new_n765), .B2(new_n767), .ZN(G1337gat));
  INV_X1    g567(.A(G99gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n595), .A2(new_n769), .A3(new_n670), .ZN(new_n770));
  NOR4_X1   g569(.A1(new_n682), .A2(new_n646), .A3(new_n365), .A4(new_n747), .ZN(new_n771));
  OAI22_X1  g570(.A1(new_n750), .A2(new_n770), .B1(new_n771), .B2(new_n769), .ZN(G1338gat));
  NAND4_X1  g571(.A1(new_n680), .A2(new_n681), .A3(new_n641), .A4(new_n758), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT108), .B(G106gat), .Z(new_n774));
  AOI21_X1  g573(.A(KEYINPUT53), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OR3_X1    g574(.A1(new_n419), .A2(G106gat), .A3(new_n365), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n750), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n773), .A2(new_n778), .A3(new_n774), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n773), .B2(new_n774), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n776), .B1(new_n743), .B2(new_n745), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(G1339gat));
  NOR2_X1   g583(.A1(new_n655), .A2(new_n594), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OR2_X1    g585(.A1(new_n350), .A2(new_n360), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT54), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n788), .B1(new_n356), .B2(new_n358), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n350), .A2(new_n360), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT98), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n350), .A2(KEYINPUT98), .A3(new_n360), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT54), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n790), .B1(new_n795), .B2(new_n345), .ZN(new_n796));
  INV_X1    g595(.A(new_n345), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT110), .B(new_n797), .C1(new_n363), .C2(KEYINPUT54), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n789), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n359), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n798), .ZN(new_n801));
  INV_X1    g600(.A(new_n789), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(new_n805), .A3(new_n684), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n615), .A2(new_n616), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n608), .B1(new_n606), .B2(new_n607), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n626), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n670), .A2(new_n629), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n335), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n629), .A2(new_n809), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n335), .A2(new_n800), .A3(new_n805), .A4(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n255), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n336), .A2(new_n718), .A3(new_n365), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n786), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n589), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n684), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n641), .B1(new_n816), .B2(new_n817), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(new_n595), .A3(new_n785), .ZN(new_n824));
  INV_X1    g623(.A(G113gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n824), .A2(new_n825), .A3(new_n638), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n822), .A2(new_n826), .ZN(G1340gat));
  AOI21_X1  g626(.A(G120gat), .B1(new_n821), .B2(new_n670), .ZN(new_n828));
  INV_X1    g627(.A(G120gat), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n824), .A2(new_n829), .A3(new_n365), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n828), .A2(new_n830), .ZN(G1341gat));
  OAI21_X1  g630(.A(G127gat), .B1(new_n824), .B2(new_n255), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n255), .A2(G127gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n820), .B2(new_n833), .ZN(G1342gat));
  OR3_X1    g633(.A1(new_n820), .A2(G134gat), .A3(new_n679), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(KEYINPUT56), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT111), .Z(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n824), .B2(new_n679), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n837), .B(new_n838), .C1(KEYINPUT56), .C2(new_n835), .ZN(G1343gat));
  NOR2_X1   g638(.A1(new_n786), .A2(new_n563), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n419), .B1(new_n816), .B2(new_n817), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT112), .B1(new_n841), .B2(KEYINPUT57), .ZN(new_n842));
  XNOR2_X1  g641(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n803), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n800), .B(new_n844), .C1(new_n636), .C2(new_n637), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n335), .B1(new_n845), .B2(new_n811), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n255), .B1(new_n846), .B2(new_n815), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n817), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n419), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n842), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n841), .A2(KEYINPUT112), .A3(KEYINPUT57), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n840), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G141gat), .B1(new_n854), .B2(new_n638), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT58), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n816), .A2(new_n817), .ZN(new_n857));
  AND4_X1   g656(.A1(new_n641), .A2(new_n857), .A3(new_n646), .A4(new_n785), .ZN(new_n858));
  INV_X1    g657(.A(G141gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n649), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n855), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n684), .B(new_n840), .C1(new_n852), .C2(new_n853), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(G141gat), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n862), .B2(G141gat), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n860), .B(KEYINPUT115), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n861), .B1(new_n867), .B2(new_n856), .ZN(G1344gat));
  INV_X1    g667(.A(G148gat), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(KEYINPUT59), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n854), .B2(new_n365), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n857), .A2(new_n850), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n366), .A2(new_n649), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n419), .B1(new_n847), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(KEYINPUT57), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n876), .A2(new_n670), .A3(new_n840), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT59), .B1(new_n877), .B2(new_n869), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n871), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n858), .A2(new_n869), .A3(new_n670), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1345gat));
  OAI21_X1  g680(.A(G155gat), .B1(new_n854), .B2(new_n255), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n858), .A2(new_n251), .A3(new_n669), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1346gat));
  NOR3_X1   g683(.A1(new_n854), .A2(new_n377), .A3(new_n679), .ZN(new_n885));
  AOI21_X1  g684(.A(G162gat), .B1(new_n858), .B2(new_n335), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1347gat));
  NAND2_X1  g686(.A1(new_n596), .A2(new_n655), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT116), .Z(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n823), .ZN(new_n890));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n638), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT117), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n655), .A2(new_n594), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n589), .B(new_n893), .C1(new_n816), .C2(new_n817), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(new_n433), .A3(new_n684), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1348gat));
  OAI21_X1  g695(.A(G176gat), .B1(new_n890), .B2(new_n365), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n421), .A3(new_n670), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1349gat));
  OAI21_X1  g698(.A(G183gat), .B1(new_n890), .B2(new_n255), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n894), .A2(new_n439), .A3(new_n669), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(KEYINPUT118), .A3(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n894), .A2(new_n440), .A3(new_n335), .ZN(new_n904));
  OAI21_X1  g703(.A(G190gat), .B1(new_n890), .B2(new_n679), .ZN(new_n905));
  XOR2_X1   g704(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n906));
  AND2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT120), .B(new_n904), .C1(new_n907), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1351gat));
  INV_X1    g712(.A(new_n841), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n563), .A2(new_n893), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n914), .A2(new_n916), .A3(G197gat), .A4(new_n718), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT121), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n876), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n915), .A2(new_n649), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G197gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT123), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT123), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n926), .B(new_n918), .C1(new_n922), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1352gat));
  NOR2_X1   g727(.A1(new_n914), .A2(new_n916), .ZN(new_n929));
  INV_X1    g728(.A(G204gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n930), .A3(new_n670), .ZN(new_n931));
  AND2_X1   g730(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n932));
  NOR2_X1   g731(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n920), .A2(new_n365), .A3(new_n916), .ZN(new_n935));
  OAI221_X1 g734(.A(new_n934), .B1(new_n932), .B2(new_n931), .C1(new_n935), .C2(new_n930), .ZN(G1353gat));
  NAND2_X1  g735(.A1(new_n915), .A2(new_n669), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n387), .A3(new_n841), .ZN(new_n939));
  INV_X1    g738(.A(new_n843), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n801), .B2(new_n802), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT91), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n628), .B1(new_n613), .B2(new_n621), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n633), .A2(new_n634), .A3(new_n627), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n629), .A2(new_n635), .A3(KEYINPUT91), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n810), .B1(new_n947), .B2(new_n800), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n814), .B1(new_n948), .B2(new_n335), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n873), .B1(new_n949), .B2(new_n255), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n849), .B1(new_n950), .B2(new_n419), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n937), .B1(new_n951), .B2(new_n872), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n387), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n876), .B2(new_n938), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n847), .A2(new_n874), .ZN(new_n958));
  AOI21_X1  g757(.A(KEYINPUT57), .B1(new_n958), .B2(new_n641), .ZN(new_n959));
  AOI211_X1 g758(.A(new_n849), .B(new_n419), .C1(new_n816), .C2(new_n817), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n953), .B(new_n938), .C1(new_n959), .C2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(G211gat), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT63), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n962), .A2(new_n963), .A3(new_n955), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n939), .B1(new_n957), .B2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI211_X1 g766(.A(KEYINPUT126), .B(new_n939), .C1(new_n957), .C2(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(G1354gat));
  AOI21_X1  g768(.A(G218gat), .B1(new_n929), .B2(new_n335), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n920), .A2(new_n916), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n335), .A2(G218gat), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT127), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n970), .B1(new_n971), .B2(new_n973), .ZN(G1355gat));
endmodule


