//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  XNOR2_X1  g000(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT33), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT28), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT66), .B(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT68), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT27), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(G183gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G183gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT27), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(G183gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n205), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n212), .A2(new_n213), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT69), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT66), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G190gat), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n219), .A2(new_n221), .A3(KEYINPUT28), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n212), .A2(new_n213), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n217), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n215), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT70), .B1(new_n227), .B2(new_n228), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n227), .A2(KEYINPUT70), .A3(new_n228), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n232), .A2(new_n233), .B1(G183gat), .B2(G190gat), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n226), .A2(KEYINPUT71), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT71), .B1(new_n226), .B2(new_n234), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT1), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT72), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT72), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n242));
  XOR2_X1   g041(.A(G127gat), .B(G134gat), .Z(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  OR3_X1    g043(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G176gat), .ZN(new_n248));
  INV_X1    g047(.A(G169gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT23), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n229), .A2(KEYINPUT23), .ZN(new_n251));
  OAI22_X1  g050(.A1(new_n248), .A2(new_n250), .B1(new_n251), .B2(new_n227), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255));
  NAND2_X1  g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n247), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(KEYINPUT65), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(G183gat), .A3(G190gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(new_n255), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n219), .A2(new_n221), .A3(new_n211), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n262), .A2(new_n263), .A3(new_n253), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n227), .B1(KEYINPUT23), .B2(new_n229), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n266), .A3(KEYINPUT23), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT25), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n264), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n264), .B2(new_n269), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n258), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n237), .A2(KEYINPUT73), .A3(new_n246), .A4(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n212), .A2(new_n213), .A3(new_n223), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n223), .B1(new_n212), .B2(new_n213), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT27), .B(G183gat), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n206), .B(new_n209), .C1(new_n279), .C2(new_n207), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n278), .A2(new_n222), .B1(new_n280), .B2(new_n205), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n232), .A2(new_n233), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n256), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n275), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n226), .A2(KEYINPUT71), .A3(new_n234), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(new_n273), .A3(new_n246), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(new_n273), .A3(new_n285), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n244), .A2(new_n245), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G227gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n292), .A2(KEYINPUT74), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT74), .B1(new_n292), .B2(new_n294), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n204), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G15gat), .B(G43gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G71gat), .B(G99gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n274), .A2(new_n288), .A3(new_n293), .A4(new_n291), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT75), .ZN(new_n304));
  OR3_X1    g103(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT34), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(KEYINPUT34), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n303), .B2(KEYINPUT34), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n203), .B1(new_n301), .B2(KEYINPUT33), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n295), .B2(new_n296), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n302), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n302), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n202), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n292), .A2(new_n294), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n292), .A2(KEYINPUT74), .A3(new_n294), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n318), .A2(new_n319), .B1(new_n203), .B2(KEYINPUT33), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n310), .B1(new_n320), .B2(new_n300), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n319), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n297), .A2(new_n301), .B1(new_n324), .B2(new_n309), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n308), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT78), .A3(new_n202), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n322), .B1(new_n325), .B2(KEYINPUT76), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n321), .A2(new_n330), .A3(new_n308), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT36), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335));
  AND2_X1   g134(.A1(G211gat), .A2(G218gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(G211gat), .A2(G218gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n336), .A2(KEYINPUT22), .ZN(new_n339));
  INV_X1    g138(.A(G197gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT79), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G197gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G204gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n341), .A2(new_n343), .A3(G204gat), .ZN(new_n347));
  AOI211_X1 g146(.A(new_n338), .B(new_n339), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n348), .B2(KEYINPUT89), .ZN(new_n349));
  INV_X1    g148(.A(new_n339), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n341), .A2(new_n343), .A3(G204gat), .ZN(new_n351));
  AOI21_X1  g150(.A(G204gat), .B1(new_n341), .B2(new_n343), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n338), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n346), .A2(new_n347), .ZN(new_n355));
  INV_X1    g154(.A(new_n338), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(new_n350), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n349), .B1(new_n358), .B2(KEYINPUT89), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n360));
  XNOR2_X1  g159(.A(G155gat), .B(G162gat), .ZN(new_n361));
  INV_X1    g160(.A(G141gat), .ZN(new_n362));
  INV_X1    g161(.A(G148gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365));
  AND2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT2), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G162gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT81), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n367), .B1(new_n374), .B2(G155gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(KEYINPUT81), .B(G162gat), .ZN(new_n379));
  INV_X1    g178(.A(G155gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT2), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n370), .A2(G155gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(G162gat), .ZN(new_n383));
  AND4_X1   g182(.A1(new_n382), .A2(new_n364), .A3(new_n383), .A4(new_n365), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT82), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n369), .B1(new_n378), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n377), .B1(new_n375), .B2(new_n376), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(new_n384), .A3(KEYINPUT82), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT84), .A3(new_n369), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n359), .A2(new_n360), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n368), .B1(new_n389), .B2(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n360), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n358), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n335), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n358), .B2(new_n396), .ZN(new_n399));
  OAI211_X1 g198(.A(G228gat), .B(G233gat), .C1(new_n399), .C2(new_n394), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n400), .A2(KEYINPUT90), .A3(new_n397), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT90), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n356), .B1(new_n355), .B2(new_n350), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n396), .B1(new_n403), .B2(new_n348), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n360), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n335), .B1(new_n405), .B2(new_n386), .ZN(new_n406));
  INV_X1    g205(.A(new_n358), .ZN(new_n407));
  AOI211_X1 g206(.A(KEYINPUT3), .B(new_n368), .C1(new_n389), .C2(new_n390), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(KEYINPUT29), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n402), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n398), .B1(new_n401), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G22gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n412), .A2(KEYINPUT91), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI221_X1 g213(.A(new_n398), .B1(KEYINPUT91), .B2(new_n412), .C1(new_n401), .C2(new_n410), .ZN(new_n415));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(G50gat), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT87), .B(KEYINPUT31), .Z(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n411), .A2(new_n412), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n398), .B(G22gat), .C1(new_n401), .C2(new_n410), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n419), .B(KEYINPUT88), .Z(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n388), .A2(new_n426), .A3(new_n246), .A4(new_n392), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n394), .A2(new_n246), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n427), .A2(KEYINPUT86), .B1(KEYINPUT4), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT84), .B1(new_n391), .B2(new_n369), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n387), .B(new_n368), .C1(new_n389), .C2(new_n390), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n430), .A2(new_n431), .A3(new_n290), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT86), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n426), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n290), .B1(new_n394), .B2(new_n360), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(new_n408), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT83), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT94), .B(KEYINPUT39), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT39), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n386), .B(new_n246), .ZN(new_n446));
  INV_X1    g245(.A(new_n441), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n437), .B1(new_n429), .B2(new_n434), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n447), .ZN(new_n450));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(KEYINPUT0), .ZN(new_n452));
  XNOR2_X1  g251(.A(G57gat), .B(G85gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  NAND4_X1  g253(.A1(new_n444), .A2(new_n450), .A3(KEYINPUT40), .A4(new_n454), .ZN(new_n455));
  AND2_X1   g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456));
  AND4_X1   g255(.A1(new_n273), .A2(new_n284), .A3(new_n285), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(KEYINPUT29), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n226), .A2(new_n234), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n273), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n358), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n289), .A2(new_n458), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n273), .A2(new_n460), .A3(new_n456), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n407), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G8gat), .B(G36gat), .ZN(new_n466));
  XNOR2_X1  g265(.A(G64gat), .B(G92gat), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n466), .B(new_n467), .Z(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n462), .A2(new_n465), .A3(KEYINPUT30), .A4(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n462), .A2(new_n465), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n468), .B(KEYINPUT80), .Z(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n471), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT93), .ZN(new_n477));
  INV_X1    g276(.A(new_n454), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT5), .B1(new_n446), .B2(new_n447), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n432), .B2(new_n426), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n388), .A2(new_n246), .A3(new_n392), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(KEYINPUT85), .A3(KEYINPUT4), .ZN(new_n483));
  INV_X1    g282(.A(new_n428), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n426), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n437), .A2(new_n441), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n479), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT5), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n438), .A2(new_n489), .A3(new_n447), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n490), .B1(new_n434), .B2(new_n429), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n478), .B1(new_n488), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n471), .A2(new_n475), .A3(new_n493), .A4(new_n472), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n455), .A2(new_n477), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n450), .A2(new_n454), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT40), .B1(new_n496), .B2(new_n444), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n425), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT6), .B(new_n478), .C1(new_n488), .C2(new_n491), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT95), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n435), .A2(new_n489), .A3(new_n487), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n438), .A2(new_n447), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n482), .A2(KEYINPUT4), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n504), .A2(new_n480), .B1(new_n426), .B2(new_n484), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n503), .B1(new_n505), .B2(new_n483), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n502), .B1(new_n506), .B2(new_n479), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT95), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT6), .A4(new_n478), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n407), .B1(new_n457), .B2(new_n461), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n463), .A2(new_n358), .A3(new_n464), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT37), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT38), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n474), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n513), .B(new_n515), .C1(new_n473), .C2(KEYINPUT37), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n469), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n473), .A2(KEYINPUT37), .ZN(new_n518));
  INV_X1    g317(.A(new_n468), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n473), .A2(KEYINPUT37), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n517), .B1(KEYINPUT38), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n454), .B(new_n502), .C1(new_n506), .C2(new_n479), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n492), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n500), .ZN(new_n527));
  INV_X1    g326(.A(new_n476), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT92), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n420), .A2(new_n424), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n530), .B1(new_n420), .B2(new_n424), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n499), .A2(new_n526), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n476), .B1(new_n525), .B2(new_n500), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n325), .A2(KEYINPUT76), .A3(new_n322), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n308), .B1(new_n321), .B2(new_n330), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n535), .B(new_n425), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n539));
  INV_X1    g338(.A(new_n327), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n425), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n477), .A2(new_n494), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n510), .A2(new_n525), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n334), .A2(new_n534), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT97), .ZN(new_n549));
  XOR2_X1   g348(.A(G169gat), .B(G197gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(KEYINPUT96), .B(KEYINPUT11), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(KEYINPUT12), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G43gat), .B(G50gat), .Z(new_n556));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT98), .B(G36gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(G29gat), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT14), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(G29gat), .B2(G36gat), .ZN(new_n562));
  OR3_X1    g361(.A1(new_n561), .A2(G29gat), .A3(G36gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n558), .B1(new_n564), .B2(KEYINPUT99), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n557), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n566), .A2(new_n560), .A3(new_n562), .A4(new_n563), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n567), .B(new_n558), .C1(KEYINPUT99), .C2(new_n564), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT100), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT16), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(G1gat), .ZN(new_n575));
  INV_X1    g374(.A(G8gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n571), .B(KEYINPUT100), .ZN(new_n577));
  INV_X1    g376(.A(G1gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n576), .B1(new_n575), .B2(new_n579), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n569), .B(new_n570), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n570), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n575), .A2(new_n579), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(G8gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n575), .A2(new_n576), .A3(new_n579), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n584), .B1(new_n569), .B2(new_n570), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n582), .B(new_n583), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT18), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n569), .A2(new_n570), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n587), .A2(new_n595), .A3(new_n588), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n582), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n583), .B(KEYINPUT13), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n599), .B1(new_n591), .B2(new_n592), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n555), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n593), .A2(KEYINPUT101), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT101), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n591), .A2(new_n603), .A3(new_n592), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n554), .B(new_n599), .C1(new_n592), .C2(new_n591), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n547), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G57gat), .B(G64gat), .Z(new_n610));
  NAND2_X1  g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT9), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G71gat), .B(G78gat), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n610), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n615), .B2(new_n614), .ZN(new_n617));
  INV_X1    g416(.A(new_n614), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n618), .A2(new_n610), .A3(KEYINPUT102), .A4(new_n613), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n620), .A2(KEYINPUT21), .ZN(new_n621));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G127gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  AOI211_X1 g424(.A(new_n581), .B(new_n580), .C1(KEYINPUT21), .C2(new_n620), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G155gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n627), .B(new_n631), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n590), .ZN(new_n634));
  NAND2_X1  g433(.A1(G85gat), .A2(G92gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT7), .ZN(new_n636));
  XNOR2_X1  g435(.A(G99gat), .B(G106gat), .ZN(new_n637));
  NAND2_X1  g436(.A1(G99gat), .A2(G106gat), .ZN(new_n638));
  INV_X1    g437(.A(G85gat), .ZN(new_n639));
  INV_X1    g438(.A(G92gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(KEYINPUT8), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n636), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n637), .B1(new_n636), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n634), .A2(new_n585), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n595), .ZN(new_n649));
  AND2_X1   g448(.A1(G232gat), .A2(G233gat), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n649), .A2(new_n644), .B1(KEYINPUT41), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G134gat), .B(G162gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G190gat), .B(G218gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT105), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n650), .A2(KEYINPUT41), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT103), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n656), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n653), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n648), .A2(new_n651), .A3(new_n660), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n654), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n654), .B2(new_n661), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n633), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n620), .A2(new_n644), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n617), .B(new_n619), .C1(new_n642), .C2(new_n643), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n645), .A2(KEYINPUT106), .A3(new_n619), .A4(new_n617), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT10), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n620), .A2(KEYINPUT10), .A3(new_n644), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n667), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n671), .A2(G230gat), .A3(G233gat), .A4(new_n672), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(G120gat), .B(G148gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n678), .B(new_n679), .Z(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(new_n676), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n609), .A2(new_n666), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n527), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n578), .ZN(G1324gat));
  INV_X1    g487(.A(new_n543), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT108), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n686), .B2(new_n689), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(G8gat), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT16), .B(G8gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT109), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n690), .A2(KEYINPUT42), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n691), .B2(new_n693), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n694), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(G1325gat));
  INV_X1    g500(.A(G15gat), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n702), .A3(new_n334), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n686), .B2(new_n327), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n703), .B1(new_n706), .B2(new_n707), .ZN(G1326gat));
  INV_X1    g507(.A(new_n533), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n686), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT43), .B(G22gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1327gat));
  NAND2_X1  g511(.A1(new_n632), .A2(new_n685), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n664), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT111), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n609), .A2(new_n715), .ZN(new_n716));
  OR3_X1    g515(.A1(new_n716), .A2(G29gat), .A3(new_n527), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n547), .B2(new_n664), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n662), .A2(new_n663), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n529), .A2(new_n533), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n510), .A2(new_n525), .A3(new_n522), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(new_n498), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n313), .A2(new_n314), .B1(new_n332), .B2(KEYINPUT36), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n328), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n327), .A2(new_n543), .A3(new_n542), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n545), .A2(new_n727), .B1(new_n538), .B2(KEYINPUT35), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT44), .B(new_n721), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n720), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n713), .A2(new_n608), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G29gat), .B1(new_n732), .B2(new_n527), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n733), .ZN(G1328gat));
  OAI21_X1  g533(.A(new_n559), .B1(new_n732), .B2(new_n689), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n716), .A2(new_n689), .A3(new_n559), .ZN(new_n736));
  NAND2_X1  g535(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT112), .B(KEYINPUT46), .Z(new_n739));
  OAI211_X1 g538(.A(new_n735), .B(new_n738), .C1(new_n736), .C2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(new_n334), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n720), .A2(new_n729), .A3(new_n741), .A4(new_n731), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G43gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n327), .A2(G43gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n609), .A2(new_n715), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n747), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n748), .A2(new_n743), .A3(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n751));
  OAI21_X1  g550(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(G1330gat));
  INV_X1    g551(.A(new_n425), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n730), .A2(new_n753), .A3(new_n731), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G50gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n716), .A2(G50gat), .A3(new_n709), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(new_n757), .A3(KEYINPUT48), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n720), .A2(new_n729), .A3(new_n533), .A4(new_n731), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(new_n760), .A3(G50gat), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n759), .B2(G50gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n761), .A2(new_n762), .A3(new_n756), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n758), .B1(new_n763), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g563(.A(KEYINPUT116), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n665), .A2(new_n607), .A3(new_n685), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n547), .B2(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT116), .B(new_n766), .C1(new_n726), .C2(new_n728), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n527), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g573(.A(KEYINPUT49), .B(G64gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n771), .A2(new_n543), .A3(new_n775), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n770), .A2(new_n689), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1333gat));
  OAI21_X1  g577(.A(G71gat), .B1(new_n770), .B2(new_n334), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n327), .A2(G71gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n771), .A2(new_n533), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g584(.A1(new_n633), .A2(new_n607), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n685), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n730), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n527), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n547), .A2(new_n664), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT51), .B1(new_n791), .B2(new_n786), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NOR4_X1   g592(.A1(new_n547), .A2(new_n793), .A3(new_n664), .A4(new_n787), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n772), .A2(new_n639), .A3(new_n684), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n790), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  NAND4_X1  g596(.A1(new_n720), .A2(new_n729), .A3(new_n543), .A4(new_n788), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G92gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n543), .A2(new_n640), .A3(new_n684), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT52), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  OAI211_X1 g602(.A(new_n803), .B(new_n799), .C1(new_n795), .C2(new_n800), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n789), .B2(new_n334), .ZN(new_n806));
  OR3_X1    g605(.A1(new_n327), .A2(G99gat), .A3(new_n685), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n795), .B2(new_n807), .ZN(G1338gat));
  NAND4_X1  g607(.A1(new_n720), .A2(new_n729), .A3(new_n753), .A4(new_n788), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G106gat), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n425), .A2(new_n685), .A3(G106gat), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n810), .B(new_n811), .C1(new_n795), .C2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n795), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n720), .A2(new_n729), .A3(new_n533), .A4(new_n788), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n815), .A2(new_n812), .B1(G106gat), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(G1339gat));
  NOR4_X1   g618(.A1(new_n632), .A2(new_n721), .A3(new_n607), .A4(new_n684), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n673), .A2(new_n667), .A3(new_n674), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(KEYINPUT54), .A3(new_n675), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n823), .B(new_n667), .C1(new_n673), .C2(new_n674), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n681), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n822), .A2(new_n825), .A3(KEYINPUT55), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n683), .ZN(new_n830));
  INV_X1    g629(.A(new_n606), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n604), .A3(new_n602), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n634), .A2(new_n587), .A3(new_n588), .A4(new_n585), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n583), .B1(new_n833), .B2(new_n582), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n597), .A2(new_n598), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n553), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT118), .B(new_n553), .C1(new_n834), .C2(new_n835), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n721), .A2(new_n828), .A3(new_n830), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n607), .A2(new_n828), .A3(new_n683), .A4(new_n829), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n832), .A2(new_n840), .A3(new_n684), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT119), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n664), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT119), .B1(new_n843), .B2(new_n844), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n820), .B1(new_n848), .B2(new_n632), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(new_n327), .A3(new_n533), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n772), .A3(new_n689), .ZN(new_n851));
  INV_X1    g650(.A(G113gat), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(new_n608), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n849), .A2(new_n527), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n854), .A2(new_n332), .A3(new_n425), .A4(new_n689), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n855), .A2(new_n608), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n853), .B1(new_n852), .B2(new_n856), .ZN(G1340gat));
  INV_X1    g656(.A(G120gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n851), .A2(new_n858), .A3(new_n685), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n855), .A2(new_n685), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n858), .B2(new_n860), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n851), .B2(new_n632), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n633), .A2(new_n624), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n862), .B1(new_n855), .B2(new_n863), .ZN(G1342gat));
  OR3_X1    g663(.A1(new_n855), .A2(G134gat), .A3(new_n664), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n851), .B2(new_n664), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n741), .A2(new_n425), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n870), .A3(new_n689), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n362), .B1(new_n871), .B2(new_n608), .ZN(new_n872));
  OR2_X1    g671(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT55), .B1(new_n822), .B2(new_n825), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n830), .A2(new_n607), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n844), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n664), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n633), .B1(new_n878), .B2(new_n842), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n533), .B1(new_n879), .B2(new_n820), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  INV_X1    g681(.A(new_n847), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n664), .A3(new_n845), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n633), .B1(new_n884), .B2(new_n842), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n882), .B(new_n753), .C1(new_n885), .C2(new_n820), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n741), .A2(new_n527), .A3(new_n543), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n607), .A2(G141gat), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n872), .B(new_n873), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(G1344gat));
  OAI21_X1  g691(.A(KEYINPUT57), .B1(new_n849), .B2(new_n425), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n882), .B(new_n533), .C1(new_n879), .C2(new_n820), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n684), .A3(new_n887), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(G148gat), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT123), .B1(new_n896), .B2(KEYINPUT59), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n898), .B(new_n899), .C1(new_n895), .C2(G148gat), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n881), .A2(new_n886), .A3(new_n684), .A4(new_n887), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n363), .A2(KEYINPUT59), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n902), .A2(new_n901), .A3(new_n903), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n897), .A2(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n871), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n363), .A3(new_n684), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n908), .ZN(G1345gat));
  NOR3_X1   g708(.A1(new_n888), .A2(new_n380), .A3(new_n632), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n633), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  AOI21_X1  g711(.A(G155gat), .B1(new_n911), .B2(KEYINPUT124), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1346gat));
  NAND3_X1  g713(.A1(new_n907), .A2(new_n379), .A3(new_n721), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n374), .B1(new_n888), .B2(new_n664), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n849), .A2(new_n772), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n332), .A2(new_n425), .A3(new_n543), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n607), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n772), .A2(new_n689), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n850), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n924), .A2(new_n249), .A3(new_n608), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n922), .A2(new_n925), .ZN(G1348gat));
  OAI21_X1  g725(.A(new_n266), .B1(new_n920), .B2(new_n685), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n684), .A2(new_n248), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT125), .Z(G1349gat));
  NAND3_X1  g729(.A1(new_n921), .A2(new_n278), .A3(new_n633), .ZN(new_n931));
  OAI21_X1  g730(.A(G183gat), .B1(new_n924), .B2(new_n632), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n921), .A2(new_n206), .A3(new_n721), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n850), .A2(new_n721), .A3(new_n923), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n938), .A3(G190gat), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n938), .B1(new_n937), .B2(G190gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(G1351gat));
  AND2_X1   g741(.A1(new_n893), .A2(new_n894), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n334), .A2(new_n923), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n608), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n741), .A2(new_n425), .A3(new_n689), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(KEYINPUT127), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n948), .A2(new_n918), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n607), .A2(new_n340), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NOR2_X1   g751(.A1(new_n685), .A2(G204gat), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n950), .A2(KEYINPUT62), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT62), .B1(new_n950), .B2(new_n954), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n943), .A2(new_n684), .A3(new_n944), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n955), .B(new_n956), .C1(new_n345), .C2(new_n957), .ZN(G1353gat));
  OR3_X1    g757(.A1(new_n950), .A2(G211gat), .A3(new_n632), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n633), .A3(new_n944), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  OAI21_X1  g762(.A(G218gat), .B1(new_n945), .B2(new_n664), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n664), .A2(G218gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n950), .B2(new_n965), .ZN(G1355gat));
endmodule


