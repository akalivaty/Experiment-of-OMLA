//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1203,
    new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT65), .Z(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(G137), .A3(new_n463), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n463), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n463), .A3(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n474), .A3(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n463), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n478), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT3), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT69), .B1(new_n487), .B2(new_n463), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n467), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n482), .B1(G124), .B2(new_n491), .ZN(G162));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n484), .A2(new_n486), .A3(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n463), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n471), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G102), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n493), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n495), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n501), .B1(new_n467), .B2(G126), .ZN(new_n502));
  OAI211_X1 g077(.A(KEYINPUT70), .B(new_n498), .C1(new_n502), .C2(new_n463), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n484), .A2(new_n486), .A3(G138), .A4(new_n463), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(KEYINPUT71), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n467), .A2(G138), .A3(new_n463), .A4(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n500), .A2(new_n503), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(G166));
  OR2_X1    g102(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(KEYINPUT72), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(G51), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT73), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  INV_X1    g110(.A(new_n522), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n533), .A2(new_n535), .B1(G89), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND2_X1  g116(.A1(new_n528), .A2(new_n529), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT74), .B(G52), .Z(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n545), .A2(new_n519), .B1(new_n546), .B2(new_n522), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n514), .A2(new_n516), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT75), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n519), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n536), .A2(G81), .ZN(new_n555));
  INV_X1    g130(.A(G43), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n542), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  INV_X1    g140(.A(new_n524), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G53), .ZN(new_n567));
  NAND2_X1  g142(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n570), .A2(new_n519), .B1(new_n522), .B2(new_n571), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n569), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(KEYINPUT78), .ZN(new_n575));
  XNOR2_X1  g150(.A(G166), .B(new_n575), .ZN(G303));
  NAND2_X1  g151(.A1(new_n536), .A2(G87), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n566), .A2(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  INV_X1    g156(.A(G48), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n522), .A2(new_n581), .B1(new_n524), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT79), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n514), .A2(new_n516), .A3(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n519), .B1(new_n591), .B2(new_n522), .ZN(new_n592));
  INV_X1    g167(.A(new_n542), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(G47), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(new_n593), .A2(G54), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n517), .A2(G92), .A3(new_n521), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT10), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(new_n519), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G284));
  OAI21_X1  g179(.A(new_n603), .B1(new_n602), .B2(G171), .ZN(G321));
  NAND2_X1  g180(.A1(G299), .A2(new_n602), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(G168), .B2(new_n602), .ZN(G280));
  AND3_X1   g183(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  OAI21_X1  g186(.A(new_n602), .B1(new_n554), .B2(new_n557), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n601), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n491), .A2(G123), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT80), .Z(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n620), .B(new_n621), .C1(G111), .C2(new_n463), .ZN(new_n622));
  INV_X1    g197(.A(new_n478), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G135), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n617), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G2096), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n472), .A2(new_n474), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n628), .A2(new_n487), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n627), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2435), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2438), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n644), .A2(new_n647), .A3(new_n645), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n647), .B1(new_n644), .B2(new_n645), .ZN(new_n649));
  OAI211_X1 g224(.A(G14), .B(new_n646), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT84), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n655), .B(KEYINPUT17), .Z(new_n658));
  OAI21_X1  g233(.A(new_n657), .B1(new_n654), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  INV_X1    g235(.A(new_n652), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n654), .A2(new_n661), .A3(new_n656), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n654), .A3(new_n652), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2096), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n626), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n632), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n670), .A3(G2100), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n680), .B1(KEYINPUT20), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n679), .A3(new_n681), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n683), .B(new_n684), .C1(KEYINPUT20), .C2(new_n682), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT87), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1981), .B(G1986), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n690), .ZN(new_n693));
  AND3_X1   g268(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G24), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n594), .B2(new_n697), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n699), .A2(G1986), .ZN(new_n700));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT32), .ZN(new_n702));
  INV_X1    g277(.A(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n697), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n697), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT89), .B(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n697), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n697), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT33), .Z(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(G1976), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(G1976), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n704), .A2(new_n708), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n491), .A2(G119), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n623), .A2(G131), .ZN(new_n722));
  OR2_X1    g297(.A1(G95), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT35), .B(G1991), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n699), .B2(G1986), .ZN(new_n730));
  AND4_X1   g305(.A1(new_n700), .A2(new_n717), .A3(new_n718), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT90), .B(KEYINPUT36), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n718), .A2(new_n730), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n735), .A2(new_n700), .A3(new_n717), .A4(new_n733), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT91), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n700), .A3(new_n717), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT36), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n734), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g315(.A1(G5), .A2(G16), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G171), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1961), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n719), .A2(G32), .ZN(new_n744));
  INV_X1    g319(.A(new_n628), .ZN(new_n745));
  AOI22_X1  g320(.A1(G141), .A2(new_n623), .B1(new_n745), .B2(G105), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n491), .A2(G129), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT94), .B(KEYINPUT26), .Z(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n744), .B1(new_n752), .B2(new_n719), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n743), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(KEYINPUT24), .A2(G34), .ZN(new_n757));
  NOR2_X1   g332(.A1(KEYINPUT24), .A2(G34), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n757), .A2(new_n758), .A3(G29), .ZN(new_n759));
  INV_X1    g334(.A(G160), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2084), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n719), .A2(G33), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n766), .A2(G2105), .B1(new_n623), .B2(G139), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n497), .A2(G103), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT25), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(new_n719), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT93), .B(G2072), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n697), .A2(G4), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n609), .B2(new_n697), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n774), .B1(new_n776), .B2(G1348), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n753), .A2(new_n755), .B1(new_n762), .B2(new_n761), .ZN(new_n778));
  INV_X1    g353(.A(new_n776), .ZN(new_n779));
  INV_X1    g354(.A(G1348), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n756), .A2(new_n763), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n719), .A2(G26), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n491), .A2(G128), .ZN(new_n784));
  OR2_X1    g359(.A1(G104), .A2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n785), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n786));
  AOI21_X1  g361(.A(KEYINPUT92), .B1(new_n623), .B2(G140), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n788));
  INV_X1    g363(.A(G140), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n478), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n784), .B(new_n786), .C1(new_n787), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n783), .B1(new_n791), .B2(G29), .ZN(new_n792));
  MUX2_X1   g367(.A(new_n783), .B(new_n792), .S(KEYINPUT28), .Z(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT31), .B(G11), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n797));
  AND3_X1   g372(.A1(new_n797), .A2(KEYINPUT95), .A3(G28), .ZN(new_n798));
  AOI21_X1  g373(.A(KEYINPUT95), .B1(new_n797), .B2(G28), .ZN(new_n799));
  OAI221_X1 g374(.A(new_n719), .B1(new_n797), .B2(G28), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n796), .B(new_n800), .C1(new_n625), .C2(new_n719), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT96), .Z(new_n802));
  NOR3_X1   g377(.A1(new_n782), .A2(new_n795), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n697), .A2(G21), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G168), .B2(new_n697), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1966), .ZN(new_n806));
  AND3_X1   g381(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n569), .A2(new_n572), .ZN(new_n808));
  OAI21_X1  g383(.A(KEYINPUT23), .B1(new_n808), .B2(new_n697), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n697), .A2(G20), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n697), .A2(G19), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n558), .B2(new_n697), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n811), .A2(new_n812), .B1(G1341), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n719), .A2(G35), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G162), .B2(new_n719), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT29), .Z(new_n818));
  INV_X1    g393(.A(G2090), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n815), .B(new_n820), .C1(new_n812), .C2(new_n811), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n818), .A2(new_n819), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n719), .A2(G27), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G164), .B2(new_n719), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G2078), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n806), .A2(new_n821), .A3(new_n822), .A4(new_n825), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n803), .B(new_n826), .C1(G1341), .C2(new_n814), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n740), .A2(new_n828), .ZN(G311));
  NAND2_X1  g404(.A1(new_n740), .A2(new_n828), .ZN(G150));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n550), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G651), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT98), .B(G93), .Z(new_n835));
  NAND2_X1  g410(.A1(new_n536), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n836), .C1(new_n542), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n558), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n838), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n557), .B2(new_n554), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n601), .A2(new_n610), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n848), .B(new_n849), .C1(new_n846), .C2(new_n845), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n838), .A2(G860), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT100), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  NAND2_X1  g429(.A1(new_n491), .A2(G130), .ZN(new_n855));
  OR2_X1    g430(.A1(G106), .A2(G2105), .ZN(new_n856));
  INV_X1    g431(.A(G118), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n483), .B1(new_n857), .B2(G2105), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n623), .A2(G142), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n630), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n630), .A2(new_n860), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n726), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n725), .B1(new_n865), .B2(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT101), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n494), .A2(new_n495), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(G2105), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n873), .A2(new_n506), .A3(new_n509), .A4(new_n498), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n791), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n791), .A2(new_n875), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(new_n770), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n770), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n751), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n880), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n752), .A3(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT102), .B1(new_n871), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n869), .A2(new_n870), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n886), .A2(new_n881), .A3(new_n887), .A4(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n871), .A2(new_n884), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n625), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n884), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n881), .A2(new_n883), .A3(KEYINPUT103), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n889), .B(new_n895), .C1(new_n867), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g477(.A(new_n842), .B(KEYINPUT104), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n613), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n609), .A2(G299), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n601), .A2(new_n808), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(KEYINPUT41), .A3(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n908), .B1(new_n913), .B2(new_n904), .ZN(new_n914));
  NOR2_X1   g489(.A1(G290), .A2(new_n710), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n594), .A2(G288), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n915), .A2(KEYINPUT105), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n594), .B(G288), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n919));
  XNOR2_X1  g494(.A(G305), .B(G166), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n914), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n924), .A2(new_n925), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n908), .B(new_n929), .C1(new_n913), .C2(new_n904), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n928), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g507(.A(G868), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n838), .A2(new_n602), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  NAND2_X1  g510(.A1(new_n933), .A2(new_n934), .ZN(G331));
  INV_X1    g511(.A(G37), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n537), .B(new_n539), .C1(G301), .C2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(G171), .A2(KEYINPUT107), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n842), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(G301), .A2(new_n938), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n839), .B2(new_n841), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n939), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n939), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n842), .A2(new_n940), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n839), .A3(new_n841), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n944), .A2(new_n948), .A3(new_n912), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n944), .A2(new_n948), .B1(new_n906), .B2(new_n905), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n921), .A2(new_n922), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n944), .A2(new_n948), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n907), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(new_n948), .A3(new_n912), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n923), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n937), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n949), .B2(new_n950), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n954), .A2(new_n923), .A3(new_n955), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n955), .A2(new_n961), .A3(new_n923), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n954), .A2(new_n961), .A3(new_n923), .A4(new_n955), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n937), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n958), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n957), .A2(new_n964), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n963), .A2(new_n937), .A3(new_n965), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n969), .B2(new_n964), .ZN(new_n970));
  MUX2_X1   g545(.A(new_n967), .B(new_n970), .S(KEYINPUT44), .Z(G397));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n511), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n498), .B1(new_n502), .B2(new_n463), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n506), .A2(new_n509), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n972), .B(new_n973), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n470), .A2(new_n475), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT109), .B(G40), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n465), .B1(G125), .B2(new_n467), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n979), .B(new_n981), .C1(new_n982), .C2(new_n463), .ZN(new_n983));
  NOR4_X1   g558(.A1(new_n974), .A2(new_n978), .A3(G2084), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n989));
  AOI21_X1  g564(.A(G1966), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n984), .A2(new_n985), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n511), .A2(new_n973), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n469), .A2(new_n476), .A3(new_n980), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n993), .A2(new_n762), .A3(new_n994), .A4(new_n977), .ZN(new_n995));
  INV_X1    g570(.A(G1966), .ZN(new_n996));
  AND3_X1   g571(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n496), .A2(new_n499), .ZN(new_n998));
  AOI21_X1  g573(.A(G1384), .B1(new_n510), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n994), .B1(new_n999), .B2(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n996), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT118), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(G168), .B1(new_n991), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n985), .B1(new_n984), .B2(new_n990), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1005), .B1(new_n537), .B2(new_n539), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n995), .A2(new_n1001), .A3(KEYINPUT118), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1003), .A2(KEYINPUT51), .A3(G8), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1006), .A2(KEYINPUT51), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n984), .B2(new_n990), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n972), .B1(new_n874), .B2(new_n973), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n983), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n511), .A2(new_n972), .A3(new_n973), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n994), .B(KEYINPUT114), .C1(new_n999), .C2(new_n972), .ZN(new_n1020));
  AND4_X1   g595(.A1(new_n819), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n983), .B1(new_n992), .B2(new_n987), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n874), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1971), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT115), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1018), .A2(new_n819), .A3(new_n1020), .A4(new_n1019), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT45), .B1(new_n511), .B2(new_n973), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1023), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n983), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1026), .B(new_n1027), .C1(G1971), .C2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1025), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G303), .A2(G8), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(KEYINPUT111), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1033), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n993), .A2(new_n994), .A3(new_n977), .ZN(new_n1042));
  OAI221_X1 g617(.A(KEYINPUT110), .B1(new_n1030), .B2(G1971), .C1(new_n1042), .C2(G2090), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1042), .A2(G2090), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(new_n1024), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1043), .A2(new_n1046), .A3(new_n1039), .A4(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n983), .A2(new_n986), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(new_n1005), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT49), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n584), .A2(new_n703), .A3(new_n588), .ZN(new_n1051));
  INV_X1    g626(.A(new_n588), .ZN(new_n1052));
  OAI21_X1  g627(.A(G1981), .B1(new_n1052), .B2(new_n583), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1054), .B2(new_n1050), .ZN(new_n1056));
  AOI211_X1 g631(.A(KEYINPUT112), .B(KEYINPUT49), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1057));
  OAI221_X1 g632(.A(new_n1049), .B1(new_n1050), .B2(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1976), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1049), .B1(new_n1059), .B2(G288), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT52), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n1059), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1049), .B(new_n1062), .C1(new_n1059), .C2(G288), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1058), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1041), .A2(new_n1047), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G2078), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n986), .A2(new_n987), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n989), .A2(new_n1067), .A3(new_n1068), .A4(new_n994), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n988), .A2(new_n989), .A3(KEYINPUT119), .A4(new_n1067), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1042), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(KEYINPUT121), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(KEYINPUT121), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1080), .B(new_n1081), .C1(new_n1082), .C2(G2078), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1073), .A2(KEYINPUT120), .A3(new_n1075), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1078), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(G171), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1015), .A2(KEYINPUT124), .A3(new_n1066), .A4(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1064), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1089), .A2(G171), .A3(new_n1047), .A4(new_n1085), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT62), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1009), .A2(KEYINPUT62), .A3(new_n1012), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1087), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1058), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n710), .A2(new_n1059), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT113), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1051), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n1049), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1047), .B2(new_n1064), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1043), .A2(new_n1046), .A3(G8), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1064), .B1(new_n1103), .B2(new_n1040), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1011), .A2(G286), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1047), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1105), .A2(KEYINPUT63), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1066), .A2(new_n1106), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1102), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n982), .B(KEYINPUT122), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(G2105), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1115), .A2(KEYINPUT53), .A3(G40), .A4(new_n1067), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1068), .A2(new_n979), .A3(new_n1023), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1083), .B(new_n1075), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT123), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1119), .A2(G301), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1085), .A2(G301), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT54), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1118), .B2(G171), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1120), .A2(new_n1122), .B1(new_n1086), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1082), .A2(G1996), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT58), .B(G1341), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1048), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n558), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n808), .B(KEYINPUT57), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n812), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1030), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1132), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(KEYINPUT61), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(KEYINPUT61), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1131), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT117), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1042), .A2(new_n780), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1048), .A2(new_n794), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1141), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1042), .A2(new_n780), .B1(new_n794), .B2(new_n1048), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1147), .A2(KEYINPUT117), .A3(KEYINPUT60), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1146), .A2(new_n609), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1141), .B(new_n601), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1140), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1132), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1147), .A2(new_n601), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1137), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1013), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1125), .A2(new_n1158), .A3(new_n1066), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1087), .A2(new_n1092), .A3(KEYINPUT125), .A4(new_n1093), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1096), .A2(new_n1113), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1068), .A2(new_n983), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n791), .B(new_n794), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n751), .A2(G1996), .ZN(new_n1164));
  INV_X1    g739(.A(G1996), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n752), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n725), .A2(new_n728), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n725), .A2(new_n728), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(G1986), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1170), .B1(new_n1171), .B2(new_n594), .ZN(new_n1172));
  NOR2_X1   g747(.A1(G290), .A2(G1986), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1162), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1161), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1162), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1163), .B2(new_n752), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1178));
  XNOR2_X1  g753(.A(KEYINPUT126), .B(KEYINPUT46), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(KEYINPUT126), .A2(KEYINPUT46), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT47), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1173), .A2(new_n1162), .ZN(new_n1184));
  XNOR2_X1  g759(.A(new_n1184), .B(KEYINPUT48), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1170), .B2(new_n1176), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1169), .ZN(new_n1187));
  OAI22_X1  g762(.A1(new_n1167), .A2(new_n1187), .B1(G2067), .B2(new_n791), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1162), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1183), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1175), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  OAI21_X1  g768(.A(G319), .B1(new_n694), .B2(new_n695), .ZN(new_n1195));
  INV_X1    g769(.A(new_n1195), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n672), .A2(new_n650), .A3(new_n673), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n894), .B2(new_n900), .ZN(new_n1198));
  AND4_X1   g772(.A1(new_n1194), .A2(new_n967), .A3(new_n1196), .A4(new_n1198), .ZN(new_n1199));
  AOI21_X1  g773(.A(new_n1195), .B1(new_n958), .B2(new_n966), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1194), .B1(new_n1200), .B2(new_n1198), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n1199), .A2(new_n1201), .ZN(G308));
  NAND3_X1  g776(.A1(new_n967), .A2(new_n1198), .A3(new_n1196), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1203), .A2(KEYINPUT127), .ZN(new_n1204));
  NAND3_X1  g778(.A1(new_n1200), .A2(new_n1194), .A3(new_n1198), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1205), .ZN(G225));
endmodule


