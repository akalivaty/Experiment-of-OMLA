

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769;

  XNOR2_X1 U373 ( .A(n495), .B(G134), .ZN(n531) );
  XOR2_X1 U374 ( .A(G116), .B(G107), .Z(n530) );
  AND2_X1 U375 ( .A1(n412), .A2(KEYINPUT44), .ZN(n410) );
  BUF_X1 U376 ( .A(n546), .Z(n582) );
  NOR2_X2 U377 ( .A1(n360), .A2(n683), .ZN(n660) );
  NOR2_X2 U378 ( .A1(n713), .A2(n595), .ZN(n427) );
  XNOR2_X2 U379 ( .A(n586), .B(n585), .ZN(n713) );
  NOR2_X2 U380 ( .A1(n666), .A2(n677), .ZN(n667) );
  INV_X1 U381 ( .A(n464), .ZN(n636) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n516) );
  NOR2_X1 U383 ( .A1(n747), .A2(n399), .ZN(n681) );
  NOR2_X1 U384 ( .A1(n571), .A2(n514), .ZN(n730) );
  INV_X1 U385 ( .A(G146), .ZN(n422) );
  NAND2_X1 U386 ( .A1(n363), .A2(n578), .ZN(n740) );
  XNOR2_X1 U387 ( .A(n609), .B(n608), .ZN(n641) );
  XNOR2_X1 U388 ( .A(n428), .B(n594), .ZN(n623) );
  OR2_X1 U389 ( .A1(n603), .A2(n621), .ZN(n586) );
  OR2_X1 U390 ( .A1(n694), .A2(n693), .ZN(n621) );
  XNOR2_X1 U391 ( .A(n582), .B(KEYINPUT38), .ZN(n566) );
  XNOR2_X1 U392 ( .A(n563), .B(KEYINPUT1), .ZN(n694) );
  XNOR2_X1 U393 ( .A(n655), .B(KEYINPUT59), .ZN(n656) );
  XNOR2_X1 U394 ( .A(n487), .B(n420), .ZN(n648) );
  NOR2_X2 U395 ( .A1(n360), .A2(n683), .ZN(n351) );
  BUF_X1 U396 ( .A(n660), .Z(n671) );
  XNOR2_X1 U397 ( .A(n365), .B(n430), .ZN(n575) );
  INV_X1 U398 ( .A(n385), .ZN(n377) );
  AND2_X1 U399 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U400 ( .A1(n526), .A2(G902), .ZN(n382) );
  NAND2_X1 U401 ( .A1(n364), .A2(n740), .ZN(n365) );
  AND2_X1 U402 ( .A1(n366), .A2(n367), .ZN(n364) );
  NOR2_X1 U403 ( .A1(n352), .A2(n552), .ZN(n366) );
  XNOR2_X1 U404 ( .A(n515), .B(KEYINPUT81), .ZN(n367) );
  INV_X1 U405 ( .A(G234), .ZN(n435) );
  INV_X1 U406 ( .A(KEYINPUT8), .ZN(n444) );
  NAND2_X1 U407 ( .A1(n444), .A2(n435), .ZN(n434) );
  XNOR2_X1 U408 ( .A(n474), .B(n518), .ZN(n423) );
  XNOR2_X1 U409 ( .A(n399), .B(KEYINPUT75), .ZN(n406) );
  INV_X1 U410 ( .A(KEYINPUT2), .ZN(n405) );
  XNOR2_X1 U411 ( .A(n456), .B(G902), .ZN(n631) );
  NOR2_X1 U412 ( .A1(n537), .A2(G902), .ZN(n386) );
  XNOR2_X1 U413 ( .A(n490), .B(n489), .ZN(n563) );
  XNOR2_X1 U414 ( .A(n393), .B(KEYINPUT12), .ZN(n392) );
  XNOR2_X1 U415 ( .A(n395), .B(KEYINPUT102), .ZN(n394) );
  INV_X1 U416 ( .A(KEYINPUT11), .ZN(n395) );
  INV_X1 U417 ( .A(KEYINPUT10), .ZN(n451) );
  XNOR2_X1 U418 ( .A(G113), .B(G143), .ZN(n519) );
  XNOR2_X1 U419 ( .A(KEYINPUT18), .B(KEYINPUT78), .ZN(n494) );
  XNOR2_X1 U420 ( .A(G146), .B(G125), .ZN(n499) );
  XNOR2_X1 U421 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n498) );
  XNOR2_X1 U422 ( .A(n506), .B(n437), .ZN(n753) );
  XNOR2_X1 U423 ( .A(n505), .B(n504), .ZN(n437) );
  INV_X1 U424 ( .A(KEYINPUT16), .ZN(n503) );
  XNOR2_X1 U425 ( .A(n570), .B(n402), .ZN(n714) );
  INV_X1 U426 ( .A(KEYINPUT41), .ZN(n402) );
  NOR2_X1 U427 ( .A1(n564), .A2(n415), .ZN(n414) );
  NAND2_X1 U428 ( .A1(n566), .A2(KEYINPUT39), .ZN(n415) );
  NAND2_X1 U429 ( .A1(n688), .A2(n419), .ZN(n417) );
  AND2_X1 U430 ( .A1(n378), .A2(n373), .ZN(n372) );
  AND2_X1 U431 ( .A1(n381), .A2(n370), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n398), .B(n397), .ZN(n396) );
  INV_X1 U433 ( .A(KEYINPUT72), .ZN(n397) );
  NAND2_X1 U434 ( .A1(n686), .A2(n551), .ZN(n398) );
  INV_X1 U435 ( .A(KEYINPUT69), .ZN(n430) );
  NOR2_X1 U436 ( .A1(n597), .A2(KEYINPUT65), .ZN(n610) );
  INV_X1 U437 ( .A(n646), .ZN(n409) );
  NAND2_X1 U438 ( .A1(n557), .A2(n736), .ZN(n686) );
  NAND2_X1 U439 ( .A1(n537), .A2(G902), .ZN(n389) );
  XNOR2_X1 U440 ( .A(G119), .B(G137), .ZN(n445) );
  NAND2_X1 U441 ( .A1(G234), .A2(G237), .ZN(n462) );
  XOR2_X1 U442 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n463) );
  INV_X1 U443 ( .A(G237), .ZN(n508) );
  NOR2_X1 U444 ( .A1(n377), .A2(n371), .ZN(n370) );
  NAND2_X1 U445 ( .A1(n379), .A2(n538), .ZN(n371) );
  NOR2_X1 U446 ( .A1(n377), .A2(n376), .ZN(n375) );
  NAND2_X1 U447 ( .A1(n388), .A2(KEYINPUT106), .ZN(n378) );
  INV_X1 U448 ( .A(n388), .ZN(n387) );
  XNOR2_X1 U449 ( .A(n506), .B(n421), .ZN(n420) );
  XNOR2_X1 U450 ( .A(n477), .B(n480), .ZN(n421) );
  NAND2_X1 U451 ( .A1(n433), .A2(n431), .ZN(n527) );
  NAND2_X1 U452 ( .A1(n636), .A2(n432), .ZN(n431) );
  INV_X1 U453 ( .A(KEYINPUT7), .ZN(n532) );
  NAND2_X1 U454 ( .A1(n361), .A2(n404), .ZN(n360) );
  INV_X1 U455 ( .A(n631), .ZN(n404) );
  NAND2_X1 U456 ( .A1(n362), .A2(n405), .ZN(n361) );
  XNOR2_X1 U457 ( .A(n392), .B(n394), .ZN(n517) );
  XOR2_X1 U458 ( .A(G101), .B(G140), .Z(n484) );
  XNOR2_X1 U459 ( .A(n507), .B(n753), .ZN(n663) );
  XOR2_X1 U460 ( .A(KEYINPUT89), .B(n637), .Z(n677) );
  INV_X1 U461 ( .A(KEYINPUT42), .ZN(n400) );
  OR2_X2 U462 ( .A1(n714), .A2(n571), .ZN(n401) );
  NOR2_X1 U463 ( .A1(n413), .A2(n416), .ZN(n565) );
  OR2_X1 U464 ( .A1(n414), .A2(n557), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n562), .B(KEYINPUT36), .ZN(n363) );
  INV_X1 U466 ( .A(n566), .ZN(n688) );
  INV_X1 U467 ( .A(G902), .ZN(n536) );
  AND2_X1 U468 ( .A1(n730), .A2(n396), .ZN(n352) );
  XOR2_X1 U469 ( .A(n450), .B(n449), .Z(n353) );
  OR2_X1 U470 ( .A1(n414), .A2(n416), .ZN(n354) );
  AND2_X1 U471 ( .A1(n643), .A2(n626), .ZN(n355) );
  AND2_X1 U472 ( .A1(n694), .A2(n619), .ZN(n356) );
  INV_X1 U473 ( .A(KEYINPUT39), .ZN(n419) );
  OR2_X1 U474 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n357) );
  XNOR2_X1 U475 ( .A(n496), .B(n497), .ZN(n502) );
  NOR2_X1 U476 ( .A1(n679), .A2(n358), .ZN(n359) );
  NAND2_X1 U477 ( .A1(n680), .A2(KEYINPUT2), .ZN(n358) );
  XNOR2_X1 U478 ( .A(n630), .B(KEYINPUT45), .ZN(n679) );
  XNOR2_X2 U479 ( .A(n359), .B(KEYINPUT76), .ZN(n683) );
  NAND2_X1 U480 ( .A1(n407), .A2(n406), .ZN(n362) );
  OR2_X1 U481 ( .A1(n669), .A2(n391), .ZN(n390) );
  OR2_X1 U482 ( .A1(n655), .A2(n384), .ZN(n383) );
  NAND2_X1 U483 ( .A1(n381), .A2(n379), .ZN(n545) );
  NAND2_X1 U484 ( .A1(n387), .A2(n385), .ZN(n569) );
  NAND2_X1 U485 ( .A1(n372), .A2(n368), .ZN(n557) );
  NAND2_X1 U486 ( .A1(n369), .A2(n387), .ZN(n368) );
  NAND2_X1 U487 ( .A1(n374), .A2(KEYINPUT106), .ZN(n373) );
  NAND2_X1 U488 ( .A1(n381), .A2(n375), .ZN(n374) );
  INV_X1 U489 ( .A(n379), .ZN(n376) );
  NAND2_X1 U490 ( .A1(n655), .A2(n380), .ZN(n379) );
  NOR2_X1 U491 ( .A1(n526), .A2(G902), .ZN(n380) );
  INV_X1 U492 ( .A(n526), .ZN(n384) );
  NAND2_X1 U493 ( .A1(n669), .A2(n386), .ZN(n385) );
  NAND2_X1 U494 ( .A1(n390), .A2(n389), .ZN(n388) );
  INV_X1 U495 ( .A(n537), .ZN(n391) );
  NAND2_X1 U496 ( .A1(n516), .A2(G214), .ZN(n393) );
  NAND2_X1 U497 ( .A1(n633), .A2(n632), .ZN(n399) );
  XNOR2_X2 U498 ( .A(n576), .B(KEYINPUT48), .ZN(n633) );
  NOR2_X1 U499 ( .A1(n768), .A2(n769), .ZN(n573) );
  XNOR2_X2 U500 ( .A(n401), .B(n400), .ZN(n769) );
  XNOR2_X2 U501 ( .A(n403), .B(G119), .ZN(n439) );
  XNOR2_X2 U502 ( .A(G116), .B(KEYINPUT3), .ZN(n403) );
  INV_X1 U503 ( .A(n679), .ZN(n407) );
  NAND2_X1 U504 ( .A1(n408), .A2(n357), .ZN(n627) );
  NAND2_X1 U505 ( .A1(n410), .A2(n409), .ZN(n408) );
  XNOR2_X2 U506 ( .A(n411), .B(KEYINPUT35), .ZN(n646) );
  NAND2_X1 U507 ( .A1(n426), .A2(n596), .ZN(n411) );
  NAND2_X1 U508 ( .A1(n612), .A2(n611), .ZN(n412) );
  NAND2_X1 U509 ( .A1(n593), .A2(n592), .ZN(n428) );
  NAND2_X1 U510 ( .A1(n418), .A2(n417), .ZN(n416) );
  NAND2_X1 U511 ( .A1(n564), .A2(n419), .ZN(n418) );
  NAND2_X1 U512 ( .A1(n544), .A2(n616), .ZN(n564) );
  XNOR2_X2 U513 ( .A(n440), .B(n439), .ZN(n506) );
  XNOR2_X2 U514 ( .A(n759), .B(n422), .ZN(n487) );
  XNOR2_X2 U515 ( .A(n531), .B(n423), .ZN(n759) );
  XNOR2_X2 U516 ( .A(n425), .B(n424), .ZN(n440) );
  XNOR2_X2 U517 ( .A(G101), .B(KEYINPUT71), .ZN(n424) );
  XNOR2_X2 U518 ( .A(KEYINPUT91), .B(G113), .ZN(n425) );
  XNOR2_X1 U519 ( .A(n427), .B(KEYINPUT34), .ZN(n426) );
  XNOR2_X2 U520 ( .A(n560), .B(n513), .ZN(n593) );
  NAND2_X1 U521 ( .A1(n559), .A2(n429), .ZN(n577) );
  INV_X1 U522 ( .A(n558), .ZN(n429) );
  NAND2_X1 U523 ( .A1(n730), .A2(n429), .ZN(n731) );
  NOR2_X1 U524 ( .A1(n444), .A2(n435), .ZN(n432) );
  AND2_X1 U525 ( .A1(n436), .A2(n434), .ZN(n433) );
  NAND2_X1 U526 ( .A1(n464), .A2(n444), .ZN(n436) );
  XNOR2_X2 U527 ( .A(G953), .B(KEYINPUT64), .ZN(n464) );
  XNOR2_X2 U528 ( .A(n438), .B(G104), .ZN(n505) );
  XNOR2_X2 U529 ( .A(G110), .B(G107), .ZN(n438) );
  NAND2_X2 U530 ( .A1(n441), .A2(n579), .ZN(n560) );
  INV_X1 U531 ( .A(n546), .ZN(n441) );
  XNOR2_X2 U532 ( .A(n510), .B(n509), .ZN(n546) );
  NAND2_X1 U533 ( .A1(n606), .A2(n694), .ZN(n613) );
  NAND2_X1 U534 ( .A1(n606), .A2(n356), .ZN(n601) );
  XNOR2_X1 U535 ( .A(n487), .B(n486), .ZN(n674) );
  XNOR2_X1 U536 ( .A(n505), .B(n485), .ZN(n486) );
  AND2_X1 U537 ( .A1(n554), .A2(n700), .ZN(n482) );
  BUF_X1 U538 ( .A(n679), .Z(n747) );
  XNOR2_X2 U539 ( .A(KEYINPUT68), .B(G131), .ZN(n518) );
  NOR2_X1 U540 ( .A1(n569), .A2(n568), .ZN(n442) );
  AND2_X1 U541 ( .A1(n639), .A2(n638), .ZN(G66) );
  INV_X1 U542 ( .A(KEYINPUT46), .ZN(n572) );
  XNOR2_X1 U543 ( .A(n533), .B(n532), .ZN(n534) );
  INV_X1 U544 ( .A(n677), .ZN(n638) );
  NAND2_X1 U545 ( .A1(G221), .A2(n527), .ZN(n455) );
  XOR2_X1 U546 ( .A(G110), .B(G128), .Z(n446) );
  XNOR2_X1 U547 ( .A(n446), .B(n445), .ZN(n450) );
  XOR2_X1 U548 ( .A(KEYINPUT24), .B(KEYINPUT82), .Z(n448) );
  XNOR2_X1 U549 ( .A(KEYINPUT23), .B(KEYINPUT94), .ZN(n447) );
  XNOR2_X1 U550 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U551 ( .A(n451), .B(G140), .ZN(n452) );
  XNOR2_X1 U552 ( .A(n499), .B(n452), .ZN(n758) );
  INV_X1 U553 ( .A(n758), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n353), .B(n453), .ZN(n454) );
  XNOR2_X1 U555 ( .A(n455), .B(n454), .ZN(n634) );
  NAND2_X1 U556 ( .A1(n634), .A2(n536), .ZN(n461) );
  XOR2_X1 U557 ( .A(KEYINPUT25), .B(KEYINPUT95), .Z(n459) );
  XNOR2_X1 U558 ( .A(KEYINPUT90), .B(KEYINPUT15), .ZN(n456) );
  NAND2_X1 U559 ( .A1(n631), .A2(G234), .ZN(n457) );
  XNOR2_X1 U560 ( .A(KEYINPUT20), .B(n457), .ZN(n470) );
  AND2_X1 U561 ( .A1(n470), .A2(G217), .ZN(n458) );
  XNOR2_X1 U562 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X2 U563 ( .A(n461), .B(n460), .ZN(n696) );
  XNOR2_X1 U564 ( .A(n463), .B(n462), .ZN(n465) );
  NAND2_X1 U565 ( .A1(G952), .A2(n465), .ZN(n712) );
  NOR2_X1 U566 ( .A1(n712), .A2(G953), .ZN(n589) );
  NAND2_X1 U567 ( .A1(n465), .A2(G902), .ZN(n466) );
  XOR2_X1 U568 ( .A(KEYINPUT92), .B(n466), .Z(n588) );
  NAND2_X1 U569 ( .A1(n464), .A2(n588), .ZN(n467) );
  NOR2_X1 U570 ( .A1(G900), .A2(n467), .ZN(n468) );
  XNOR2_X1 U571 ( .A(n468), .B(KEYINPUT108), .ZN(n469) );
  NOR2_X1 U572 ( .A1(n589), .A2(n469), .ZN(n542) );
  AND2_X1 U573 ( .A1(n470), .A2(G221), .ZN(n471) );
  XNOR2_X1 U574 ( .A(n471), .B(KEYINPUT21), .ZN(n697) );
  INV_X1 U575 ( .A(n697), .ZN(n472) );
  OR2_X1 U576 ( .A1(n542), .A2(n472), .ZN(n473) );
  NOR2_X1 U577 ( .A1(n696), .A2(n473), .ZN(n554) );
  XNOR2_X2 U578 ( .A(G143), .B(G128), .ZN(n495) );
  XNOR2_X1 U579 ( .A(G137), .B(KEYINPUT4), .ZN(n474) );
  XOR2_X1 U580 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n476) );
  NAND2_X1 U581 ( .A1(n516), .A2(G210), .ZN(n475) );
  XNOR2_X1 U582 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U583 ( .A(KEYINPUT98), .B(KEYINPUT74), .Z(n479) );
  XNOR2_X1 U584 ( .A(KEYINPUT101), .B(KEYINPUT100), .ZN(n478) );
  XNOR2_X1 U585 ( .A(n479), .B(n478), .ZN(n480) );
  NAND2_X1 U586 ( .A1(n648), .A2(n536), .ZN(n481) );
  XNOR2_X2 U587 ( .A(n481), .B(G472), .ZN(n700) );
  XNOR2_X1 U588 ( .A(n482), .B(KEYINPUT28), .ZN(n492) );
  NAND2_X1 U589 ( .A1(G227), .A2(n636), .ZN(n483) );
  XNOR2_X1 U590 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U591 ( .A1(n674), .A2(n536), .ZN(n490) );
  INV_X1 U592 ( .A(KEYINPUT70), .ZN(n488) );
  XNOR2_X1 U593 ( .A(n488), .B(G469), .ZN(n489) );
  INV_X1 U594 ( .A(n563), .ZN(n491) );
  NAND2_X1 U595 ( .A1(n492), .A2(n491), .ZN(n571) );
  INV_X1 U596 ( .A(G224), .ZN(n493) );
  NOR2_X1 U597 ( .A1(n464), .A2(n493), .ZN(n497) );
  XNOR2_X1 U598 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U599 ( .A(n498), .B(KEYINPUT87), .ZN(n500) );
  XNOR2_X1 U600 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U601 ( .A(n502), .B(n501), .ZN(n507) );
  XNOR2_X1 U602 ( .A(n503), .B(G122), .ZN(n504) );
  NAND2_X1 U603 ( .A1(n663), .A2(n631), .ZN(n510) );
  NAND2_X1 U604 ( .A1(n536), .A2(n508), .ZN(n511) );
  NAND2_X1 U605 ( .A1(n511), .A2(G210), .ZN(n509) );
  NAND2_X1 U606 ( .A1(n511), .A2(G214), .ZN(n579) );
  INV_X1 U607 ( .A(n579), .ZN(n687) );
  INV_X1 U608 ( .A(KEYINPUT77), .ZN(n512) );
  XNOR2_X1 U609 ( .A(n512), .B(KEYINPUT19), .ZN(n513) );
  INV_X1 U610 ( .A(n593), .ZN(n514) );
  INV_X1 U611 ( .A(KEYINPUT47), .ZN(n550) );
  NOR2_X1 U612 ( .A1(n730), .A2(n550), .ZN(n515) );
  XNOR2_X1 U613 ( .A(n518), .B(n517), .ZN(n523) );
  XOR2_X1 U614 ( .A(G122), .B(G104), .Z(n520) );
  XNOR2_X1 U615 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U616 ( .A(n521), .B(n758), .Z(n522) );
  XNOR2_X1 U617 ( .A(n523), .B(n522), .ZN(n655) );
  XOR2_X1 U618 ( .A(KEYINPUT13), .B(KEYINPUT103), .Z(n525) );
  XNOR2_X1 U619 ( .A(KEYINPUT104), .B(G475), .ZN(n524) );
  XNOR2_X1 U620 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U621 ( .A(G122), .B(KEYINPUT9), .Z(n529) );
  NAND2_X1 U622 ( .A1(G217), .A2(n527), .ZN(n528) );
  XNOR2_X1 U623 ( .A(n529), .B(n528), .ZN(n535) );
  XNOR2_X1 U624 ( .A(n531), .B(n530), .ZN(n533) );
  XNOR2_X1 U625 ( .A(n535), .B(n534), .ZN(n669) );
  XOR2_X1 U626 ( .A(KEYINPUT105), .B(G478), .Z(n537) );
  INV_X1 U627 ( .A(KEYINPUT106), .ZN(n538) );
  NAND2_X1 U628 ( .A1(n569), .A2(n545), .ZN(n736) );
  NOR2_X1 U629 ( .A1(n686), .A2(n550), .ZN(n549) );
  NAND2_X1 U630 ( .A1(n700), .A2(n579), .ZN(n540) );
  XOR2_X1 U631 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n539) );
  XOR2_X1 U632 ( .A(n540), .B(n539), .Z(n541) );
  NOR2_X1 U633 ( .A1(n542), .A2(n541), .ZN(n544) );
  NAND2_X1 U634 ( .A1(n696), .A2(n697), .ZN(n693) );
  NOR2_X1 U635 ( .A1(n693), .A2(n563), .ZN(n543) );
  XNOR2_X1 U636 ( .A(n543), .B(KEYINPUT96), .ZN(n616) );
  INV_X1 U637 ( .A(n545), .ZN(n568) );
  AND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n596) );
  INV_X1 U639 ( .A(n582), .ZN(n547) );
  NAND2_X1 U640 ( .A1(n596), .A2(n547), .ZN(n548) );
  NOR2_X1 U641 ( .A1(n564), .A2(n548), .ZN(n640) );
  OR2_X1 U642 ( .A1(n549), .A2(n640), .ZN(n552) );
  XOR2_X1 U643 ( .A(KEYINPUT67), .B(n550), .Z(n551) );
  INV_X1 U644 ( .A(KEYINPUT6), .ZN(n553) );
  XNOR2_X1 U645 ( .A(n700), .B(n553), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n554), .A2(n584), .ZN(n555) );
  XNOR2_X1 U647 ( .A(n555), .B(KEYINPUT109), .ZN(n559) );
  INV_X1 U648 ( .A(KEYINPUT107), .ZN(n556) );
  XNOR2_X1 U649 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U650 ( .A(KEYINPUT112), .B(n577), .ZN(n561) );
  NOR2_X1 U651 ( .A1(n561), .A2(n560), .ZN(n562) );
  INV_X1 U652 ( .A(n694), .ZN(n578) );
  XNOR2_X1 U653 ( .A(n565), .B(KEYINPUT40), .ZN(n768) );
  NAND2_X1 U654 ( .A1(n566), .A2(n579), .ZN(n567) );
  XNOR2_X1 U655 ( .A(n567), .B(KEYINPUT111), .ZN(n685) );
  NAND2_X1 U656 ( .A1(n685), .A2(n442), .ZN(n570) );
  XNOR2_X1 U657 ( .A(n573), .B(n572), .ZN(n574) );
  NOR2_X2 U658 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U659 ( .A1(n354), .A2(n736), .ZN(n742) );
  NOR2_X1 U660 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U662 ( .A(n581), .B(KEYINPUT43), .ZN(n583) );
  AND2_X1 U663 ( .A1(n583), .A2(n582), .ZN(n642) );
  NOR2_X1 U664 ( .A1(n742), .A2(n642), .ZN(n632) );
  INV_X1 U665 ( .A(n584), .ZN(n603) );
  INV_X1 U666 ( .A(KEYINPUT33), .ZN(n585) );
  INV_X1 U667 ( .A(G953), .ZN(n587) );
  NOR2_X1 U668 ( .A1(G898), .A2(n587), .ZN(n751) );
  NAND2_X1 U669 ( .A1(n588), .A2(n751), .ZN(n591) );
  INV_X1 U670 ( .A(n589), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U672 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n594) );
  XNOR2_X1 U673 ( .A(n623), .B(KEYINPUT93), .ZN(n617) );
  INV_X1 U674 ( .A(n617), .ZN(n595) );
  NOR2_X1 U675 ( .A1(n646), .A2(KEYINPUT44), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n442), .A2(n697), .ZN(n598) );
  OR2_X2 U677 ( .A1(n623), .A2(n598), .ZN(n600) );
  INV_X1 U678 ( .A(KEYINPUT22), .ZN(n599) );
  XNOR2_X2 U679 ( .A(n600), .B(n599), .ZN(n606) );
  INV_X1 U680 ( .A(n700), .ZN(n619) );
  XNOR2_X1 U681 ( .A(n601), .B(KEYINPUT66), .ZN(n602) );
  OR2_X2 U682 ( .A1(n602), .A2(n696), .ZN(n645) );
  OR2_X1 U683 ( .A1(n694), .A2(n696), .ZN(n604) );
  NOR2_X1 U684 ( .A1(n604), .A2(n584), .ZN(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n609) );
  INV_X1 U686 ( .A(KEYINPUT79), .ZN(n607) );
  XNOR2_X1 U687 ( .A(n607), .B(KEYINPUT32), .ZN(n608) );
  NAND2_X2 U688 ( .A1(n645), .A2(n641), .ZN(n612) );
  NOR2_X1 U689 ( .A1(n610), .A2(n612), .ZN(n629) );
  INV_X1 U690 ( .A(KEYINPUT65), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n613), .A2(n584), .ZN(n614) );
  XNOR2_X1 U692 ( .A(n614), .B(KEYINPUT84), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n615), .A2(n696), .ZN(n643) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n618), .B(KEYINPUT97), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n723) );
  INV_X1 U697 ( .A(n621), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n622), .A2(n700), .ZN(n704) );
  NOR2_X1 U699 ( .A1(n704), .A2(n623), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n624), .B(KEYINPUT31), .ZN(n735) );
  NAND2_X1 U701 ( .A1(n723), .A2(n735), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n625), .A2(n686), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n355), .ZN(n628) );
  NOR2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  AND2_X2 U705 ( .A1(n633), .A2(n632), .ZN(n680) );
  NAND2_X1 U706 ( .A1(n671), .A2(G217), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n635), .B(n634), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n636), .A2(G952), .ZN(n637) );
  XOR2_X1 U709 ( .A(G143), .B(n640), .Z(G45) );
  XNOR2_X1 U710 ( .A(n641), .B(G119), .ZN(G21) );
  XOR2_X1 U711 ( .A(n642), .B(G140), .Z(G42) );
  XNOR2_X1 U712 ( .A(n643), .B(G101), .ZN(G3) );
  XNOR2_X1 U713 ( .A(G110), .B(KEYINPUT114), .ZN(n644) );
  XNOR2_X1 U714 ( .A(n645), .B(n644), .ZN(G12) );
  XOR2_X1 U715 ( .A(n646), .B(G122), .Z(G24) );
  NAND2_X1 U716 ( .A1(n351), .A2(G472), .ZN(n650) );
  XNOR2_X1 U717 ( .A(KEYINPUT113), .B(KEYINPUT62), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X2 U720 ( .A1(n651), .A2(n677), .ZN(n654) );
  XNOR2_X1 U721 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n652) );
  XNOR2_X1 U722 ( .A(n652), .B(KEYINPUT85), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n654), .B(n653), .ZN(G57) );
  NAND2_X1 U724 ( .A1(n351), .A2(G475), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n658) );
  NOR2_X2 U726 ( .A1(n658), .A2(n677), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n659), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U728 ( .A1(n660), .A2(G210), .ZN(n665) );
  XNOR2_X1 U729 ( .A(KEYINPUT80), .B(KEYINPUT54), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT55), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n667), .B(KEYINPUT56), .ZN(G51) );
  AND2_X1 U734 ( .A1(n671), .A2(G478), .ZN(n668) );
  XNOR2_X1 U735 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U736 ( .A1(n670), .A2(n677), .ZN(G63) );
  NAND2_X1 U737 ( .A1(n671), .A2(G469), .ZN(n676) );
  XNOR2_X1 U738 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT58), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U741 ( .A(n676), .B(n675), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(G54) );
  NOR2_X1 U743 ( .A1(n681), .A2(KEYINPUT2), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n684), .B(KEYINPUT83), .ZN(n720) );
  NAND2_X1 U746 ( .A1(n686), .A2(n685), .ZN(n691) );
  NAND2_X1 U747 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U748 ( .A1(n689), .A2(n442), .ZN(n690) );
  AND2_X1 U749 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U750 ( .A1(n692), .A2(n713), .ZN(n709) );
  NAND2_X1 U751 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U752 ( .A(KEYINPUT50), .B(n695), .ZN(n702) );
  NOR2_X1 U753 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U754 ( .A(KEYINPUT49), .B(n698), .Z(n699) );
  NOR2_X1 U755 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(KEYINPUT120), .ZN(n705) );
  NAND2_X1 U758 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U759 ( .A(KEYINPUT51), .B(n706), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n707), .A2(n714), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U762 ( .A(n710), .B(KEYINPUT52), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U764 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U765 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U766 ( .A(n717), .B(KEYINPUT121), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n718), .A2(G953), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U769 ( .A(KEYINPUT53), .B(n721), .Z(G75) );
  NOR2_X1 U770 ( .A1(n558), .A2(n723), .ZN(n722) );
  XOR2_X1 U771 ( .A(G104), .B(n722), .Z(G6) );
  NOR2_X1 U772 ( .A1(n736), .A2(n723), .ZN(n725) );
  XNOR2_X1 U773 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U775 ( .A(G107), .B(n726), .ZN(G9) );
  XOR2_X1 U776 ( .A(G128), .B(KEYINPUT29), .Z(n729) );
  INV_X1 U777 ( .A(n736), .ZN(n727) );
  NAND2_X1 U778 ( .A1(n730), .A2(n727), .ZN(n728) );
  XNOR2_X1 U779 ( .A(n729), .B(n728), .ZN(G30) );
  XOR2_X1 U780 ( .A(G146), .B(KEYINPUT115), .Z(n732) );
  XNOR2_X1 U781 ( .A(n732), .B(n731), .ZN(G48) );
  NOR2_X1 U782 ( .A1(n558), .A2(n735), .ZN(n733) );
  XOR2_X1 U783 ( .A(KEYINPUT116), .B(n733), .Z(n734) );
  XNOR2_X1 U784 ( .A(G113), .B(n734), .ZN(G15) );
  NOR2_X1 U785 ( .A1(n736), .A2(n735), .ZN(n738) );
  XNOR2_X1 U786 ( .A(G116), .B(KEYINPUT117), .ZN(n737) );
  XNOR2_X1 U787 ( .A(n738), .B(n737), .ZN(G18) );
  XOR2_X1 U788 ( .A(KEYINPUT118), .B(KEYINPUT37), .Z(n739) );
  XNOR2_X1 U789 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U790 ( .A(G125), .B(n741), .ZN(G27) );
  XNOR2_X1 U791 ( .A(G134), .B(n742), .ZN(n743) );
  XNOR2_X1 U792 ( .A(n743), .B(KEYINPUT119), .ZN(G36) );
  NAND2_X1 U793 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U794 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U795 ( .A1(n745), .A2(G898), .ZN(n746) );
  XNOR2_X1 U796 ( .A(KEYINPUT123), .B(n746), .ZN(n750) );
  NOR2_X1 U797 ( .A1(n747), .A2(G953), .ZN(n748) );
  XNOR2_X1 U798 ( .A(n748), .B(KEYINPUT124), .ZN(n749) );
  NOR2_X1 U799 ( .A1(n750), .A2(n749), .ZN(n757) );
  XNOR2_X1 U800 ( .A(KEYINPUT125), .B(KEYINPUT126), .ZN(n755) );
  INV_X1 U801 ( .A(n751), .ZN(n752) );
  NAND2_X1 U802 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U803 ( .A(n755), .B(n754), .Z(n756) );
  XNOR2_X1 U804 ( .A(n757), .B(n756), .ZN(G69) );
  XOR2_X1 U805 ( .A(n759), .B(n758), .Z(n763) );
  INV_X1 U806 ( .A(n763), .ZN(n760) );
  XOR2_X1 U807 ( .A(n760), .B(n399), .Z(n761) );
  NOR2_X1 U808 ( .A1(n464), .A2(n761), .ZN(n762) );
  XNOR2_X1 U809 ( .A(KEYINPUT127), .B(n762), .ZN(n767) );
  XOR2_X1 U810 ( .A(G227), .B(n763), .Z(n764) );
  NAND2_X1 U811 ( .A1(n764), .A2(G900), .ZN(n765) );
  NAND2_X1 U812 ( .A1(n765), .A2(G953), .ZN(n766) );
  NAND2_X1 U813 ( .A1(n767), .A2(n766), .ZN(G72) );
  XOR2_X1 U814 ( .A(G131), .B(n768), .Z(G33) );
  XOR2_X1 U815 ( .A(G137), .B(n769), .Z(G39) );
endmodule

