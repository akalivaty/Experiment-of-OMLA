

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  XOR2_X1 U325 ( .A(n352), .B(n351), .Z(n530) );
  XNOR2_X1 U326 ( .A(n447), .B(n446), .ZN(n449) );
  XNOR2_X1 U327 ( .A(n477), .B(KEYINPUT64), .ZN(n478) );
  XOR2_X1 U328 ( .A(n352), .B(n309), .Z(n539) );
  NOR2_X1 U329 ( .A1(n584), .A2(n588), .ZN(n293) );
  XOR2_X1 U330 ( .A(G204GAT), .B(KEYINPUT75), .Z(n294) );
  INV_X1 U331 ( .A(KEYINPUT98), .ZN(n336) );
  XNOR2_X1 U332 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U333 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U334 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U335 ( .A(n450), .B(n294), .ZN(n451) );
  OR2_X1 U336 ( .A1(n539), .A2(n537), .ZN(n378) );
  XNOR2_X1 U337 ( .A(n452), .B(n451), .ZN(n456) );
  XNOR2_X1 U338 ( .A(n479), .B(n478), .ZN(n538) );
  XOR2_X1 U339 ( .A(KEYINPUT38), .B(n460), .Z(n512) );
  XNOR2_X1 U340 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U341 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U342 ( .A(n493), .B(n492), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n464), .B(n463), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n296) );
  XNOR2_X1 U345 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n295) );
  XNOR2_X1 U346 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U347 ( .A(G169GAT), .B(n297), .Z(n352) );
  XOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .Z(n319) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n454) );
  XOR2_X1 U350 ( .A(n319), .B(n454), .Z(n299) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G127GAT), .Z(n388) );
  XOR2_X1 U354 ( .A(n300), .B(n388), .Z(n308) );
  XOR2_X1 U355 ( .A(G99GAT), .B(G134GAT), .Z(n302) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U358 ( .A(G176GAT), .B(G183GAT), .Z(n304) );
  XNOR2_X1 U359 ( .A(KEYINPUT20), .B(KEYINPUT85), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U363 ( .A(KEYINPUT4), .B(G57GAT), .Z(n311) );
  XNOR2_X1 U364 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n310) );
  XNOR2_X1 U365 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U366 ( .A(KEYINPUT1), .B(KEYINPUT95), .Z(n313) );
  XNOR2_X1 U367 ( .A(KEYINPUT96), .B(KEYINPUT5), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U369 ( .A(n315), .B(n314), .Z(n321) );
  XOR2_X1 U370 ( .A(G134GAT), .B(KEYINPUT79), .Z(n412) );
  XOR2_X1 U371 ( .A(KEYINPUT6), .B(n412), .Z(n317) );
  NAND2_X1 U372 ( .A1(G225GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G162GAT), .Z(n323) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(G148GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U379 ( .A(n325), .B(n324), .Z(n333) );
  XOR2_X1 U380 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U383 ( .A(G141GAT), .B(n328), .Z(n364) );
  XOR2_X1 U384 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n330) );
  XNOR2_X1 U385 ( .A(G127GAT), .B(G120GAT), .ZN(n329) );
  XNOR2_X1 U386 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n364), .B(n331), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n528) );
  INV_X1 U389 ( .A(n539), .ZN(n488) );
  XOR2_X1 U390 ( .A(KEYINPUT102), .B(KEYINPUT100), .Z(n335) );
  XNOR2_X1 U391 ( .A(KEYINPUT97), .B(KEYINPUT101), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n339) );
  NAND2_X1 U393 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XOR2_X1 U394 ( .A(n340), .B(KEYINPUT99), .Z(n346) );
  XNOR2_X1 U395 ( .A(G211GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n341), .B(KEYINPUT89), .ZN(n342) );
  XOR2_X1 U397 ( .A(n342), .B(KEYINPUT21), .Z(n344) );
  XNOR2_X1 U398 ( .A(G197GAT), .B(G204GAT), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n365) );
  XNOR2_X1 U400 ( .A(n365), .B(G92GAT), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(G8GAT), .B(G183GAT), .Z(n381) );
  XOR2_X1 U403 ( .A(n347), .B(n381), .Z(n350) );
  XOR2_X1 U404 ( .A(G176GAT), .B(G64GAT), .Z(n448) );
  XNOR2_X1 U405 ( .A(G36GAT), .B(G190GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n348), .B(KEYINPUT80), .ZN(n416) );
  XNOR2_X1 U407 ( .A(n448), .B(n416), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  INV_X1 U409 ( .A(n530), .ZN(n480) );
  NOR2_X1 U410 ( .A1(n488), .A2(n480), .ZN(n353) );
  XNOR2_X1 U411 ( .A(KEYINPUT105), .B(n353), .ZN(n368) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n355) );
  XNOR2_X1 U413 ( .A(KEYINPUT22), .B(KEYINPUT91), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(n356), .B(KEYINPUT24), .Z(n358) );
  XOR2_X1 U416 ( .A(G50GAT), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(n404), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n363) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(G78GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n359), .B(G148GAT), .ZN(n453) );
  XOR2_X1 U421 ( .A(n453), .B(KEYINPUT87), .Z(n361) );
  NAND2_X1 U422 ( .A1(G228GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U424 ( .A(n363), .B(n362), .Z(n367) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n485) );
  NAND2_X1 U427 ( .A1(n368), .A2(n485), .ZN(n369) );
  XNOR2_X1 U428 ( .A(KEYINPUT25), .B(n369), .ZN(n373) );
  NOR2_X1 U429 ( .A1(n485), .A2(n539), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n370), .B(KEYINPUT26), .ZN(n575) );
  XNOR2_X1 U431 ( .A(KEYINPUT27), .B(n530), .ZN(n376) );
  NAND2_X1 U432 ( .A1(n575), .A2(n376), .ZN(n371) );
  XOR2_X1 U433 ( .A(KEYINPUT104), .B(n371), .Z(n372) );
  NOR2_X1 U434 ( .A1(n373), .A2(n372), .ZN(n374) );
  NOR2_X1 U435 ( .A1(n528), .A2(n374), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n485), .B(KEYINPUT67), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n375), .B(KEYINPUT28), .ZN(n541) );
  NAND2_X1 U438 ( .A1(n376), .A2(n528), .ZN(n377) );
  XOR2_X1 U439 ( .A(n377), .B(KEYINPUT103), .Z(n537) );
  NOR2_X1 U440 ( .A1(n541), .A2(n378), .ZN(n379) );
  NOR2_X1 U441 ( .A1(n380), .A2(n379), .ZN(n497) );
  INV_X1 U442 ( .A(n497), .ZN(n422) );
  XOR2_X1 U443 ( .A(G57GAT), .B(KEYINPUT13), .Z(n450) );
  XOR2_X1 U444 ( .A(n381), .B(n450), .Z(n383) );
  XNOR2_X1 U445 ( .A(G211GAT), .B(G78GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U447 ( .A(G64GAT), .B(KEYINPUT83), .Z(n385) );
  NAND2_X1 U448 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U450 ( .A(n387), .B(n386), .Z(n390) );
  XOR2_X1 U451 ( .A(G22GAT), .B(G1GAT), .Z(n435) );
  XNOR2_X1 U452 ( .A(n435), .B(n388), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n398) );
  XOR2_X1 U454 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n392) );
  XNOR2_X1 U455 ( .A(G71GAT), .B(G155GAT), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U457 ( .A(KEYINPUT82), .B(KEYINPUT15), .Z(n394) );
  XNOR2_X1 U458 ( .A(KEYINPUT84), .B(KEYINPUT81), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U460 ( .A(n396), .B(n395), .Z(n397) );
  XOR2_X1 U461 ( .A(n398), .B(n397), .Z(n584) );
  INV_X1 U462 ( .A(n584), .ZN(n494) );
  XOR2_X1 U463 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n400) );
  XNOR2_X1 U464 ( .A(G43GAT), .B(G29GAT), .ZN(n399) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U466 ( .A(KEYINPUT7), .B(n401), .Z(n441) );
  INV_X1 U467 ( .A(n441), .ZN(n408) );
  XOR2_X1 U468 ( .A(G92GAT), .B(KEYINPUT73), .Z(n403) );
  XNOR2_X1 U469 ( .A(G99GAT), .B(G85GAT), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n403), .B(n402), .ZN(n447) );
  XOR2_X1 U471 ( .A(n447), .B(n404), .Z(n406) );
  NAND2_X1 U472 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U473 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U474 ( .A(n408), .B(n407), .Z(n420) );
  XOR2_X1 U475 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n410) );
  XNOR2_X1 U476 ( .A(G106GAT), .B(KEYINPUT66), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U478 ( .A(n411), .B(KEYINPUT9), .Z(n414) );
  XNOR2_X1 U479 ( .A(G218GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U481 ( .A(n415), .B(KEYINPUT78), .Z(n418) );
  XNOR2_X1 U482 ( .A(n416), .B(KEYINPUT77), .ZN(n417) );
  XNOR2_X1 U483 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U484 ( .A(n420), .B(n419), .Z(n470) );
  XOR2_X1 U485 ( .A(KEYINPUT36), .B(KEYINPUT108), .Z(n421) );
  XOR2_X1 U486 ( .A(n470), .B(n421), .Z(n588) );
  NAND2_X1 U487 ( .A1(n422), .A2(n293), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n423), .B(KEYINPUT37), .ZN(n527) );
  XOR2_X1 U489 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n425) );
  XNOR2_X1 U490 ( .A(KEYINPUT30), .B(KEYINPUT71), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n439) );
  XOR2_X1 U492 ( .A(G141GAT), .B(G197GAT), .Z(n427) );
  XNOR2_X1 U493 ( .A(G36GAT), .B(G50GAT), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U495 ( .A(G8GAT), .B(G113GAT), .Z(n429) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(G15GAT), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U498 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U499 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n433) );
  NAND2_X1 U500 ( .A1(G229GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U501 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U502 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U504 ( .A(n439), .B(n438), .Z(n440) );
  XOR2_X1 U505 ( .A(n441), .B(n440), .Z(n577) );
  XOR2_X1 U506 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n443) );
  XNOR2_X1 U507 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n442) );
  XNOR2_X1 U508 ( .A(n443), .B(n442), .ZN(n458) );
  AND2_X1 U509 ( .A1(G230GAT), .A2(G233GAT), .ZN(n445) );
  INV_X1 U510 ( .A(KEYINPUT33), .ZN(n444) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(n468) );
  INV_X1 U515 ( .A(n468), .ZN(n459) );
  INV_X1 U516 ( .A(n459), .ZN(n581) );
  NOR2_X1 U517 ( .A1(n577), .A2(n581), .ZN(n498) );
  NAND2_X1 U518 ( .A1(n527), .A2(n498), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n539), .A2(n512), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n462) );
  XNOR2_X1 U521 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n461) );
  INV_X1 U522 ( .A(KEYINPUT54), .ZN(n482) );
  NOR2_X1 U523 ( .A1(n588), .A2(n494), .ZN(n465) );
  XOR2_X1 U524 ( .A(KEYINPUT45), .B(n465), .Z(n466) );
  NOR2_X1 U525 ( .A1(n581), .A2(n466), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n467), .A2(n577), .ZN(n476) );
  XOR2_X1 U527 ( .A(KEYINPUT41), .B(n468), .Z(n568) );
  INV_X1 U528 ( .A(n577), .ZN(n566) );
  AND2_X1 U529 ( .A1(n568), .A2(n566), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT46), .ZN(n472) );
  INV_X1 U531 ( .A(n470), .ZN(n563) );
  OR2_X1 U532 ( .A1(n584), .A2(n563), .ZN(n471) );
  OR2_X1 U533 ( .A1(n472), .A2(n471), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT47), .B(KEYINPUT116), .Z(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n479) );
  INV_X1 U537 ( .A(KEYINPUT48), .ZN(n477) );
  NOR2_X1 U538 ( .A1(n538), .A2(n480), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  NOR2_X1 U540 ( .A1(n528), .A2(n483), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT65), .B(n484), .Z(n576) );
  NAND2_X1 U542 ( .A1(n576), .A2(n485), .ZN(n487) );
  XOR2_X1 U543 ( .A(KEYINPUT124), .B(KEYINPUT55), .Z(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(n489) );
  NOR2_X2 U545 ( .A1(n489), .A2(n488), .ZN(n572) );
  AND2_X1 U546 ( .A1(n572), .A2(n563), .ZN(n493) );
  XNOR2_X1 U547 ( .A(KEYINPUT126), .B(KEYINPUT58), .ZN(n491) );
  INV_X1 U548 ( .A(G190GAT), .ZN(n490) );
  XOR2_X1 U549 ( .A(KEYINPUT34), .B(KEYINPUT106), .Z(n500) );
  NOR2_X1 U550 ( .A1(n563), .A2(n494), .ZN(n495) );
  XOR2_X1 U551 ( .A(KEYINPUT16), .B(n495), .Z(n496) );
  NOR2_X1 U552 ( .A1(n497), .A2(n496), .ZN(n516) );
  AND2_X1 U553 ( .A1(n498), .A2(n516), .ZN(n505) );
  NAND2_X1 U554 ( .A1(n505), .A2(n528), .ZN(n499) );
  XNOR2_X1 U555 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U556 ( .A(G1GAT), .B(n501), .Z(G1324GAT) );
  NAND2_X1 U557 ( .A1(n505), .A2(n530), .ZN(n502) );
  XNOR2_X1 U558 ( .A(n502), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .Z(n504) );
  NAND2_X1 U560 ( .A1(n505), .A2(n539), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n504), .B(n503), .ZN(G1326GAT) );
  NAND2_X1 U562 ( .A1(n505), .A2(n541), .ZN(n506) );
  XNOR2_X1 U563 ( .A(n506), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U564 ( .A1(n512), .A2(n528), .ZN(n510) );
  XOR2_X1 U565 ( .A(KEYINPUT109), .B(KEYINPUT39), .Z(n508) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT107), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U568 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  NAND2_X1 U569 ( .A1(n530), .A2(n512), .ZN(n511) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n511), .ZN(G1329GAT) );
  NAND2_X1 U571 ( .A1(n512), .A2(n541), .ZN(n513) );
  XNOR2_X1 U572 ( .A(n513), .B(KEYINPUT112), .ZN(n514) );
  XNOR2_X1 U573 ( .A(G50GAT), .B(n514), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n518) );
  INV_X1 U575 ( .A(n568), .ZN(n515) );
  NOR2_X1 U576 ( .A1(n515), .A2(n566), .ZN(n526) );
  AND2_X1 U577 ( .A1(n526), .A2(n516), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n523), .A2(n528), .ZN(n517) );
  XNOR2_X1 U579 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n523), .A2(n530), .ZN(n520) );
  XNOR2_X1 U582 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n523), .A2(n539), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n521), .B(KEYINPUT114), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G71GAT), .B(n522), .ZN(G1334GAT) );
  XOR2_X1 U586 ( .A(G78GAT), .B(KEYINPUT43), .Z(n525) );
  NAND2_X1 U587 ( .A1(n523), .A2(n541), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1335GAT) );
  AND2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n528), .A2(n534), .ZN(n529) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n529), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n534), .A2(n530), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT115), .Z(n533) );
  NAND2_X1 U595 ( .A1(n534), .A2(n539), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n534), .A2(n541), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT44), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  XOR2_X1 U600 ( .A(G113GAT), .B(KEYINPUT117), .Z(n543) );
  NOR2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n553) );
  NAND2_X1 U602 ( .A1(n539), .A2(n553), .ZN(n540) );
  NOR2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n549), .A2(n566), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n545) );
  NAND2_X1 U607 ( .A1(n549), .A2(n568), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n546), .ZN(G1341GAT) );
  NAND2_X1 U610 ( .A1(n549), .A2(n584), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U614 ( .A1(n549), .A2(n563), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n575), .ZN(n554) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(n554), .Z(n564) );
  NAND2_X1 U619 ( .A1(n564), .A2(n566), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT121), .B(n558), .Z(n560) );
  NAND2_X1 U625 ( .A1(n564), .A2(n568), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  XOR2_X1 U627 ( .A(G155GAT), .B(KEYINPUT123), .Z(n562) );
  NAND2_X1 U628 ( .A1(n584), .A2(n564), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n572), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n570) );
  NAND2_X1 U635 ( .A1(n572), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(n571), .ZN(G1349GAT) );
  XOR2_X1 U638 ( .A(G183GAT), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U639 ( .A1(n572), .A2(n584), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n587) );
  NOR2_X1 U642 ( .A1(n577), .A2(n587), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  INV_X1 U647 ( .A(n587), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

