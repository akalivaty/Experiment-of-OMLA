//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1349, new_n1350, new_n1351;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n204), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G238), .ZN(new_n215));
  AND2_X1   g0015(.A1(new_n215), .A2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G116), .A2(G270), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n209), .B(new_n214), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G107), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  NAND3_X1  g0040(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(new_n212), .ZN(new_n242));
  INV_X1    g0042(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(KEYINPUT67), .A2(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT8), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n246), .A2(G20), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  INV_X1    g0050(.A(G68), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n252), .A2(G20), .B1(G150), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n243), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(new_n249), .B2(new_n257), .ZN(new_n258));
  AOI211_X1 g0058(.A(new_n242), .B(new_n257), .C1(new_n203), .C2(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G50), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT9), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n267), .A3(G274), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n265), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G226), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n268), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT66), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n246), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(G222), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G223), .A3(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n284), .B(new_n285), .C1(new_n286), .C2(new_n282), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n273), .B1(new_n287), .B2(new_n269), .ZN(new_n288));
  INV_X1    g0088(.A(G200), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(G190), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n262), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n262), .A2(new_n294), .A3(new_n290), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n253), .A2(G50), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n204), .A2(G33), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n297), .B1(new_n204), .B2(G68), .C1(new_n286), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT11), .B1(new_n299), .B2(new_n242), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G68), .B2(new_n259), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n257), .A2(new_n251), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT12), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n299), .A2(KEYINPUT11), .A3(new_n242), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n270), .A2(G238), .ZN(new_n307));
  INV_X1    g0107(.A(G274), .ZN(new_n308));
  AND2_X1   g0108(.A1(G1), .A2(G13), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n266), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(KEYINPUT70), .A3(new_n265), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT70), .B1(new_n310), .B2(new_n265), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n307), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  MUX2_X1   g0114(.A(G226), .B(G232), .S(G1698), .Z(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT66), .B1(new_n274), .B2(new_n275), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n279), .A2(new_n277), .A3(new_n280), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n267), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT13), .B1(new_n314), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n319), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n269), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT70), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n268), .A2(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(new_n311), .B1(G238), .B2(new_n270), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT13), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n323), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n321), .A2(new_n328), .A3(G190), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n306), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n289), .B1(new_n321), .B2(new_n328), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n314), .A2(new_n320), .A3(KEYINPUT13), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n327), .B1(new_n323), .B2(new_n326), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G169), .ZN(new_n336));
  OAI211_X1 g0136(.A(KEYINPUT71), .B(KEYINPUT14), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT71), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n336), .B1(new_n321), .B2(new_n328), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(G179), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT72), .B(KEYINPUT14), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n337), .A2(new_n341), .A3(new_n342), .A4(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n332), .B1(new_n345), .B2(new_n305), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT68), .B(G179), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n288), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n348), .B(new_n261), .C1(G169), .C2(new_n288), .ZN(new_n349));
  INV_X1    g0149(.A(G244), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n268), .B1(new_n271), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G232), .A2(G1698), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n215), .A2(new_n283), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n282), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n316), .A2(new_n317), .ZN(new_n355));
  INV_X1    g0155(.A(G107), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n267), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n351), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n336), .ZN(new_n360));
  XOR2_X1   g0160(.A(KEYINPUT15), .B(G87), .Z(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n247), .B1(G20), .B2(G77), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT8), .B(G58), .Z(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n253), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n243), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n256), .A2(G77), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n259), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n367), .B1(new_n286), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n358), .A2(new_n347), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n360), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT69), .ZN(new_n372));
  INV_X1    g0172(.A(G190), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n359), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n367), .B1(new_n286), .B2(new_n368), .C1(new_n358), .C2(new_n289), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n359), .B2(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n296), .A2(new_n346), .A3(new_n349), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n245), .A2(new_n256), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n259), .B2(new_n245), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  XNOR2_X1  g0182(.A(G58), .B(G68), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G20), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n253), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n279), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n280), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n204), .B1(new_n276), .B2(new_n281), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n387), .B1(new_n392), .B2(new_n251), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n279), .A2(new_n204), .A3(new_n280), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n391), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n388), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n386), .B1(new_n398), .B2(G68), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n243), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n382), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n272), .A2(G1698), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(G223), .B2(G1698), .C1(new_n274), .C2(new_n275), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n267), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n267), .A2(G232), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n268), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n289), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n405), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n268), .A2(new_n407), .A3(KEYINPUT73), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT73), .B1(new_n268), .B2(new_n407), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n409), .B1(new_n413), .B2(G190), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(G20), .B1(new_n316), .B2(new_n317), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n388), .B1(new_n416), .B2(KEYINPUT7), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n386), .B1(new_n417), .B2(G68), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n400), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(new_n381), .A3(new_n414), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n415), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n410), .B(new_n347), .C1(new_n411), .C2(new_n412), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n336), .B1(new_n405), .B2(new_n408), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI211_X1 g0227(.A(new_n424), .B(new_n427), .C1(new_n419), .C2(new_n381), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n427), .B1(new_n419), .B2(new_n381), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT74), .B1(new_n429), .B2(KEYINPUT18), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT74), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(new_n424), .C1(new_n401), .C2(new_n427), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n379), .A2(new_n423), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n283), .A2(G244), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n279), .B2(new_n280), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT76), .B1(new_n436), .B2(KEYINPUT4), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G283), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT76), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT4), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n274), .A2(new_n275), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n439), .B(new_n440), .C1(new_n441), .C2(new_n435), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n316), .A2(new_n317), .A3(G250), .A4(G1698), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n440), .A2(new_n350), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n316), .A2(new_n317), .A3(new_n283), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n269), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n264), .A2(G1), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT5), .B(G41), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n310), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n267), .ZN(new_n455));
  INV_X1    g0255(.A(G257), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G200), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n203), .A2(G33), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n256), .A2(new_n461), .A3(new_n212), .A4(new_n241), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G97), .ZN(new_n463));
  INV_X1    g0263(.A(G97), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n256), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(KEYINPUT75), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT75), .B1(new_n463), .B2(new_n465), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n253), .A2(G77), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT6), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n471), .A2(new_n464), .A3(G107), .ZN(new_n472));
  XNOR2_X1  g0272(.A(G97), .B(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n470), .B1(new_n474), .B2(new_n204), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n392), .B2(new_n356), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n469), .B1(new_n477), .B2(new_n242), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n448), .A2(G190), .A3(new_n458), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n460), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n468), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n466), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n475), .B1(new_n417), .B2(G107), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(new_n243), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n448), .A2(new_n347), .A3(new_n458), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n440), .B1(new_n441), .B2(new_n435), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n486), .A2(KEYINPUT76), .B1(G33), .B2(G283), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n487), .A2(new_n442), .A3(new_n444), .A4(new_n446), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n457), .B1(new_n488), .B2(new_n269), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n484), .B(new_n485), .C1(new_n489), .C2(G169), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n361), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n257), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n492), .A2(new_n462), .ZN(new_n494));
  OR2_X1    g0294(.A1(KEYINPUT78), .A2(G87), .ZN(new_n495));
  NOR2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NAND2_X1  g0296(.A1(KEYINPUT78), .A2(G87), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n319), .B2(new_n204), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n298), .B2(new_n464), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n279), .A2(new_n280), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n204), .A4(G68), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n504), .A2(new_n204), .A3(G68), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT79), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n503), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n493), .B(new_n494), .C1(new_n509), .C2(new_n243), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT80), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n508), .A2(new_n506), .ZN(new_n513));
  INV_X1    g0313(.A(new_n503), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n242), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(KEYINPUT80), .A3(new_n493), .A4(new_n494), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(G238), .A2(G1698), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n350), .B2(G1698), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n504), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n246), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n269), .ZN(new_n526));
  INV_X1    g0326(.A(new_n347), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n449), .A2(new_n308), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n528), .B(new_n267), .C1(G250), .C2(new_n449), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT77), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n523), .B1(new_n520), .B2(new_n504), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n532), .B2(new_n267), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(G169), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n531), .B1(new_n530), .B2(new_n534), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(G264), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n455), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G294), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n246), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n456), .B1(new_n279), .B2(new_n280), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n542), .B2(G1698), .ZN(new_n543));
  INV_X1    g0343(.A(G250), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G1698), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT85), .B1(new_n504), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n545), .B(KEYINPUT85), .C1(new_n275), .C2(new_n274), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n539), .B1(new_n549), .B2(new_n269), .ZN(new_n550));
  AOI21_X1  g0350(.A(G169), .B1(new_n550), .B2(new_n451), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n545), .B1(new_n274), .B2(new_n275), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT85), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n547), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n267), .B1(new_n555), .B2(new_n543), .ZN(new_n556));
  INV_X1    g0356(.A(new_n451), .ZN(new_n557));
  NOR4_X1   g0357(.A1(new_n556), .A2(G179), .A3(new_n557), .A4(new_n539), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n204), .B(G87), .C1(new_n274), .C2(new_n275), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT22), .ZN(new_n561));
  INV_X1    g0361(.A(G87), .ZN(new_n562));
  OR3_X1    g0362(.A1(new_n562), .A2(KEYINPUT22), .A3(G20), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n561), .B1(new_n355), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT24), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n204), .B2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n356), .A2(KEYINPUT23), .A3(G20), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n567), .A2(new_n568), .B1(new_n523), .B2(new_n204), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n564), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n565), .B1(new_n564), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n242), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT25), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n256), .B2(G107), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n256), .A2(new_n573), .A3(G107), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n575), .A2(new_n576), .B1(new_n356), .B2(new_n462), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n518), .A2(new_n537), .B1(new_n559), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n533), .A2(G200), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n373), .B2(new_n533), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n243), .B1(new_n513), .B2(new_n514), .ZN(new_n583));
  INV_X1    g0383(.A(new_n493), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n462), .A2(new_n562), .ZN(new_n585));
  NOR4_X1   g0385(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NOR4_X1   g0386(.A1(new_n556), .A2(new_n373), .A3(new_n557), .A4(new_n539), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n550), .A2(new_n451), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n587), .B1(G200), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n572), .A2(new_n578), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n491), .A2(new_n580), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n454), .A2(G270), .A3(new_n267), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT81), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n593), .A2(new_n594), .A3(new_n451), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n593), .B2(new_n451), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n538), .A2(new_n283), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n355), .A2(G303), .B1(new_n504), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(G257), .B(new_n283), .C1(new_n274), .C2(new_n275), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n504), .A2(KEYINPUT82), .A3(G257), .A4(new_n283), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n267), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G190), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n355), .A2(G303), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n504), .A2(new_n598), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n269), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n593), .A2(new_n451), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n593), .A2(new_n451), .A3(new_n594), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G200), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n241), .A2(new_n212), .B1(G20), .B2(new_n522), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n438), .B(new_n204), .C1(G33), .C2(new_n464), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n618), .A2(KEYINPUT20), .A3(new_n619), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n257), .A2(new_n522), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n462), .B2(new_n522), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n607), .A2(new_n617), .A3(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n618), .A2(KEYINPUT20), .A3(new_n619), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT20), .B1(new_n618), .B2(new_n619), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(G169), .B1(new_n633), .B2(new_n626), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n634), .B1(new_n611), .B2(new_n615), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n628), .A2(G179), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n635), .A2(KEYINPUT21), .B1(new_n606), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n336), .B1(new_n624), .B2(new_n627), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n597), .B2(new_n605), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT83), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n630), .B(new_n638), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(KEYINPUT84), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n640), .A2(new_n642), .B1(new_n616), .B2(new_n636), .ZN(new_n648));
  OAI21_X1  g0448(.A(KEYINPUT83), .B1(new_n635), .B2(KEYINPUT21), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n648), .B1(new_n649), .B2(new_n643), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n630), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n592), .B1(new_n647), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n434), .A2(new_n653), .ZN(G372));
  INV_X1    g0454(.A(KEYINPUT86), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n490), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n530), .A2(new_n534), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n518), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n586), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n459), .A2(new_n336), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n660), .A2(KEYINPUT86), .A3(new_n485), .A4(new_n484), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n656), .A2(new_n658), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n518), .A2(new_n537), .ZN(new_n665));
  INV_X1    g0465(.A(new_n490), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n659), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n663), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n588), .A2(G200), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n550), .A2(G190), .A3(new_n451), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n572), .A3(new_n578), .A4(new_n670), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n659), .A2(new_n671), .A3(new_n480), .A4(new_n490), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n559), .A2(new_n579), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n674), .B(new_n638), .C1(new_n644), .C2(new_n645), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n673), .A2(new_n675), .B1(new_n518), .B2(new_n657), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n434), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n349), .ZN(new_n679));
  INV_X1    g0479(.A(new_n332), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n680), .A2(new_n371), .B1(new_n345), .B2(new_n305), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n417), .A2(G68), .ZN(new_n682));
  AOI21_X1  g0482(.A(KEYINPUT16), .B1(new_n682), .B2(new_n387), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n399), .A2(KEYINPUT16), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n242), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n381), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n427), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT18), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n681), .A2(new_n423), .B1(new_n428), .B2(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n679), .B1(new_n689), .B2(new_n296), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n678), .A2(new_n690), .ZN(G369));
  NAND3_X1  g0491(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(KEYINPUT87), .B(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n647), .A2(new_n652), .B1(new_n628), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n697), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n650), .A2(new_n629), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n579), .A2(new_n697), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n671), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n674), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n699), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n701), .A2(G330), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n638), .B1(new_n644), .B2(new_n645), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n703), .A2(new_n710), .A3(new_n674), .A4(new_n699), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n709), .A2(new_n706), .A3(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n207), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n498), .A2(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n210), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT28), .ZN(new_n719));
  AOI211_X1 g0519(.A(KEYINPUT29), .B(new_n697), .C1(new_n668), .C2(new_n676), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n662), .A2(KEYINPUT26), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n675), .A2(new_n491), .A3(new_n591), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n665), .A2(new_n666), .A3(new_n663), .A4(new_n659), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n722), .A2(new_n723), .A3(new_n658), .A4(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n721), .B1(new_n725), .B2(new_n699), .ZN(new_n726));
  INV_X1    g0526(.A(G330), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n665), .A2(new_n674), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n672), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n646), .A2(KEYINPUT84), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n651), .B1(new_n650), .B2(new_n630), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n729), .B(new_n699), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  INV_X1    g0533(.A(G179), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n533), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n611), .A2(new_n550), .A3(new_n615), .A4(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n733), .B1(new_n736), .B2(new_n459), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n527), .B1(new_n526), .B2(new_n529), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n616), .A2(new_n459), .A3(new_n588), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT88), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n737), .A2(KEYINPUT88), .A3(new_n739), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n550), .A2(new_n735), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n489), .A3(new_n606), .A4(KEYINPUT30), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n742), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT31), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n699), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n737), .A2(new_n745), .A3(new_n739), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n697), .ZN(new_n750));
  AOI22_X1  g0550(.A1(new_n746), .A2(new_n748), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n727), .B1(new_n732), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n720), .A2(new_n726), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n719), .B1(new_n753), .B2(G1), .ZN(G364));
  NAND2_X1  g0554(.A1(new_n701), .A2(G330), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n204), .A2(G13), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n203), .B1(new_n756), .B2(G45), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n714), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n698), .A2(new_n700), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n727), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n755), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT89), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n212), .B1(G20), .B2(new_n336), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n204), .A2(G190), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n772), .A2(new_n734), .A3(G200), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT91), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G107), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n734), .A2(G20), .A3(G190), .A4(G200), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n495), .B2(new_n497), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n355), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT92), .Z(new_n784));
  NOR2_X1   g0584(.A1(new_n347), .A2(new_n204), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n373), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G190), .A2(G200), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G58), .A2(new_n788), .B1(new_n791), .B2(G77), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n249), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT32), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n734), .A2(new_n289), .A3(KEYINPUT90), .ZN(new_n796));
  AOI21_X1  g0596(.A(KEYINPUT90), .B1(new_n734), .B2(new_n289), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n772), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n798), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(KEYINPUT32), .A3(G159), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n794), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n784), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n796), .A2(new_n797), .ZN(new_n805));
  OAI21_X1  g0605(.A(G20), .B1(new_n805), .B2(new_n373), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G97), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n785), .A2(new_n373), .A3(G200), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n251), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n778), .A2(G283), .B1(new_n801), .B2(G329), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n812), .B2(new_n790), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  INV_X1    g0614(.A(G322), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n355), .B1(new_n814), .B2(new_n780), .C1(new_n787), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n793), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(G326), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n806), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT94), .B(KEYINPUT33), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(G317), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n818), .B1(new_n540), .B2(new_n819), .C1(new_n808), .C2(new_n821), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n804), .A2(new_n810), .B1(new_n813), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n771), .B1(new_n823), .B2(KEYINPUT95), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(KEYINPUT95), .B2(new_n823), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n713), .A2(new_n504), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(new_n264), .B2(new_n211), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n236), .B2(new_n264), .ZN(new_n829));
  INV_X1    g0629(.A(G355), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n282), .A2(new_n207), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n829), .B1(G116), .B2(new_n207), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n768), .A2(new_n770), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n760), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n769), .A2(new_n825), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n765), .A2(new_n835), .ZN(G396));
  NAND2_X1  g0636(.A1(new_n369), .A2(new_n697), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n371), .A2(KEYINPUT97), .A3(new_n697), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT97), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n360), .A2(new_n369), .A3(new_n370), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n699), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n378), .A2(new_n837), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n677), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n697), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n378), .A2(new_n837), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n838), .A2(new_n841), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g0647(.A1(KEYINPUT26), .A2(new_n665), .A3(new_n666), .A4(new_n659), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(new_n663), .B2(new_n662), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n723), .A2(new_n658), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n699), .B(new_n847), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n752), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n759), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n853), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n771), .A2(new_n767), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n759), .B1(G77), .B2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(G143), .A2(new_n788), .B1(new_n791), .B2(G159), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  INV_X1    g0659(.A(G150), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n859), .B2(new_n793), .C1(new_n860), .C2(new_n808), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT34), .Z(new_n862));
  OAI21_X1  g0662(.A(new_n504), .B1(new_n249), .B2(new_n780), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(new_n801), .B2(G132), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n864), .B1(new_n777), .B2(new_n251), .C1(new_n819), .C2(new_n250), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT96), .Z(new_n866));
  NOR2_X1   g0666(.A1(new_n777), .A2(new_n562), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n868), .B1(new_n522), .B2(new_n790), .C1(new_n812), .C2(new_n798), .ZN(new_n869));
  INV_X1    g0669(.A(new_n808), .ZN(new_n870));
  AOI22_X1  g0670(.A1(G283), .A2(new_n870), .B1(new_n817), .B2(G303), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n355), .B1(new_n356), .B2(new_n780), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n788), .B2(G294), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n807), .A3(new_n873), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n862), .A2(new_n866), .B1(new_n869), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n857), .B1(new_n875), .B2(new_n770), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n847), .B2(new_n767), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n855), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(G384));
  NAND2_X1  g0679(.A1(new_n473), .A2(new_n471), .ZN(new_n880));
  INV_X1    g0680(.A(new_n472), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n883), .A2(G116), .A3(new_n213), .A4(new_n884), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT36), .Z(new_n886));
  NOR2_X1   g0686(.A1(new_n251), .A2(G50), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT98), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n211), .B(G77), .C1(new_n250), .C2(new_n251), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n203), .B(G13), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n399), .A2(KEYINPUT16), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n381), .B1(new_n685), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n695), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n433), .B2(new_n423), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n686), .A2(new_n687), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n686), .A2(new_n894), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT37), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n420), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n893), .B1(new_n687), .B2(new_n894), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n420), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n901), .B1(new_n903), .B2(new_n900), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n897), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n750), .A2(new_n747), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n653), .B2(new_n699), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n305), .B(new_n697), .C1(new_n345), .C2(new_n332), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n306), .A2(new_n699), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n916), .B(new_n332), .C1(new_n345), .C2(new_n305), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n847), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n909), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n910), .A2(new_n911), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n732), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n916), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n346), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n842), .B1(new_n925), .B2(new_n914), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(new_n899), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n428), .A2(new_n688), .ZN(new_n929));
  OAI211_X1 g0729(.A(KEYINPUT99), .B(new_n928), .C1(new_n929), .C2(new_n423), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n898), .A2(new_n899), .A3(new_n420), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(KEYINPUT37), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n901), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n422), .B(new_n415), .C1(new_n428), .C2(new_n688), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT99), .B1(new_n935), .B2(new_n928), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n906), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n927), .B1(new_n908), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n921), .B1(new_n938), .B2(new_n920), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT100), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n434), .A2(new_n923), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n942), .A2(new_n943), .A3(new_n727), .ZN(new_n944));
  AND3_X1   g0744(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT38), .B1(new_n897), .B2(new_n904), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT39), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n937), .A2(new_n908), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT39), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n345), .A2(new_n305), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(new_n697), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n948), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n915), .A2(new_n917), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n371), .A2(new_n699), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n955), .B1(new_n851), .B2(new_n956), .ZN(new_n957));
  AOI22_X1  g0757(.A1(new_n957), .A2(new_n909), .B1(new_n929), .B2(new_n695), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n434), .B1(new_n720), .B2(new_n726), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n690), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT101), .B1(new_n944), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n944), .A2(new_n962), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n203), .C2(new_n756), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n944), .A2(KEYINPUT101), .A3(new_n962), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n891), .B1(new_n965), .B2(new_n966), .ZN(G367));
  NAND2_X1  g0767(.A1(new_n826), .A2(new_n232), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n968), .B(new_n833), .C1(new_n207), .C2(new_n492), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n793), .A2(new_n812), .B1(new_n787), .B2(new_n814), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT104), .Z(new_n971));
  INV_X1    g0771(.A(G283), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n441), .B1(new_n790), .B2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n777), .A2(new_n464), .B1(new_n974), .B2(new_n798), .ZN(new_n975));
  OAI21_X1  g0775(.A(KEYINPUT105), .B1(new_n780), .B2(new_n522), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT46), .Z(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n540), .B2(new_n808), .C1(new_n819), .C2(new_n356), .ZN(new_n978));
  NOR4_X1   g0778(.A1(new_n971), .A2(new_n973), .A3(new_n975), .A4(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT106), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n817), .A2(G143), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n860), .B2(new_n787), .C1(new_n251), .C2(new_n819), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT107), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT107), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n282), .B1(new_n790), .B2(new_n249), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n777), .A2(new_n286), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G159), .C2(new_n870), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n798), .A2(new_n859), .B1(new_n250), .B2(new_n780), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT108), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n984), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n980), .B1(new_n983), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT47), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n991), .B(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n759), .B(new_n969), .C1(new_n993), .C2(new_n771), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT109), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n516), .A2(new_n493), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n697), .B1(new_n997), .B2(new_n585), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n658), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n658), .A2(new_n659), .A3(new_n998), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n768), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n994), .A2(new_n995), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n996), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n753), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n711), .A2(new_n706), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT102), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n666), .A2(new_n1009), .A3(new_n697), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT102), .B1(new_n490), .B2(new_n699), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n484), .A2(new_n697), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1010), .A2(new_n1011), .B1(new_n491), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n709), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n709), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n707), .B1(new_n650), .B2(new_n697), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n755), .A2(new_n711), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n711), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(G330), .A3(new_n701), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1007), .B1(new_n1022), .B2(new_n1027), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n714), .B(KEYINPUT41), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n757), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n1013), .A2(new_n711), .A3(KEYINPUT42), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT42), .B1(new_n1013), .B2(new_n711), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT43), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1013), .A2(new_n674), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n699), .B1(new_n1036), .B2(new_n666), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1002), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1002), .A2(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1037), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1039), .B(new_n1040), .C1(new_n1041), .C2(new_n1033), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n709), .B2(new_n1013), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n709), .A2(new_n1013), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1038), .A2(new_n1042), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT103), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1038), .A2(new_n1042), .A3(new_n1045), .A4(KEYINPUT103), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1044), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1006), .B1(new_n1030), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(G387));
  NAND2_X1  g0853(.A1(new_n1027), .A2(new_n753), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n714), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT111), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1007), .A2(new_n1026), .A3(new_n1024), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(KEYINPUT111), .A3(new_n714), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n826), .B1(new_n229), .B2(new_n264), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n716), .B2(new_n831), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n363), .A2(new_n249), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1064));
  XNOR2_X1  g0864(.A(new_n1063), .B(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n716), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1062), .A2(new_n1067), .B1(new_n356), .B2(new_n713), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n833), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n759), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G317), .A2(new_n788), .B1(new_n791), .B2(G303), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n812), .B2(new_n808), .C1(new_n815), .C2(new_n793), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT48), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n780), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n806), .A2(G283), .B1(G294), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT49), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n777), .A2(new_n522), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n504), .B(new_n1082), .C1(G326), .C2(new_n801), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n780), .A2(new_n286), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n441), .B(new_n1085), .C1(new_n778), .C2(G97), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n787), .A2(new_n249), .B1(new_n860), .B2(new_n798), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G68), .B2(new_n791), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n806), .A2(new_n361), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G159), .A2(new_n817), .B1(new_n870), .B2(new_n245), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1086), .A2(new_n1088), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n771), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1070), .B(new_n1092), .C1(new_n707), .C2(new_n768), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1027), .B2(new_n758), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1060), .A2(new_n1094), .ZN(G393));
  OAI221_X1 g0895(.A(new_n833), .B1(new_n464), .B2(new_n207), .C1(new_n827), .C2(new_n239), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n819), .A2(new_n286), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n791), .A2(new_n363), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n801), .A2(G143), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n441), .B1(new_n1076), .B2(G68), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n868), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1097), .B(new_n1101), .C1(G50), .C2(new_n870), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n793), .A2(new_n860), .B1(new_n787), .B2(new_n799), .ZN(new_n1103));
  XOR2_X1   g0903(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1104));
  XNOR2_X1  g0904(.A(new_n1103), .B(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n793), .A2(new_n974), .B1(new_n787), .B2(new_n812), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n870), .A2(G303), .B1(G116), .B2(new_n806), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n282), .B1(G283), .B2(new_n1076), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n791), .A2(G294), .B1(G322), .B2(new_n801), .ZN(new_n1110));
  AND4_X1   g0910(.A1(new_n779), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1102), .A2(new_n1105), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n759), .B(new_n1096), .C1(new_n1112), .C2(new_n771), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1013), .B2(new_n768), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n1022), .B2(new_n758), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1021), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1116), .A2(new_n753), .A3(new_n1027), .A4(new_n1019), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n714), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1116), .A2(new_n1019), .B1(new_n753), .B2(new_n1027), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1115), .B1(new_n1118), .B2(new_n1119), .ZN(G390));
  NOR2_X1   g0920(.A1(new_n913), .A2(new_n727), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n434), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n960), .A2(new_n1122), .A3(new_n690), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n851), .A2(new_n956), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n923), .A2(G330), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n918), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n955), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n752), .B2(new_n847), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1124), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n955), .B1(new_n1125), .B2(new_n842), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n752), .A2(new_n1127), .A3(new_n847), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n725), .A2(new_n699), .A3(new_n847), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1130), .A2(new_n956), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1123), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1126), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT113), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n953), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n951), .A2(new_n948), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1132), .A2(new_n956), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1127), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n953), .B1(new_n937), .B2(new_n908), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1136), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n948), .A2(new_n951), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1131), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT113), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1135), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1148), .A2(new_n1151), .A3(new_n1143), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1134), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(new_n715), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1145), .A2(new_n1152), .A3(new_n1134), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1145), .A2(new_n1152), .A3(new_n758), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n767), .B1(new_n948), .B2(new_n951), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n282), .B1(new_n777), .B2(new_n249), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G125), .B2(new_n801), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT114), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n780), .A2(new_n860), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G132), .A2(new_n788), .B1(new_n791), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n819), .A2(new_n799), .B1(new_n1167), .B2(new_n793), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(G137), .B2(new_n870), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1161), .A2(new_n1163), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n787), .A2(new_n522), .B1(new_n540), .B2(new_n798), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n791), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n355), .B1(new_n562), .B2(new_n780), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n778), .B2(G68), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1097), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G107), .A2(new_n870), .B1(new_n817), .B2(G283), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n771), .B1(new_n1170), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n759), .B1(new_n245), .B2(new_n856), .ZN(new_n1179));
  OR3_X1    g0979(.A1(new_n1158), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1156), .A2(new_n1157), .A3(new_n1180), .ZN(G378));
  NAND2_X1  g0981(.A1(new_n954), .A2(new_n958), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n296), .A2(new_n349), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n261), .A2(new_n894), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT55), .Z(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1183), .A3(new_n1188), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n939), .B2(G330), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n920), .B1(new_n949), .B2(new_n919), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n923), .A2(new_n926), .A3(new_n920), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n947), .A2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G330), .B(new_n1194), .C1(new_n1196), .C2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1182), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1194), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n727), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n959), .A3(new_n1199), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1201), .A2(KEYINPUT119), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1123), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1155), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT119), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1209), .B(new_n1182), .C1(new_n1195), .C2(new_n1200), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT57), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1155), .B2(new_n1207), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1201), .A2(new_n1205), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n715), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1206), .A2(new_n758), .A3(new_n1210), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1202), .A2(new_n766), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n759), .B1(G50), .B2(new_n856), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n788), .A2(G107), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT115), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1221), .A2(new_n1222), .B1(new_n464), .B2(new_n808), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G116), .B2(new_n817), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n777), .A2(new_n250), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n790), .A2(new_n492), .B1(new_n972), .B2(new_n798), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n441), .A2(new_n263), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1085), .A4(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1221), .A2(new_n1222), .B1(G68), .B2(new_n806), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1224), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT58), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(G33), .A2(G41), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(G50), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1230), .A2(new_n1231), .B1(new_n1227), .B2(new_n1233), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n787), .A2(new_n1167), .B1(new_n780), .B2(new_n1164), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT116), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n817), .A2(G125), .B1(new_n791), .B2(G137), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n870), .A2(G132), .B1(G150), .B2(new_n806), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  XOR2_X1   g1039(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1240));
  XNOR2_X1  g1040(.A(new_n1239), .B(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n801), .A2(G124), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1232), .C1(new_n777), .C2(new_n799), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1234), .B1(new_n1231), .B2(new_n1230), .C1(new_n1241), .C2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1220), .B1(new_n1244), .B2(new_n770), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1219), .A2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1218), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1217), .A2(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n1133), .A2(new_n1129), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(new_n1207), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(new_n1029), .A3(new_n1134), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT120), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n759), .B1(G68), .B2(new_n856), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n282), .B(new_n986), .C1(G97), .C2(new_n1076), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n787), .A2(new_n972), .B1(new_n814), .B2(new_n798), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1255), .B1(G107), .B2(new_n791), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G116), .A2(new_n870), .B1(new_n817), .B2(G294), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1089), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT121), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n441), .B(new_n1225), .C1(G159), .C2(new_n1076), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n787), .A2(new_n859), .B1(new_n1167), .B2(new_n798), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G150), .B2(new_n791), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n806), .A2(G50), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(G132), .A2(new_n817), .B1(new_n870), .B2(new_n1165), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1261), .A2(new_n1263), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1260), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1253), .B1(new_n1268), .B2(new_n770), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n1127), .B2(new_n767), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1249), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n757), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1252), .A2(new_n1273), .ZN(G381));
  INV_X1    g1074(.A(G390), .ZN(new_n1275));
  INV_X1    g1075(.A(G396), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1059), .A2(new_n1058), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT111), .B1(new_n1054), .B2(new_n714), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1276), .B(new_n1094), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1052), .A2(new_n878), .A3(new_n1275), .A4(new_n1280), .ZN(new_n1281));
  OR4_X1    g1081(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1281), .ZN(G407));
  AND3_X1   g1082(.A1(new_n1156), .A2(new_n1157), .A3(new_n1180), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n696), .A2(G213), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT122), .Z(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(G407), .B(G213), .C1(G375), .C2(new_n1286), .ZN(G409));
  AOI21_X1  g1087(.A(new_n1276), .B1(new_n1060), .B2(new_n1094), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n1052), .A2(G390), .B1(new_n1280), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1290), .B1(new_n1052), .B2(G390), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1029), .B1(new_n1117), .B2(new_n753), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1051), .B1(new_n1293), .B2(new_n758), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(new_n1005), .A3(G390), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1290), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1280), .A2(new_n1288), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G390), .B1(new_n1294), .B2(new_n1005), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1298), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1292), .A2(new_n1297), .B1(new_n1300), .B2(KEYINPUT125), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1300), .A2(KEYINPUT125), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT60), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1250), .B(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1134), .A2(new_n715), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1273), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n878), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(G384), .A3(new_n1273), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1310), .A2(new_n1311), .B1(G2897), .B2(new_n1285), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1284), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1314), .A2(G2897), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1312), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1217), .A2(G378), .A3(new_n1247), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1215), .A2(new_n758), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1318), .A2(KEYINPUT123), .A3(new_n1246), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT123), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n757), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1246), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1320), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1029), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1206), .A2(new_n1208), .A3(new_n1210), .A4(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1319), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1283), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1314), .B1(new_n1317), .B2(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1303), .B(new_n1304), .C1(new_n1316), .C2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1285), .B1(new_n1317), .B2(new_n1327), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1330), .A2(KEYINPUT63), .A3(new_n1313), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1317), .A2(new_n1327), .ZN(new_n1334));
  AND4_X1   g1134(.A1(KEYINPUT124), .A2(new_n1334), .A3(new_n1284), .A4(new_n1313), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT124), .B1(new_n1328), .B2(new_n1313), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1333), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1332), .A2(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1304), .B1(new_n1316), .B2(new_n1330), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT62), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1340), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1330), .A2(KEYINPUT62), .A3(new_n1313), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1339), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1303), .A2(KEYINPUT127), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT127), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1301), .A2(new_n1345), .A3(new_n1302), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1338), .B1(new_n1343), .B2(new_n1347), .ZN(G405));
  NAND2_X1  g1148(.A1(G375), .A2(new_n1283), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1349), .A2(new_n1317), .ZN(new_n1350));
  XOR2_X1   g1150(.A(new_n1350), .B(new_n1313), .Z(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(new_n1347), .ZN(G402));
endmodule


