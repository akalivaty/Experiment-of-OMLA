//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT92), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n192), .A2(new_n195), .A3(new_n193), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n192), .B2(new_n193), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n194), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT18), .A3(G131), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n204), .A2(KEYINPUT93), .A3(G146), .ZN(new_n205));
  INV_X1    g019(.A(new_n204), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT93), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G146), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT18), .A2(G131), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n194), .B(new_n211), .C1(new_n196), .C2(new_n197), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT16), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n200), .A3(G125), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n204), .B2(new_n214), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n198), .A2(G131), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(new_n194), .C1(new_n196), .C2(new_n197), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n189), .B(new_n213), .C1(new_n220), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n189), .ZN(new_n225));
  OAI211_X1 g039(.A(G146), .B(new_n215), .C1(new_n204), .C2(new_n214), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n204), .B(KEYINPUT19), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(G146), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n228), .B1(new_n218), .B2(new_n222), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n199), .A2(new_n210), .A3(new_n212), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n225), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT94), .ZN(new_n233));
  NOR2_X1   g047(.A1(G475), .A2(G902), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT94), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n224), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NOR3_X1   g051(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n237), .A2(KEYINPUT20), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G475), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT95), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n224), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n213), .B1(new_n220), .B2(new_n223), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n225), .ZN(new_n244));
  AOI21_X1  g058(.A(G902), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(KEYINPUT95), .A3(new_n225), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n240), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT81), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(KEYINPUT81), .ZN(new_n251));
  INV_X1    g065(.A(G107), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G104), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G101), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n188), .A2(G107), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n249), .A2(new_n252), .A3(KEYINPUT81), .A4(G104), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n207), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n193), .A2(G146), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n259), .B(new_n260), .C1(KEYINPUT1), .C2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n193), .B2(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n193), .A2(G146), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n207), .A2(G143), .ZN(new_n265));
  OAI211_X1 g079(.A(G128), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n253), .A2(new_n256), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G101), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n258), .A2(new_n262), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT10), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n262), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n273), .A2(KEYINPUT10), .A3(new_n258), .A4(new_n268), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT82), .ZN(new_n276));
  INV_X1    g090(.A(G137), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G134), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(KEYINPUT11), .A3(G134), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n281), .B1(new_n282), .B2(G137), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G131), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n279), .A2(new_n221), .A3(new_n280), .A4(new_n283), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g104(.A(new_n253), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(KEYINPUT3), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n257), .A2(new_n256), .ZN(new_n294));
  OAI21_X1  g108(.A(G101), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT4), .A3(new_n258), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT64), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n299), .B(new_n300), .C1(new_n264), .C2(new_n265), .ZN(new_n301));
  XNOR2_X1  g115(.A(G143), .B(G146), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT0), .B(G128), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT64), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n297), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n307), .B(G101), .C1(new_n293), .C2(new_n294), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n296), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n275), .A2(new_n276), .A3(new_n288), .A4(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n309), .A2(new_n288), .A3(new_n271), .A4(new_n274), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT82), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n258), .A2(new_n268), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(new_n273), .ZN(new_n316));
  INV_X1    g130(.A(new_n269), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n287), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT12), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(KEYINPUT12), .B(new_n287), .C1(new_n316), .C2(new_n317), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(G110), .B(G140), .ZN(new_n324));
  INV_X1    g138(.A(G227), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  XOR2_X1   g140(.A(new_n324), .B(new_n326), .Z(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n310), .B2(new_n312), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n275), .A2(new_n309), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n287), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n323), .A2(new_n328), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G469), .B1(new_n332), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(G469), .ZN(new_n334));
  INV_X1    g148(.A(G902), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n329), .A2(new_n322), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n327), .B1(new_n313), .B2(new_n331), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n334), .B(new_n335), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n261), .A2(G143), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n193), .A2(G128), .ZN(new_n341));
  OR3_X1    g155(.A1(new_n340), .A2(new_n341), .A3(G134), .ZN(new_n342));
  OAI21_X1  g156(.A(G134), .B1(new_n340), .B2(new_n341), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G122), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G116), .ZN(new_n346));
  INV_X1    g160(.A(G116), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G122), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n252), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n347), .A2(G122), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n348), .B1(new_n352), .B2(KEYINPUT14), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(KEYINPUT14), .B2(new_n348), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT96), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT96), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n357), .A3(G107), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n351), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n349), .B(new_n252), .ZN(new_n360));
  INV_X1    g174(.A(new_n341), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n340), .B1(new_n361), .B2(KEYINPUT13), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n363));
  OAI21_X1  g177(.A(G134), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n360), .A2(new_n364), .A3(new_n342), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  INV_X1    g181(.A(G217), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(G953), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT97), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n359), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n359), .B2(new_n366), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n335), .ZN(new_n374));
  INV_X1    g188(.A(G478), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT15), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g191(.A(new_n373), .B(new_n335), .C1(KEYINPUT15), .C2(new_n375), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G952), .ZN(new_n380));
  AOI211_X1 g194(.A(G953), .B(new_n380), .C1(G234), .C2(G237), .ZN(new_n381));
  AOI211_X1 g195(.A(new_n335), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT21), .B(G898), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(KEYINPUT80), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AND4_X1   g202(.A1(new_n248), .A2(new_n339), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n263), .A2(G128), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(new_n302), .ZN(new_n391));
  INV_X1    g205(.A(new_n262), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n202), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n272), .A2(KEYINPUT86), .A3(new_n202), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G125), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(KEYINPUT87), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(G224), .A3(new_n191), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n191), .A2(G224), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n410));
  INV_X1    g224(.A(G119), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(G116), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G113), .ZN(new_n413));
  XNOR2_X1  g227(.A(G116), .B(G119), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n413), .B1(KEYINPUT5), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT2), .A2(G113), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT65), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT65), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT2), .A3(G113), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(KEYINPUT2), .A2(G113), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n422), .A3(new_n414), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT67), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n421), .B1(new_n417), .B2(new_n419), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n414), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n415), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT84), .B1(new_n428), .B2(new_n315), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n315), .A3(KEYINPUT84), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND4_X1   g246(.A1(new_n426), .A2(new_n420), .A3(new_n422), .A4(new_n414), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n426), .B1(new_n425), .B2(new_n414), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n420), .A2(new_n422), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n437));
  INV_X1    g251(.A(new_n414), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(KEYINPUT66), .B1(new_n425), .B2(new_n414), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT68), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n424), .A2(new_n427), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT68), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n440), .A4(new_n439), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n296), .A2(new_n308), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n432), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(KEYINPUT85), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n438), .A2(new_n410), .ZN(new_n454));
  OAI22_X1  g268(.A1(new_n433), .A2(new_n434), .B1(new_n454), .B2(new_n413), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n455), .A2(new_n456), .A3(new_n314), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n429), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n447), .B1(new_n442), .B2(new_n445), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n453), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n409), .B1(new_n451), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n432), .A2(new_n449), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT6), .B1(new_n462), .B2(new_n453), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n408), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n408), .B(KEYINPUT88), .C1(new_n461), .C2(new_n463), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n395), .B2(new_n396), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT86), .B1(new_n272), .B2(new_n202), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n394), .B(G125), .C1(new_n266), .C2(new_n262), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT89), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n399), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n406), .A2(KEYINPUT7), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n468), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n399), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n395), .A2(new_n469), .A3(new_n396), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT89), .B1(new_n471), .B2(new_n472), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n475), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n480), .A2(KEYINPUT90), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n450), .B(KEYINPUT8), .Z(new_n484));
  NAND2_X1  g298(.A1(new_n455), .A2(new_n314), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n428), .A2(new_n315), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n399), .B(new_n481), .C1(new_n471), .C2(new_n472), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n397), .A2(KEYINPUT91), .A3(new_n399), .A4(new_n481), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n451), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n335), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n466), .A2(new_n467), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G210), .B1(G237), .B2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n494), .B1(new_n464), .B2(new_n465), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n497), .A3(new_n467), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G214), .B1(G237), .B2(G902), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT83), .Z(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n389), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(KEYINPUT23), .B1(new_n261), .B2(G119), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n261), .A2(G119), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT76), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n261), .A2(G119), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT76), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT23), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G110), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT77), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n411), .A2(G128), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT24), .B(G110), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n520), .B(KEYINPUT75), .Z(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(new_n217), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n516), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT78), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(G110), .B2(new_n513), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n526), .B(new_n226), .C1(G146), .C2(new_n204), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G137), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n529), .B(new_n530), .Z(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n523), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT79), .B1(new_n532), .B2(new_n534), .ZN(new_n538));
  OR2_X1    g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n368), .B1(G234), .B2(new_n335), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n540), .A2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n540), .ZN(new_n543));
  AOI21_X1  g357(.A(G902), .B1(new_n532), .B2(new_n534), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n545), .B2(new_n544), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n306), .A2(new_n287), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n282), .A2(G137), .ZN(new_n551));
  OAI21_X1  g365(.A(G131), .B1(new_n551), .B2(new_n278), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n273), .A2(new_n286), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n446), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n446), .A2(KEYINPUT70), .A3(new_n554), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n442), .A2(new_n560), .A3(new_n445), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n560), .B1(new_n442), .B2(new_n445), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n561), .A2(new_n562), .A3(new_n554), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT28), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n561), .A2(new_n562), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n554), .B(KEYINPUT71), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT28), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n190), .A2(new_n191), .A3(G210), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n570), .B(KEYINPUT27), .Z(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT26), .B(G101), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT29), .ZN(new_n576));
  INV_X1    g390(.A(new_n554), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT30), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n550), .A2(new_n578), .A3(new_n553), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n446), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n446), .A2(KEYINPUT69), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n442), .A2(new_n560), .A3(new_n445), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n577), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n576), .B1(new_n587), .B2(new_n573), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n335), .B1(new_n575), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT28), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n554), .B1(new_n561), .B2(new_n562), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(new_n585), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n567), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n574), .A2(new_n576), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT74), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(KEYINPUT74), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(G472), .B1(new_n589), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT32), .ZN(new_n601));
  NOR2_X1   g415(.A1(G472), .A2(G902), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT73), .Z(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  AOI221_X4 g418(.A(new_n556), .B1(new_n550), .B2(new_n553), .C1(new_n442), .C2(new_n445), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT70), .B1(new_n446), .B2(new_n554), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n590), .B1(new_n607), .B2(new_n585), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT72), .B(new_n574), .C1(new_n608), .C2(new_n567), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n582), .A2(new_n585), .A3(new_n573), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT31), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n582), .A2(new_n585), .A3(KEYINPUT31), .A4(new_n573), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT72), .B1(new_n569), .B2(new_n574), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n601), .B(new_n604), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT72), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n585), .A2(new_n557), .A3(new_n558), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n567), .B1(KEYINPUT28), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n619), .B1(new_n621), .B2(new_n573), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n609), .A3(new_n614), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n601), .B1(new_n623), .B2(new_n604), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n600), .B1(new_n618), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n506), .A2(new_n549), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  AOI211_X1 g441(.A(new_n504), .B(new_n384), .C1(new_n499), .C2(new_n501), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n373), .A2(new_n375), .A3(new_n335), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n372), .B2(KEYINPUT98), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n373), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n371), .B(new_n372), .C1(KEYINPUT98), .C2(new_n630), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n629), .B1(new_n634), .B2(new_n375), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n248), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n628), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(G472), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n623), .B2(new_n335), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n604), .B1(new_n615), .B2(new_n616), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n339), .A2(new_n388), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n548), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT34), .B(G104), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  AOI21_X1  g462(.A(new_n504), .B1(new_n499), .B2(new_n501), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT20), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT99), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n237), .A2(new_n653), .A3(KEYINPUT20), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n651), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n384), .ZN(new_n657));
  INV_X1    g471(.A(new_n379), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n247), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n656), .A2(KEYINPUT100), .A3(new_n657), .A4(new_n659), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n649), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT101), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n649), .A2(new_n662), .A3(new_n666), .A4(new_n663), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n645), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT35), .B(G107), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  AOI21_X1  g484(.A(KEYINPUT102), .B1(new_n523), .B2(new_n527), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n523), .A2(KEYINPUT102), .A3(new_n527), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n533), .A2(KEYINPUT36), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n541), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n547), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n639), .A2(new_n641), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n506), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT103), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT37), .B(G110), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  AND4_X1   g499(.A1(new_n497), .A2(new_n466), .A3(new_n467), .A4(new_n495), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n497), .B1(new_n500), .B2(new_n467), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n504), .A3(new_n680), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(new_n625), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n381), .B1(new_n382), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AND3_X1   g507(.A1(new_n656), .A2(new_n659), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n694), .A2(new_n339), .A3(new_n388), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  XNOR2_X1  g511(.A(new_n502), .B(KEYINPUT38), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n640), .A2(KEYINPUT32), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n617), .ZN(new_n700));
  INV_X1    g514(.A(new_n610), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n573), .B1(new_n591), .B2(new_n585), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n335), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G472), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n505), .B(new_n379), .C1(new_n239), .C2(new_n247), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n698), .A2(new_n680), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  XOR2_X1   g525(.A(new_n692), .B(KEYINPUT39), .Z(new_n712));
  AND3_X1   g526(.A1(new_n339), .A2(new_n388), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT40), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n710), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  NAND2_X1  g530(.A1(new_n636), .A2(new_n693), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n643), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n690), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  NAND2_X1  g534(.A1(new_n313), .A2(new_n331), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n721), .A2(new_n328), .B1(new_n329), .B2(new_n322), .ZN(new_n722));
  OAI21_X1  g536(.A(G469), .B1(new_n722), .B2(G902), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n723), .A2(new_n338), .A3(new_n386), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n625), .A2(new_n549), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n637), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT41), .B(G113), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G15));
  AOI21_X1  g542(.A(new_n725), .B1(new_n667), .B2(new_n665), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n347), .ZN(G18));
  AND3_X1   g544(.A1(new_n724), .A2(new_n248), .A3(new_n385), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n689), .A2(new_n625), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G119), .ZN(G21));
  XOR2_X1   g547(.A(KEYINPUT105), .B(G472), .Z(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n623), .B2(new_n335), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n574), .B1(new_n592), .B2(new_n567), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n603), .B1(new_n614), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n735), .A2(new_n548), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n723), .A2(new_n338), .A3(new_n657), .A4(new_n386), .ZN(new_n739));
  AOI211_X1 g553(.A(new_n706), .B(new_n739), .C1(new_n499), .C2(new_n501), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NOR4_X1   g556(.A1(new_n717), .A2(new_n735), .A3(new_n680), .A4(new_n737), .ZN(new_n743));
  INV_X1    g557(.A(new_n724), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n688), .A2(new_n504), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(new_n386), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n748), .B1(new_n333), .B2(new_n338), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n505), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n499), .A2(new_n505), .A3(new_n501), .A4(new_n749), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT106), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n548), .B1(new_n700), .B2(new_n600), .ZN(new_n755));
  INV_X1    g569(.A(new_n717), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n754), .A2(new_n755), .A3(KEYINPUT42), .A4(new_n756), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NAND3_X1  g576(.A1(new_n754), .A2(new_n755), .A3(new_n694), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  NOR2_X1   g578(.A1(new_n502), .A2(new_n504), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n332), .B(KEYINPUT45), .Z(new_n767));
  OAI21_X1  g581(.A(G469), .B1(new_n767), .B2(G902), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n338), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n386), .A3(new_n712), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n642), .A2(new_n680), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(KEYINPUT107), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(KEYINPUT107), .ZN(new_n775));
  INV_X1    g589(.A(new_n635), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n248), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT43), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n766), .B(new_n772), .C1(new_n779), .C2(KEYINPUT44), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(KEYINPUT44), .B2(new_n779), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G137), .ZN(G39));
  NOR4_X1   g596(.A1(new_n766), .A2(new_n625), .A3(new_n549), .A4(new_n717), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT108), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n771), .A2(new_n386), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT47), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NAND2_X1  g602(.A1(new_n549), .A2(new_n381), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n705), .A2(new_n766), .A3(new_n744), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT114), .ZN(new_n791));
  INV_X1    g605(.A(new_n248), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n776), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT115), .ZN(new_n795));
  INV_X1    g609(.A(new_n381), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n778), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n724), .A3(new_n765), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n798), .A2(new_n680), .A3(new_n737), .A4(new_n735), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n698), .A2(new_n505), .A3(new_n744), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n797), .A2(new_n738), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT113), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n802), .B(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n723), .A2(new_n338), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n387), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n786), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n801), .A2(new_n765), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT112), .ZN(new_n810));
  AOI211_X1 g624(.A(new_n799), .B(new_n805), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n795), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n795), .A2(new_n811), .A3(KEYINPUT51), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n801), .A2(new_n745), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(G952), .A3(new_n191), .ZN(new_n817));
  INV_X1    g631(.A(new_n755), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n798), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT48), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n817), .B(new_n820), .C1(new_n636), .C2(new_n791), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n814), .A2(new_n815), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT116), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n689), .B(new_n625), .C1(new_n695), .C2(new_n718), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n680), .A2(new_n693), .A3(new_n749), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n705), .A2(new_n502), .A3(new_n707), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n746), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT111), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT110), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(KEYINPUT111), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT110), .B1(new_n827), .B2(new_n831), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n506), .A2(new_n681), .B1(new_n738), .B2(new_n740), .ZN(new_n835));
  INV_X1    g649(.A(new_n636), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n792), .B2(new_n658), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n628), .A2(new_n642), .A3(new_n644), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n835), .A2(new_n626), .A3(new_n732), .A4(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n729), .A3(new_n726), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n658), .A2(new_n693), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n680), .A2(new_n643), .A3(new_n247), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n625), .A3(new_n656), .A4(new_n765), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n754), .A2(new_n743), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n763), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n759), .B2(new_n760), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n834), .A2(KEYINPUT53), .A3(new_n840), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n827), .B(KEYINPUT52), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT109), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n763), .A2(new_n843), .A3(new_n844), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n761), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n835), .A2(new_n626), .ZN(new_n853));
  INV_X1    g667(.A(new_n726), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n665), .A2(new_n667), .ZN(new_n855));
  INV_X1    g669(.A(new_n725), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n732), .A2(new_n838), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n854), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n850), .B1(new_n852), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n846), .A2(new_n840), .A3(KEYINPUT109), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n849), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n847), .B(new_n848), .C1(new_n862), .C2(KEYINPUT53), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n852), .A2(new_n859), .A3(new_n850), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT109), .B1(new_n846), .B2(new_n840), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n834), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n864), .B2(new_n862), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n863), .B1(new_n868), .B2(new_n848), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n823), .A2(new_n869), .B1(G952), .B2(G953), .ZN(new_n870));
  OR4_X1    g684(.A1(new_n548), .A2(new_n777), .A3(new_n504), .A4(new_n387), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n806), .B(KEYINPUT49), .Z(new_n872));
  OR4_X1    g686(.A1(new_n698), .A2(new_n705), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(new_n873), .ZN(G75));
  OAI21_X1  g688(.A(new_n847), .B1(new_n862), .B2(KEYINPUT53), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(G902), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n875), .B2(G902), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n498), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n461), .A2(new_n463), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(new_n408), .ZN(new_n883));
  XNOR2_X1  g697(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n191), .A2(G952), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n875), .A2(G902), .A3(new_n498), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n885), .B1(new_n889), .B2(new_n881), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n886), .B(new_n888), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(G51));
  NAND2_X1  g709(.A1(new_n767), .A2(G469), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n877), .A2(new_n878), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(G469), .A2(G902), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n899), .B1(new_n900), .B2(new_n863), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n722), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n899), .ZN(new_n904));
  INV_X1    g718(.A(new_n849), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(new_n865), .B2(new_n866), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n864), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n848), .B1(new_n907), .B2(new_n847), .ZN(new_n908));
  INV_X1    g722(.A(new_n863), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT120), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n897), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT121), .B1(new_n912), .B2(new_n887), .ZN(new_n913));
  OR3_X1    g727(.A1(new_n877), .A2(new_n878), .A3(new_n896), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n902), .B(new_n904), .C1(new_n908), .C2(new_n909), .ZN(new_n915));
  INV_X1    g729(.A(new_n722), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n901), .A2(new_n902), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT121), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n888), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n913), .A2(new_n921), .ZN(G54));
  NAND3_X1  g736(.A1(new_n879), .A2(KEYINPUT58), .A3(G475), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n233), .A2(new_n236), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n887), .ZN(G60));
  NAND2_X1  g742(.A1(new_n632), .A2(new_n633), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT122), .Z(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT59), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n930), .B1(new_n869), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n932), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n900), .B2(new_n863), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n933), .A2(new_n887), .A3(new_n935), .ZN(G63));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT60), .Z(new_n939));
  NAND3_X1  g753(.A1(new_n875), .A2(new_n677), .A3(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT123), .Z(new_n941));
  AOI21_X1  g755(.A(new_n539), .B1(new_n875), .B2(new_n939), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(new_n887), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(KEYINPUT124), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n937), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n940), .A2(KEYINPUT61), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n937), .A2(KEYINPUT124), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(G224), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n383), .A2(new_n950), .A3(new_n191), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n859), .B(KEYINPUT125), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n191), .ZN(new_n953));
  INV_X1    g767(.A(G898), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n882), .B1(new_n954), .B2(G953), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n953), .B(new_n955), .Z(G69));
  NOR2_X1   g770(.A1(new_n579), .A2(new_n581), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(new_n227), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n824), .A2(new_n746), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n715), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT62), .Z(new_n961));
  NAND4_X1  g775(.A1(new_n755), .A2(new_n713), .A3(new_n765), .A4(new_n837), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n961), .A2(new_n781), .A3(new_n787), .A4(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n958), .B1(new_n963), .B2(new_n191), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n958), .B1(new_n691), .B2(new_n191), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n787), .A2(new_n959), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n772), .A2(new_n818), .A3(new_n688), .A4(new_n706), .ZN(new_n967));
  INV_X1    g781(.A(new_n763), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND4_X1   g783(.A1(new_n761), .A2(new_n966), .A3(new_n781), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n965), .B1(new_n970), .B2(new_n191), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(G953), .B1(new_n325), .B2(new_n691), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(G72));
  XOR2_X1   g788(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n975));
  NOR2_X1   g789(.A1(new_n638), .A2(new_n335), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n587), .A2(new_n574), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n586), .A2(new_n573), .ZN(new_n979));
  NOR4_X1   g793(.A1(new_n868), .A2(new_n977), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n888), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n970), .A2(new_n979), .ZN(new_n983));
  INV_X1    g797(.A(new_n978), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n963), .B2(new_n984), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n980), .B(new_n982), .C1(new_n985), .C2(new_n952), .ZN(G57));
endmodule


