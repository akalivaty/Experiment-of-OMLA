//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT23), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT73), .B1(new_n189), .B2(G128), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(new_n187), .A3(G119), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n188), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT65), .A2(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(KEYINPUT65), .A2(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(G119), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G110), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(G119), .B2(new_n187), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT72), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT72), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n196), .B(new_n202), .C1(G119), .C2(new_n187), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n208), .B2(KEYINPUT16), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT16), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n210), .A2(new_n207), .A3(KEYINPUT75), .A4(G125), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G125), .B(G140), .ZN(new_n213));
  AOI21_X1  g027(.A(KEYINPUT74), .B1(new_n213), .B2(KEYINPUT16), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G140), .ZN(new_n216));
  AND4_X1   g030(.A1(KEYINPUT74), .A2(new_n208), .A3(new_n216), .A4(KEYINPUT16), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n208), .A2(new_n216), .A3(KEYINPUT16), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT74), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n213), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(G146), .B1(new_n225), .B2(new_n212), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n199), .B(new_n205), .C1(new_n220), .C2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(G146), .A3(new_n212), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n213), .A2(new_n219), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n204), .B1(new_n201), .B2(new_n203), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n198), .A2(G110), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n228), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G953), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(G221), .A3(G234), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n237), .B(KEYINPUT22), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(G137), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n227), .A2(new_n234), .A3(new_n239), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT25), .B1(new_n243), .B2(G902), .ZN(new_n244));
  INV_X1    g058(.A(G217), .ZN(new_n245));
  INV_X1    g059(.A(G902), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n245), .B1(G234), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n241), .A2(new_n248), .A3(new_n246), .A4(new_n242), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n244), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n247), .A2(G902), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n241), .A2(new_n242), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  INV_X1    g068(.A(G116), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G119), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(G119), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n189), .A2(KEYINPUT66), .A3(G116), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G113), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT2), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT2), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G113), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n261), .A2(new_n263), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n266), .A2(new_n257), .A3(new_n258), .A4(new_n256), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT67), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT67), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT11), .ZN(new_n272));
  INV_X1    g086(.A(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n273), .B2(G137), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(G137), .ZN(new_n275));
  INV_X1    g089(.A(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT11), .A3(G134), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G131), .ZN(new_n279));
  INV_X1    g093(.A(G131), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n274), .A2(new_n277), .A3(new_n280), .A4(new_n275), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n219), .A2(G143), .ZN(new_n283));
  AND2_X1   g097(.A1(KEYINPUT0), .A2(G128), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT64), .B(G143), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n219), .ZN(new_n286));
  INV_X1    g100(.A(G143), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT64), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G143), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n290), .A3(new_n219), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(G146), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n282), .A2(new_n286), .A3(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n276), .A2(G134), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n273), .A2(G137), .ZN(new_n299));
  OAI21_X1  g113(.A(G131), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n281), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n219), .B1(new_n288), .B2(new_n290), .ZN(new_n302));
  INV_X1    g116(.A(new_n283), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n194), .A2(new_n195), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n283), .A2(KEYINPUT1), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n291), .A2(new_n292), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n301), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AOI211_X1 g124(.A(KEYINPUT68), .B(new_n271), .C1(new_n297), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT30), .ZN(new_n314));
  AND4_X1   g128(.A1(new_n297), .A2(new_n310), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n270), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n297), .B(new_n310), .C1(new_n268), .C2(new_n269), .ZN(new_n317));
  XOR2_X1   g131(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n318));
  NOR2_X1   g132(.A1(G237), .A2(G953), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G210), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n318), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT26), .B(G101), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n316), .A2(new_n317), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT31), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n297), .A2(new_n310), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n270), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(new_n317), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n317), .A2(new_n327), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G472), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n316), .A2(KEYINPUT31), .A3(new_n317), .A4(new_n324), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n246), .A4(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT32), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n246), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n340), .A2(KEYINPUT32), .A3(new_n334), .A4(new_n333), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(KEYINPUT70), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT70), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(new_n343), .A3(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n265), .A2(new_n267), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT67), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(new_n297), .B2(new_n310), .ZN(new_n351));
  INV_X1    g165(.A(new_n317), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT28), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n331), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n324), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n328), .A2(new_n313), .A3(KEYINPUT30), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n297), .A2(new_n310), .A3(new_n312), .A4(new_n314), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n350), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n323), .B1(new_n358), .B2(new_n352), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT29), .A4(new_n324), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n246), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G472), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT71), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n366), .A3(G472), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n253), .B1(new_n345), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT87), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n220), .B2(new_n226), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n288), .A2(new_n290), .B1(new_n319), .B2(G214), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n319), .A2(G143), .A3(G214), .ZN(new_n373));
  OAI21_X1  g187(.A(G131), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n319), .A2(G143), .A3(G214), .ZN(new_n376));
  INV_X1    g190(.A(G214), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n377), .A2(G237), .A3(G953), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n280), .B(new_n376), .C1(new_n285), .C2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n372), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n381), .A2(KEYINPUT84), .A3(new_n280), .A4(new_n376), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n374), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n218), .A2(new_n219), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT87), .A3(new_n228), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n371), .A2(new_n385), .A3(new_n387), .A4(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n231), .B1(new_n219), .B2(new_n213), .ZN(new_n394));
  OR3_X1    g208(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT18), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n379), .A4(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n390), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n393), .B1(new_n390), .B2(new_n397), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n246), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G475), .ZN(new_n401));
  NOR2_X1   g215(.A1(G475), .A2(G902), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n383), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT86), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n213), .A2(new_n405), .A3(KEYINPUT19), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT19), .B1(new_n213), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n219), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n228), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT85), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n404), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n393), .B1(new_n411), .B2(new_n397), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n402), .B1(new_n398), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n412), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n390), .A2(new_n393), .A3(new_n397), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT20), .A3(new_n402), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n401), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n195), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT65), .A2(G128), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n287), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n187), .B1(new_n288), .B2(new_n290), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n273), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G143), .B1(new_n194), .B2(new_n195), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(G134), .C1(new_n187), .C2(new_n285), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT13), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n428), .A3(G134), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G122), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n255), .A2(G122), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT88), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT88), .B1(new_n432), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g249(.A(G107), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n433), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G107), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT88), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n424), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n444), .A2(new_n428), .A3(G134), .A4(new_n426), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n430), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n255), .A2(KEYINPUT14), .A3(G122), .ZN(new_n447));
  OAI211_X1 g261(.A(G107), .B(new_n447), .C1(new_n437), .C2(KEYINPUT14), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n425), .A2(new_n442), .A3(new_n427), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(new_n245), .A3(G953), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n452), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n449), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n453), .A2(new_n246), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n459));
  OR2_X1    g273(.A1(new_n459), .A2(KEYINPUT15), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(KEYINPUT15), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G478), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n453), .A2(KEYINPUT90), .A3(new_n246), .A4(new_n455), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n456), .A2(new_n457), .A3(new_n462), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n420), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G214), .B1(G237), .B2(G902), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n440), .A2(KEYINPUT77), .A3(G104), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n392), .A2(G107), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n473), .A2(new_n440), .A3(KEYINPUT77), .A4(G104), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g290(.A(G101), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n471), .A2(new_n477), .A3(new_n472), .A4(new_n474), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(KEYINPUT4), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n475), .A2(new_n480), .A3(G101), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n479), .A2(new_n348), .A3(new_n481), .A4(new_n349), .ZN(new_n482));
  INV_X1    g296(.A(new_n472), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n392), .A2(G107), .ZN(new_n484));
  OAI21_X1  g298(.A(G101), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT78), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT78), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n478), .A2(new_n488), .A3(new_n485), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT5), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n189), .A3(G116), .ZN(new_n491));
  OAI211_X1 g305(.A(G113), .B(new_n491), .C1(new_n259), .C2(new_n490), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n489), .A3(new_n267), .A4(new_n492), .ZN(new_n493));
  XNOR2_X1  g307(.A(G110), .B(G122), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n494), .B(KEYINPUT8), .Z(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n267), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n486), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n497), .B1(new_n493), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n306), .A2(new_n309), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n215), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n296), .A2(new_n286), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G125), .ZN(new_n505));
  NAND2_X1  g319(.A1(KEYINPUT82), .A2(KEYINPUT7), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G224), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n508), .A2(G953), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n507), .B(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n501), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n482), .A2(new_n493), .ZN(new_n514));
  INV_X1    g328(.A(new_n494), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n495), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n503), .A2(new_n505), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n509), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n514), .A2(new_n520), .A3(new_n515), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(G210), .B1(G237), .B2(G902), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n513), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n523), .B1(new_n513), .B2(new_n522), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n469), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT83), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G952), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(G953), .ZN(new_n530));
  NAND2_X1  g344(.A1(G234), .A2(G237), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  XOR2_X1   g347(.A(KEYINPUT21), .B(G898), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n531), .A2(G902), .A3(G953), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(KEYINPUT83), .B(new_n469), .C1(new_n524), .C2(new_n525), .ZN(new_n540));
  AND4_X1   g354(.A1(new_n468), .A2(new_n528), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G221), .B1(new_n451), .B2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  XOR2_X1   g357(.A(G110), .B(G140), .Z(new_n544));
  INV_X1    g358(.A(G227), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n544), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n478), .A2(new_n488), .A3(new_n485), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n488), .B1(new_n478), .B2(new_n485), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n502), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n283), .B(new_n304), .C1(new_n285), .C2(new_n219), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n187), .B1(new_n291), .B2(KEYINPUT1), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n302), .A2(new_n303), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n486), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n502), .B(KEYINPUT80), .C1(new_n549), .C2(new_n550), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n553), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n561), .A2(KEYINPUT12), .A3(new_n282), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT12), .B1(new_n561), .B2(new_n282), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT10), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n307), .A2(new_n308), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n293), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n566), .B2(new_n554), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n487), .A3(new_n489), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT79), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n559), .A2(new_n564), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n296), .A2(new_n286), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n571), .A2(new_n479), .A3(new_n481), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT79), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n567), .A2(new_n487), .A3(new_n573), .A4(new_n489), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n569), .A2(new_n570), .A3(new_n572), .A4(new_n574), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n562), .A2(new_n563), .B1(new_n282), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n549), .A2(new_n550), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(new_n577), .B2(new_n567), .ZN(new_n578));
  AND4_X1   g392(.A1(new_n573), .A2(new_n567), .A3(new_n487), .A4(new_n489), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n479), .A2(new_n481), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n581), .A2(new_n571), .B1(new_n564), .B2(new_n559), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT81), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n569), .A2(new_n574), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT81), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n572), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n282), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n575), .A2(new_n282), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n589), .A2(new_n548), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n548), .A2(new_n576), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G469), .B1(new_n591), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n282), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n575), .A2(new_n585), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n582), .A2(KEYINPUT81), .A3(new_n569), .A4(new_n574), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n548), .B1(new_n596), .B2(new_n589), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n590), .B1(new_n562), .B2(new_n563), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(G469), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n599), .A2(new_n600), .A3(new_n246), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n543), .B1(new_n592), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n369), .A2(new_n541), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT91), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(new_n477), .ZN(G3));
  AND3_X1   g419(.A1(new_n325), .A2(new_n326), .A3(new_n332), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT92), .B1(new_n606), .B2(new_n339), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n340), .A2(new_n608), .A3(new_n333), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT93), .A4(G472), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n607), .A2(new_n609), .A3(G472), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n336), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n576), .A2(new_n548), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n588), .A2(new_n590), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n600), .B1(new_n618), .B2(new_n246), .ZN(new_n619));
  AOI211_X1 g433(.A(G469), .B(G902), .C1(new_n597), .C2(new_n598), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n542), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n250), .A2(new_n252), .ZN(new_n623));
  INV_X1    g437(.A(new_n526), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n539), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n453), .A2(new_n626), .A3(new_n455), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n453), .A2(KEYINPUT94), .A3(new_n626), .A4(new_n455), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n454), .B1(new_n450), .B2(new_n631), .ZN(new_n632));
  AOI211_X1 g446(.A(KEYINPUT95), .B(new_n452), .C1(new_n446), .C2(new_n449), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n629), .A2(new_n630), .B1(new_n634), .B2(KEYINPUT33), .ZN(new_n635));
  INV_X1    g449(.A(G478), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n456), .A2(new_n636), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n420), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n625), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n622), .A2(new_n623), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT96), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n644), .B(new_n646), .ZN(G6));
  NAND4_X1  g461(.A1(new_n467), .A2(new_n401), .A3(new_n415), .A4(new_n419), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n625), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n622), .A2(new_n623), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT97), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n650), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n240), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n235), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n251), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n250), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n541), .A2(new_n614), .A3(new_n602), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G110), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(new_n657), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n345), .B2(new_n368), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n536), .A2(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n532), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT99), .B1(new_n648), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n401), .A2(new_n415), .A3(new_n419), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(new_n669), .A3(new_n467), .A4(new_n665), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  AOI211_X1 g485(.A(new_n543), .B(new_n526), .C1(new_n592), .C2(new_n601), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n663), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  XOR2_X1   g488(.A(new_n665), .B(KEYINPUT103), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT39), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n602), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT104), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT40), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n334), .A2(new_n246), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n324), .B1(new_n329), .B2(new_n317), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n683), .B2(KEYINPUT100), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n358), .A2(new_n352), .A3(new_n323), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT100), .ZN(new_n687));
  AOI211_X1 g501(.A(new_n687), .B(new_n324), .C1(new_n317), .C2(new_n329), .ZN(new_n688));
  OAI211_X1 g502(.A(new_n680), .B(new_n682), .C1(new_n686), .C2(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n690));
  OAI21_X1  g504(.A(KEYINPUT101), .B1(new_n690), .B2(new_n681), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n342), .B2(new_n344), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n524), .A2(new_n525), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT38), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n662), .A2(new_n467), .A3(new_n420), .A4(new_n469), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT102), .Z(new_n698));
  NAND3_X1  g512(.A1(new_n679), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n285), .ZN(G45));
  NAND2_X1  g514(.A1(new_n345), .A2(new_n368), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n642), .A2(new_n666), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n672), .A2(new_n701), .A3(new_n657), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  AOI21_X1  g518(.A(new_n600), .B1(new_n599), .B2(new_n246), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n620), .A3(new_n543), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n369), .A2(new_n643), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND3_X1  g523(.A1(new_n369), .A2(new_n649), .A3(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NOR4_X1   g525(.A1(new_n705), .A2(new_n620), .A3(new_n543), .A4(new_n526), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n663), .A2(new_n712), .A3(new_n468), .A4(new_n539), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n420), .A2(new_n715), .A3(new_n467), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n715), .B1(new_n420), .B2(new_n467), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n716), .A2(new_n717), .A3(new_n526), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n606), .B2(new_n339), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n336), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n719), .B1(new_n721), .B2(new_n253), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n623), .A2(KEYINPUT105), .A3(new_n336), .A4(new_n720), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n718), .A2(new_n539), .A3(new_n706), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR2_X1   g540(.A1(new_n662), .A2(new_n721), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n706), .A2(new_n624), .A3(new_n727), .A4(new_n702), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n694), .A2(new_n469), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n730), .B1(new_n621), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n731), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n602), .A2(KEYINPUT107), .A3(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n369), .A3(new_n702), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n368), .A2(new_n338), .A3(new_n341), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(KEYINPUT42), .A3(new_n623), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n702), .A3(new_n732), .A4(new_n734), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  NAND4_X1  g556(.A1(new_n732), .A2(new_n369), .A3(new_n671), .A4(new_n734), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  XNOR2_X1  g558(.A(new_n618), .B(KEYINPUT45), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(G469), .ZN(new_n746));
  NAND2_X1  g560(.A1(G469), .A2(G902), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT46), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n620), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n746), .A2(KEYINPUT46), .A3(new_n747), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n543), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT108), .B1(new_n668), .B2(new_n641), .ZN(new_n754));
  XOR2_X1   g568(.A(new_n754), .B(KEYINPUT43), .Z(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n615), .A3(new_n657), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n752), .B(new_n676), .C1(new_n753), .C2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n756), .A2(new_n753), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n731), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n276), .ZN(G39));
  NAND2_X1  g574(.A1(new_n750), .A2(new_n751), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT47), .B1(new_n761), .B2(new_n542), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT47), .ZN(new_n763));
  AOI211_X1 g577(.A(new_n763), .B(new_n543), .C1(new_n750), .C2(new_n751), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n765), .A2(new_n642), .A3(new_n666), .A4(new_n731), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n701), .A2(new_n623), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  NAND2_X1  g583(.A1(new_n755), .A2(new_n533), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n738), .A2(new_n623), .ZN(new_n772));
  INV_X1    g586(.A(new_n706), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n731), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT48), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n236), .A2(G952), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n623), .A3(new_n533), .A4(new_n693), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n642), .ZN(new_n779));
  INV_X1    g593(.A(new_n724), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n770), .A2(new_n780), .ZN(new_n781));
  AOI211_X1 g595(.A(new_n777), .B(new_n779), .C1(new_n712), .C2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n776), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n776), .B2(new_n782), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n705), .A2(new_n620), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n787), .B(KEYINPUT110), .Z(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n543), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n731), .B1(new_n765), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n469), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n780), .A2(new_n773), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n771), .A2(new_n791), .A3(new_n695), .A4(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n790), .A2(new_n781), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n778), .A2(new_n420), .A3(new_n641), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n771), .A2(new_n727), .A3(new_n774), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT118), .Z(new_n801));
  NAND4_X1  g615(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n762), .ZN(new_n803));
  INV_X1    g617(.A(new_n764), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n789), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n733), .A3(new_n781), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n796), .A2(new_n795), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n806), .A2(new_n801), .A3(new_n799), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n786), .B1(new_n802), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n692), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n345), .A2(new_n811), .ZN(new_n812));
  OR3_X1    g626(.A1(new_n657), .A2(KEYINPUT112), .A3(new_n666), .ZN(new_n813));
  OAI21_X1  g627(.A(KEYINPUT112), .B1(new_n657), .B2(new_n666), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n718), .A2(new_n812), .A3(new_n602), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n693), .A2(new_n621), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(KEYINPUT113), .A3(new_n718), .A4(new_n815), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n673), .A2(new_n703), .A3(new_n728), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT52), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n821), .A2(new_n822), .A3(KEYINPUT52), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(new_n821), .B2(new_n822), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n825), .B1(new_n828), .B2(new_n824), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n528), .A2(new_n539), .A3(new_n540), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n642), .A2(new_n648), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n602), .A3(new_n623), .A4(new_n614), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n603), .A3(new_n658), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT111), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT111), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n658), .A3(new_n603), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n713), .A2(new_n707), .A3(new_n710), .A4(new_n725), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n737), .B2(new_n740), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n621), .A2(new_n731), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n701), .A3(new_n468), .A4(new_n665), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n732), .A2(new_n702), .A3(new_n734), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n842), .B1(new_n843), .B2(new_n721), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n657), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n838), .A2(new_n840), .A3(new_n743), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT53), .B1(new_n829), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n846), .A2(new_n828), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT54), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n846), .B2(new_n828), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n821), .A2(new_n822), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n824), .A3(new_n823), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n826), .A2(KEYINPUT114), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n840), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n839), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n741), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT117), .ZN(new_n865));
  INV_X1    g679(.A(new_n743), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n835), .B2(new_n837), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n845), .A4(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n853), .B(new_n854), .C1(new_n862), .C2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT116), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n852), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(KEYINPUT116), .B(KEYINPUT54), .C1(new_n848), .C2(new_n851), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n810), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n529), .A2(new_n236), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n810), .A2(new_n871), .A3(KEYINPUT120), .A4(new_n872), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n788), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT49), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n668), .A2(new_n542), .A3(new_n641), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n881), .A2(new_n253), .A3(new_n791), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(KEYINPUT109), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n879), .B2(KEYINPUT49), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n812), .B1(new_n882), .B2(KEYINPUT109), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n880), .A2(new_n884), .A3(new_n695), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n878), .A2(new_n886), .ZN(G75));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n853), .B1(new_n862), .B2(new_n868), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G902), .ZN(new_n890));
  INV_X1    g704(.A(G210), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n517), .A2(new_n521), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(new_n519), .Z(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n892), .A2(new_n895), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n236), .A2(G952), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n889), .A2(KEYINPUT54), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n869), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n747), .B(KEYINPUT57), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n901), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n599), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n890), .A2(new_n746), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n898), .B1(new_n908), .B2(new_n909), .ZN(G54));
  NAND4_X1  g724(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(new_n418), .Z(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n898), .ZN(G60));
  NAND2_X1  g727(.A1(new_n871), .A2(new_n872), .ZN(new_n914));
  XNOR2_X1  g728(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n636), .A2(new_n246), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n915), .B(new_n916), .Z(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n635), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n901), .A2(new_n635), .A3(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n898), .A3(new_n920), .ZN(G63));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT60), .Z(new_n924));
  AND3_X1   g738(.A1(new_n889), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n889), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n898), .B1(new_n927), .B2(new_n243), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n655), .B1(new_n925), .B2(new_n926), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n928), .B(new_n929), .C1(KEYINPUT124), .C2(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n889), .A2(new_n924), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT123), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n889), .A2(new_n922), .A3(new_n924), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n243), .A3(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n898), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n934), .A2(KEYINPUT124), .A3(new_n935), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n930), .A2(new_n939), .ZN(G66));
  NAND2_X1  g754(.A1(new_n838), .A2(new_n863), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT125), .Z(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n236), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n535), .B2(new_n508), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n893), .B1(G898), .B2(new_n236), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G69));
  NAND2_X1  g761(.A1(new_n699), .A2(new_n822), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  INV_X1    g763(.A(new_n369), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(new_n831), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n831), .A2(new_n951), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n678), .A2(new_n733), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n759), .B1(new_n766), .B2(new_n767), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n949), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n356), .A2(new_n357), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n406), .A2(new_n407), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n956), .A2(new_n236), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(G900), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n959), .B2(new_n545), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n963));
  INV_X1    g777(.A(new_n822), .ZN(new_n964));
  OR3_X1    g778(.A1(new_n759), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n759), .B2(new_n964), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n866), .B1(new_n766), .B2(new_n767), .ZN(new_n968));
  AND4_X1   g782(.A1(new_n676), .A2(new_n752), .A3(new_n718), .A4(new_n772), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n967), .A2(new_n968), .A3(new_n741), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n236), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(G227), .B2(new_n236), .ZN(new_n973));
  OAI221_X1 g787(.A(new_n960), .B1(new_n236), .B2(new_n962), .C1(new_n973), .C2(new_n959), .ZN(G72));
  XNOR2_X1  g788(.A(new_n681), .B(KEYINPUT63), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n956), .B2(new_n942), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n316), .A2(new_n317), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n978), .A2(new_n323), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n975), .B1(new_n971), .B2(new_n942), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n977), .A2(new_n324), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n898), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n848), .A2(new_n851), .ZN(new_n984));
  INV_X1    g798(.A(new_n979), .ZN(new_n985));
  INV_X1    g799(.A(new_n982), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n984), .A2(new_n975), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n980), .A2(new_n983), .A3(new_n987), .ZN(G57));
endmodule


