

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U323 ( .A(n365), .B(n364), .ZN(n385) );
  NAND2_X1 U324 ( .A1(n470), .A2(n469), .ZN(n484) );
  XNOR2_X1 U325 ( .A(n418), .B(n291), .ZN(n323) );
  XOR2_X1 U326 ( .A(n310), .B(n309), .Z(n557) );
  XOR2_X1 U327 ( .A(G99GAT), .B(G190GAT), .Z(n291) );
  XOR2_X1 U328 ( .A(G134GAT), .B(G106GAT), .Z(n292) );
  XOR2_X1 U329 ( .A(G92GAT), .B(KEYINPUT72), .Z(n293) );
  XOR2_X1 U330 ( .A(n329), .B(KEYINPUT64), .Z(n294) );
  XNOR2_X1 U331 ( .A(n363), .B(KEYINPUT111), .ZN(n364) );
  INV_X1 U332 ( .A(KEYINPUT31), .ZN(n326) );
  XNOR2_X1 U333 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U334 ( .A(G15GAT), .B(G127GAT), .Z(n367) );
  XNOR2_X1 U335 ( .A(n301), .B(n292), .ZN(n302) );
  NOR2_X1 U336 ( .A1(n583), .A2(n486), .ZN(n487) );
  XNOR2_X1 U337 ( .A(n458), .B(KEYINPUT26), .ZN(n568) );
  XNOR2_X1 U338 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U339 ( .A(n324), .B(n323), .ZN(n325) );
  NOR2_X1 U340 ( .A1(n518), .A2(n450), .ZN(n561) );
  XNOR2_X1 U341 ( .A(n512), .B(KEYINPUT107), .ZN(n522) );
  INV_X1 U342 ( .A(n527), .ZN(n518) );
  XNOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n451) );
  XNOR2_X1 U344 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n296) );
  XNOR2_X1 U346 ( .A(KEYINPUT9), .B(KEYINPUT76), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n305) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G85GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n293), .B(n297), .ZN(n329) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n294), .B(n298), .ZN(n303) );
  XOR2_X1 U352 ( .A(G36GAT), .B(G190GAT), .Z(n402) );
  XOR2_X1 U353 ( .A(KEYINPUT75), .B(n402), .Z(n300) );
  XOR2_X1 U354 ( .A(G50GAT), .B(G162GAT), .Z(n444) );
  XNOR2_X1 U355 ( .A(G218GAT), .B(n444), .ZN(n299) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n305), .B(n304), .ZN(n310) );
  XOR2_X1 U358 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n307) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G29GAT), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U361 ( .A(KEYINPUT67), .B(n308), .ZN(n358) );
  INV_X1 U362 ( .A(n358), .ZN(n309) );
  XOR2_X1 U363 ( .A(KEYINPUT82), .B(KEYINPUT18), .Z(n312) );
  XNOR2_X1 U364 ( .A(KEYINPUT19), .B(KEYINPUT83), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U366 ( .A(n313), .B(KEYINPUT17), .Z(n315) );
  XNOR2_X1 U367 ( .A(G169GAT), .B(G183GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n408) );
  XOR2_X1 U369 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n317) );
  XNOR2_X1 U370 ( .A(G43GAT), .B(G113GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(G120GAT), .B(G71GAT), .Z(n334) );
  XNOR2_X1 U373 ( .A(n318), .B(n334), .ZN(n322) );
  XOR2_X1 U374 ( .A(n367), .B(G176GAT), .Z(n320) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U378 ( .A(G134GAT), .B(KEYINPUT0), .Z(n418) );
  XNOR2_X1 U379 ( .A(n408), .B(n325), .ZN(n527) );
  XNOR2_X1 U380 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n394) );
  NAND2_X1 U381 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U383 ( .A(KEYINPUT74), .B(KEYINPUT70), .Z(n331) );
  XNOR2_X1 U384 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(n333), .B(n332), .Z(n336) );
  XOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT13), .Z(n366) );
  XNOR2_X1 U388 ( .A(n334), .B(n366), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U390 ( .A(G78GAT), .B(G148GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n435) );
  XOR2_X1 U393 ( .A(G64GAT), .B(KEYINPUT73), .Z(n340) );
  XNOR2_X1 U394 ( .A(G176GAT), .B(G204GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n401) );
  XNOR2_X1 U396 ( .A(n435), .B(n401), .ZN(n342) );
  NAND2_X1 U397 ( .A1(n341), .A2(n342), .ZN(n346) );
  INV_X1 U398 ( .A(n341), .ZN(n344) );
  INV_X1 U399 ( .A(n342), .ZN(n343) );
  NAND2_X1 U400 ( .A1(n344), .A2(n343), .ZN(n345) );
  NAND2_X1 U401 ( .A1(n346), .A2(n345), .ZN(n573) );
  XOR2_X1 U402 ( .A(KEYINPUT41), .B(n573), .Z(n550) );
  XOR2_X1 U403 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n348) );
  XNOR2_X1 U404 ( .A(G15GAT), .B(KEYINPUT29), .ZN(n347) );
  XNOR2_X1 U405 ( .A(n348), .B(n347), .ZN(n362) );
  XOR2_X1 U406 ( .A(G22GAT), .B(G141GAT), .Z(n350) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G50GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U409 ( .A(n351), .B(G197GAT), .Z(n353) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G1GAT), .Z(n413) );
  XNOR2_X1 U411 ( .A(G169GAT), .B(n413), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U413 ( .A(KEYINPUT66), .B(KEYINPUT69), .Z(n355) );
  NAND2_X1 U414 ( .A1(G229GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U416 ( .A(n357), .B(n356), .Z(n360) );
  XOR2_X1 U417 ( .A(KEYINPUT68), .B(G8GAT), .Z(n374) );
  XOR2_X1 U418 ( .A(n358), .B(n374), .Z(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n529) );
  INV_X1 U421 ( .A(n529), .ZN(n570) );
  NAND2_X1 U422 ( .A1(n550), .A2(n570), .ZN(n365) );
  XOR2_X1 U423 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n363) );
  XOR2_X1 U424 ( .A(n366), .B(G78GAT), .Z(n369) );
  XNOR2_X1 U425 ( .A(n367), .B(G211GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U427 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n371) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U430 ( .A(n373), .B(n372), .Z(n376) );
  XOR2_X1 U431 ( .A(G22GAT), .B(G155GAT), .Z(n443) );
  XNOR2_X1 U432 ( .A(n374), .B(n443), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n384) );
  XOR2_X1 U434 ( .A(G64GAT), .B(G71GAT), .Z(n378) );
  XNOR2_X1 U435 ( .A(G1GAT), .B(G183GAT), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n380) );
  XNOR2_X1 U438 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U440 ( .A(n382), .B(n381), .Z(n383) );
  XOR2_X1 U441 ( .A(n384), .B(n383), .Z(n576) );
  INV_X1 U442 ( .A(n576), .ZN(n536) );
  NAND2_X1 U443 ( .A1(n385), .A2(n536), .ZN(n386) );
  NOR2_X1 U444 ( .A1(n557), .A2(n386), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n387), .B(KEYINPUT47), .ZN(n392) );
  XOR2_X1 U446 ( .A(KEYINPUT36), .B(n557), .Z(n583) );
  NOR2_X1 U447 ( .A1(n583), .A2(n536), .ZN(n388) );
  XOR2_X1 U448 ( .A(KEYINPUT45), .B(n388), .Z(n389) );
  NOR2_X1 U449 ( .A1(n573), .A2(n389), .ZN(n390) );
  NAND2_X1 U450 ( .A1(n390), .A2(n529), .ZN(n391) );
  NAND2_X1 U451 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n544) );
  XOR2_X1 U453 ( .A(KEYINPUT88), .B(G218GAT), .Z(n396) );
  XNOR2_X1 U454 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U456 ( .A(G197GAT), .B(n397), .Z(n448) );
  XOR2_X1 U457 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n399) );
  XNOR2_X1 U458 ( .A(G8GAT), .B(G92GAT), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n448), .B(n400), .ZN(n406) );
  XOR2_X1 U461 ( .A(n402), .B(n401), .Z(n404) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n516) );
  NOR2_X1 U466 ( .A1(n544), .A2(n516), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n409), .B(KEYINPUT54), .ZN(n431) );
  XOR2_X1 U468 ( .A(G85GAT), .B(G162GAT), .Z(n411) );
  XNOR2_X1 U469 ( .A(G120GAT), .B(G148GAT), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U471 ( .A(n412), .B(G155GAT), .Z(n415) );
  XNOR2_X1 U472 ( .A(G29GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n422) );
  XOR2_X1 U474 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n417) );
  XNOR2_X1 U475 ( .A(G141GAT), .B(KEYINPUT89), .ZN(n416) );
  XNOR2_X1 U476 ( .A(n417), .B(n416), .ZN(n436) );
  XOR2_X1 U477 ( .A(n436), .B(n418), .Z(n420) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U480 ( .A(n422), .B(n421), .Z(n430) );
  XOR2_X1 U481 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n424) );
  XNOR2_X1 U482 ( .A(G127GAT), .B(G57GAT), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U484 ( .A(KEYINPUT4), .B(KEYINPUT90), .Z(n426) );
  XNOR2_X1 U485 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n513) );
  NAND2_X1 U489 ( .A1(n431), .A2(n513), .ZN(n567) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n433) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U493 ( .A(n434), .B(KEYINPUT22), .Z(n438) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U496 ( .A(G204GAT), .B(KEYINPUT86), .Z(n440) );
  XNOR2_X1 U497 ( .A(KEYINPUT23), .B(KEYINPUT85), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U499 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n467) );
  NOR2_X1 U503 ( .A1(n567), .A2(n467), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  NAND2_X1 U505 ( .A1(n557), .A2(n561), .ZN(n452) );
  NAND2_X1 U506 ( .A1(n561), .A2(n550), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  XNOR2_X1 U508 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XOR2_X1 U510 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n457) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n457), .B(n456), .ZN(n476) );
  NOR2_X1 U513 ( .A1(n573), .A2(n529), .ZN(n488) );
  XNOR2_X1 U514 ( .A(KEYINPUT27), .B(n516), .ZN(n465) );
  NAND2_X1 U515 ( .A1(n467), .A2(n518), .ZN(n458) );
  NOR2_X1 U516 ( .A1(n465), .A2(n568), .ZN(n459) );
  XOR2_X1 U517 ( .A(KEYINPUT96), .B(n459), .Z(n463) );
  NOR2_X1 U518 ( .A1(n518), .A2(n516), .ZN(n460) );
  NOR2_X1 U519 ( .A1(n467), .A2(n460), .ZN(n461) );
  XNOR2_X1 U520 ( .A(KEYINPUT25), .B(n461), .ZN(n462) );
  NAND2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n464), .A2(n513), .ZN(n470) );
  NOR2_X1 U523 ( .A1(n465), .A2(n513), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n466), .B(KEYINPUT94), .ZN(n546) );
  XOR2_X1 U525 ( .A(KEYINPUT28), .B(n467), .Z(n523) );
  NAND2_X1 U526 ( .A1(n546), .A2(n523), .ZN(n526) );
  XNOR2_X1 U527 ( .A(KEYINPUT95), .B(n526), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n518), .A2(n468), .ZN(n469) );
  XOR2_X1 U529 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n472) );
  INV_X1 U530 ( .A(n557), .ZN(n541) );
  NAND2_X1 U531 ( .A1(n576), .A2(n541), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  AND2_X1 U534 ( .A1(n484), .A2(n474), .ZN(n499) );
  NAND2_X1 U535 ( .A1(n488), .A2(n499), .ZN(n482) );
  NOR2_X1 U536 ( .A1(n513), .A2(n482), .ZN(n475) );
  XOR2_X1 U537 ( .A(n476), .B(n475), .Z(G1324GAT) );
  NOR2_X1 U538 ( .A1(n516), .A2(n482), .ZN(n477) );
  XOR2_X1 U539 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U540 ( .A1(n482), .A2(n518), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n479) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT100), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U545 ( .A1(n523), .A2(n482), .ZN(n483) );
  XOR2_X1 U546 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  NAND2_X1 U548 ( .A1(n536), .A2(n484), .ZN(n485) );
  XOR2_X1 U549 ( .A(KEYINPUT101), .B(n485), .Z(n486) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(n487), .Z(n511) );
  NAND2_X1 U551 ( .A1(n511), .A2(n488), .ZN(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT38), .B(n489), .ZN(n497) );
  NOR2_X1 U553 ( .A1(n513), .A2(n497), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U555 ( .A1(n497), .A2(n516), .ZN(n492) );
  XOR2_X1 U556 ( .A(KEYINPUT102), .B(n492), .Z(n493) );
  XNOR2_X1 U557 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n495) );
  NOR2_X1 U559 ( .A1(n518), .A2(n497), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n496), .ZN(G1330GAT) );
  NOR2_X1 U562 ( .A1(n497), .A2(n523), .ZN(n498) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n498), .Z(G1331GAT) );
  INV_X1 U564 ( .A(n550), .ZN(n531) );
  NOR2_X1 U565 ( .A1(n570), .A2(n531), .ZN(n510) );
  NAND2_X1 U566 ( .A1(n510), .A2(n499), .ZN(n505) );
  NOR2_X1 U567 ( .A1(n513), .A2(n505), .ZN(n501) );
  XNOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT104), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U570 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NOR2_X1 U571 ( .A1(n516), .A2(n505), .ZN(n503) );
  XOR2_X1 U572 ( .A(G64GAT), .B(n503), .Z(G1333GAT) );
  NOR2_X1 U573 ( .A1(n518), .A2(n505), .ZN(n504) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n504), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n505), .A2(n523), .ZN(n509) );
  XOR2_X1 U576 ( .A(KEYINPUT105), .B(KEYINPUT43), .Z(n507) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U578 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U579 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  AND2_X1 U580 ( .A1(n511), .A2(n510), .ZN(n512) );
  NOR2_X1 U581 ( .A1(n513), .A2(n522), .ZN(n514) );
  XOR2_X1 U582 ( .A(n514), .B(KEYINPUT108), .Z(n515) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n516), .A2(n522), .ZN(n517) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n518), .A2(n522), .ZN(n519) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n521) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U590 ( .A(n521), .B(n520), .ZN(n525) );
  NOR2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U592 ( .A(n525), .B(n524), .Z(G1339GAT) );
  NOR2_X1 U593 ( .A1(n544), .A2(n526), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n529), .A2(n540), .ZN(n530) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  NOR2_X1 U597 ( .A1(n540), .A2(n531), .ZN(n535) );
  XOR2_X1 U598 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n533) );
  XNOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U602 ( .A1(n536), .A2(n540), .ZN(n538) );
  XNOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n568), .A2(n544), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(KEYINPUT117), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n558), .A2(n570), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(KEYINPUT118), .ZN(n549) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n552) );
  NAND2_X1 U616 ( .A1(n558), .A2(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n554) );
  XOR2_X1 U618 ( .A(G148GAT), .B(KEYINPUT52), .Z(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U620 ( .A1(n558), .A2(n576), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  XOR2_X1 U623 ( .A(G162GAT), .B(KEYINPUT121), .Z(n560) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n570), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n561), .A2(n576), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT124), .ZN(n566) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(n566), .Z(n572) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(KEYINPUT123), .B(n569), .ZN(n582) );
  INV_X1 U636 ( .A(n582), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n577), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U640 ( .A1(n577), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n581) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n585) );
  NOR2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U649 ( .A(n585), .B(n584), .Z(G1355GAT) );
endmodule

