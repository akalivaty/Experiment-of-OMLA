

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U556 ( .A(n713), .ZN(n733) );
  AND2_X1 U557 ( .A1(n679), .A2(n678), .ZN(n795) );
  BUF_X1 U558 ( .A(n681), .Z(n560) );
  AND2_X1 U559 ( .A1(G101), .A2(G2104), .ZN(n536) );
  XOR2_X1 U560 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  XNOR2_X1 U561 ( .A(n538), .B(n537), .ZN(n539) );
  NOR2_X1 U562 ( .A1(n709), .A2(n708), .ZN(n710) );
  INV_X1 U563 ( .A(KEYINPUT96), .ZN(n730) );
  INV_X1 U564 ( .A(KEYINPUT23), .ZN(n537) );
  NOR2_X1 U565 ( .A1(n526), .A2(n639), .ZN(n527) );
  NOR2_X1 U566 ( .A1(n639), .A2(G651), .ZN(n522) );
  BUF_X1 U567 ( .A(n522), .Z(n646) );
  NAND2_X1 U568 ( .A1(G47), .A2(n646), .ZN(n525) );
  INV_X1 U569 ( .A(G651), .ZN(n526) );
  NOR2_X1 U570 ( .A1(G543), .A2(n526), .ZN(n523) );
  XOR2_X2 U571 ( .A(KEYINPUT1), .B(n523), .Z(n647) );
  NAND2_X1 U572 ( .A1(G60), .A2(n647), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n531) );
  NOR2_X2 U574 ( .A1(G543), .A2(G651), .ZN(n642) );
  NAND2_X1 U575 ( .A1(G85), .A2(n642), .ZN(n529) );
  XNOR2_X2 U576 ( .A(KEYINPUT66), .B(n527), .ZN(n643) );
  NAND2_X1 U577 ( .A1(G72), .A2(n643), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U579 ( .A1(n531), .A2(n530), .ZN(G290) );
  NOR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT17), .B(n532), .Z(n681) );
  NAND2_X1 U582 ( .A1(n681), .A2(G137), .ZN(n534) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n902) );
  NAND2_X1 U584 ( .A1(n902), .A2(G113), .ZN(n533) );
  AND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n678) );
  INV_X1 U586 ( .A(G2105), .ZN(n535) );
  NOR2_X4 U587 ( .A1(n535), .A2(G2104), .ZN(n901) );
  NAND2_X1 U588 ( .A1(n901), .A2(G125), .ZN(n540) );
  INV_X1 U589 ( .A(G2105), .ZN(n561) );
  NAND2_X1 U590 ( .A1(n536), .A2(n561), .ZN(n538) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n541), .B(KEYINPUT65), .ZN(n677) );
  AND2_X1 U593 ( .A1(n678), .A2(n677), .ZN(G160) );
  NAND2_X1 U594 ( .A1(G52), .A2(n646), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G64), .A2(n647), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G90), .A2(n642), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G77), .A2(n643), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  NAND2_X1 U604 ( .A1(G51), .A2(n646), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G63), .A2(n647), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U607 ( .A(KEYINPUT6), .B(n551), .ZN(n557) );
  NAND2_X1 U608 ( .A1(n642), .A2(G89), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G76), .A2(n643), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U612 ( .A(n555), .B(KEYINPUT5), .Z(n556) );
  NOR2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U614 ( .A(KEYINPUT7), .B(n558), .Z(n559) );
  XOR2_X1 U615 ( .A(KEYINPUT73), .B(n559), .Z(G168) );
  XOR2_X1 U616 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U617 ( .A1(G138), .A2(n560), .ZN(n566) );
  AND2_X1 U618 ( .A1(n561), .A2(G2104), .ZN(n905) );
  NAND2_X1 U619 ( .A1(G102), .A2(n905), .ZN(n565) );
  NAND2_X1 U620 ( .A1(G126), .A2(n901), .ZN(n563) );
  NAND2_X1 U621 ( .A1(G114), .A2(n902), .ZN(n562) );
  AND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n682) );
  NOR2_X1 U624 ( .A1(n566), .A2(n682), .ZN(G164) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT10), .ZN(n568) );
  XNOR2_X1 U627 ( .A(KEYINPUT68), .B(n568), .ZN(G223) );
  INV_X1 U628 ( .A(G223), .ZN(n840) );
  NAND2_X1 U629 ( .A1(n840), .A2(G567), .ZN(n569) );
  XNOR2_X1 U630 ( .A(n569), .B(KEYINPUT69), .ZN(n570) );
  XNOR2_X1 U631 ( .A(KEYINPUT11), .B(n570), .ZN(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n647), .ZN(n571) );
  XNOR2_X1 U633 ( .A(n571), .B(KEYINPUT14), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G43), .A2(n646), .ZN(n572) );
  XNOR2_X1 U635 ( .A(n572), .B(KEYINPUT70), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n642), .A2(G81), .ZN(n575) );
  XNOR2_X1 U638 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U639 ( .A1(G68), .A2(n643), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT13), .B(n578), .Z(n579) );
  NOR2_X1 U642 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X2 U643 ( .A(KEYINPUT71), .B(n581), .ZN(n949) );
  INV_X1 U644 ( .A(n949), .ZN(n703) );
  NAND2_X1 U645 ( .A1(n703), .A2(G860), .ZN(G153) );
  INV_X1 U646 ( .A(G171), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G92), .A2(n642), .ZN(n583) );
  NAND2_X1 U648 ( .A1(G79), .A2(n643), .ZN(n582) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G54), .A2(n646), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G66), .A2(n647), .ZN(n584) );
  NAND2_X1 U652 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n588), .B(KEYINPUT15), .ZN(n942) );
  INV_X1 U655 ( .A(G868), .ZN(n661) );
  NAND2_X1 U656 ( .A1(n942), .A2(n661), .ZN(n589) );
  XNOR2_X1 U657 ( .A(n589), .B(KEYINPUT72), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U660 ( .A1(G53), .A2(n646), .ZN(n593) );
  NAND2_X1 U661 ( .A1(G65), .A2(n647), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G91), .A2(n642), .ZN(n594) );
  XNOR2_X1 U664 ( .A(KEYINPUT67), .B(n594), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G78), .A2(n643), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(G299) );
  NOR2_X1 U668 ( .A1(G286), .A2(n661), .ZN(n600) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U670 ( .A1(n600), .A2(n599), .ZN(G297) );
  INV_X1 U671 ( .A(G559), .ZN(n605) );
  NOR2_X1 U672 ( .A1(G860), .A2(n605), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n942), .A2(n601), .ZN(n604) );
  XNOR2_X1 U674 ( .A(KEYINPUT16), .B(KEYINPUT74), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT75), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(G148) );
  INV_X1 U677 ( .A(n942), .ZN(n658) );
  NAND2_X1 U678 ( .A1(n605), .A2(n658), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n606), .A2(G868), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n949), .A2(n661), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U682 ( .A1(G123), .A2(n901), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n905), .A2(G99), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U686 ( .A1(G135), .A2(n560), .ZN(n613) );
  NAND2_X1 U687 ( .A1(G111), .A2(n902), .ZN(n612) );
  NAND2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n615), .A2(n614), .ZN(n1014) );
  XNOR2_X1 U690 ( .A(n1014), .B(G2096), .ZN(n616) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT76), .ZN(n618) );
  INV_X1 U692 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U694 ( .A1(n646), .A2(G50), .ZN(n619) );
  XNOR2_X1 U695 ( .A(KEYINPUT81), .B(n619), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n647), .A2(G62), .ZN(n620) );
  XOR2_X1 U697 ( .A(KEYINPUT80), .B(n620), .Z(n621) );
  NOR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U699 ( .A(KEYINPUT82), .B(n623), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n643), .A2(G75), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G88), .A2(n642), .ZN(n624) );
  AND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(G303) );
  INV_X1 U704 ( .A(G303), .ZN(G166) );
  NAND2_X1 U705 ( .A1(G48), .A2(n646), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G61), .A2(n647), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n643), .A2(G73), .ZN(n630) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  NOR2_X1 U710 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n642), .A2(G86), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G49), .A2(n646), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U716 ( .A1(n647), .A2(n637), .ZN(n638) );
  XOR2_X1 U717 ( .A(KEYINPUT79), .B(n638), .Z(n641) );
  NAND2_X1 U718 ( .A1(n639), .A2(G87), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(G288) );
  INV_X1 U720 ( .A(G299), .ZN(n718) );
  XNOR2_X1 U721 ( .A(n718), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U722 ( .A(G166), .B(G305), .ZN(n653) );
  NAND2_X1 U723 ( .A1(G93), .A2(n642), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G80), .A2(n643), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G55), .A2(n646), .ZN(n649) );
  NAND2_X1 U727 ( .A1(G67), .A2(n647), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U730 ( .A(n652), .B(KEYINPUT78), .Z(n846) );
  XOR2_X1 U731 ( .A(n653), .B(n846), .Z(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(G288), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U734 ( .A(n657), .B(n656), .ZN(n915) );
  NAND2_X1 U735 ( .A1(G559), .A2(n658), .ZN(n659) );
  XOR2_X1 U736 ( .A(n949), .B(n659), .Z(n844) );
  XOR2_X1 U737 ( .A(n915), .B(n844), .Z(n660) );
  NOR2_X1 U738 ( .A1(n661), .A2(n660), .ZN(n663) );
  NOR2_X1 U739 ( .A1(n846), .A2(G868), .ZN(n662) );
  NOR2_X1 U740 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n664) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n665), .ZN(n666) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n667), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U747 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n669) );
  NAND2_X1 U748 ( .A1(G132), .A2(G82), .ZN(n668) );
  XNOR2_X1 U749 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U750 ( .A1(n670), .A2(G218), .ZN(n671) );
  NAND2_X1 U751 ( .A1(G96), .A2(n671), .ZN(n848) );
  NAND2_X1 U752 ( .A1(n848), .A2(G2106), .ZN(n675) );
  NAND2_X1 U753 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U754 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U755 ( .A1(G108), .A2(n673), .ZN(n849) );
  NAND2_X1 U756 ( .A1(n849), .A2(G567), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n675), .A2(n674), .ZN(n850) );
  NAND2_X1 U758 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U759 ( .A1(n850), .A2(n676), .ZN(n843) );
  NAND2_X1 U760 ( .A1(n843), .A2(G36), .ZN(G176) );
  AND2_X1 U761 ( .A1(G40), .A2(n677), .ZN(n679) );
  INV_X1 U762 ( .A(G1384), .ZN(n683) );
  AND2_X1 U763 ( .A1(G138), .A2(n683), .ZN(n680) );
  AND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n685) );
  AND2_X1 U765 ( .A1(n683), .A2(n682), .ZN(n684) );
  OR2_X1 U766 ( .A1(n685), .A2(n684), .ZN(n796) );
  NAND2_X1 U767 ( .A1(n795), .A2(n796), .ZN(n686) );
  XNOR2_X1 U768 ( .A(n686), .B(KEYINPUT64), .ZN(n687) );
  INV_X2 U769 ( .A(n687), .ZN(n713) );
  NOR2_X1 U770 ( .A1(n733), .A2(G2084), .ZN(n745) );
  NAND2_X1 U771 ( .A1(n733), .A2(G8), .ZN(n779) );
  NOR2_X1 U772 ( .A1(G1966), .A2(n779), .ZN(n747) );
  NOR2_X1 U773 ( .A1(n745), .A2(n747), .ZN(n688) );
  NAND2_X1 U774 ( .A1(G8), .A2(n688), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT30), .B(n689), .ZN(n690) );
  NOR2_X1 U776 ( .A1(G168), .A2(n690), .ZN(n694) );
  XNOR2_X1 U777 ( .A(KEYINPUT25), .B(G2078), .ZN(n995) );
  NAND2_X1 U778 ( .A1(n713), .A2(n995), .ZN(n692) );
  XNOR2_X1 U779 ( .A(G1961), .B(KEYINPUT91), .ZN(n972) );
  NAND2_X1 U780 ( .A1(n733), .A2(n972), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n725) );
  NOR2_X1 U782 ( .A1(G171), .A2(n725), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U784 ( .A(n695), .B(KEYINPUT31), .ZN(n729) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n713), .ZN(n696) );
  XNOR2_X1 U786 ( .A(n696), .B(KEYINPUT26), .ZN(n698) );
  NAND2_X1 U787 ( .A1(G1341), .A2(n733), .ZN(n697) );
  NAND2_X1 U788 ( .A1(n698), .A2(n697), .ZN(n700) );
  INV_X1 U789 ( .A(KEYINPUT93), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n700), .B(n699), .ZN(n706) );
  NAND2_X1 U791 ( .A1(G2067), .A2(n713), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n733), .A2(G1348), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n707) );
  NAND2_X1 U794 ( .A1(n707), .A2(n942), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U796 ( .A1(n706), .A2(n705), .ZN(n709) );
  NOR2_X1 U797 ( .A1(n707), .A2(n942), .ZN(n708) );
  XNOR2_X1 U798 ( .A(n710), .B(KEYINPUT94), .ZN(n717) );
  NAND2_X1 U799 ( .A1(n713), .A2(G2072), .ZN(n712) );
  XNOR2_X1 U800 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n711) );
  XNOR2_X1 U801 ( .A(n712), .B(n711), .ZN(n715) );
  INV_X1 U802 ( .A(G1956), .ZN(n962) );
  NOR2_X1 U803 ( .A1(n713), .A2(n962), .ZN(n714) );
  NOR2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n722) );
  NOR2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U808 ( .A(n720), .B(KEYINPUT28), .Z(n721) );
  NAND2_X1 U809 ( .A1(n722), .A2(n721), .ZN(n724) );
  XOR2_X1 U810 ( .A(KEYINPUT95), .B(KEYINPUT29), .Z(n723) );
  XNOR2_X1 U811 ( .A(n724), .B(n723), .ZN(n727) );
  AND2_X1 U812 ( .A1(n725), .A2(G171), .ZN(n726) );
  NOR2_X1 U813 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X2 U814 ( .A1(n729), .A2(n728), .ZN(n731) );
  XNOR2_X1 U815 ( .A(n731), .B(n730), .ZN(n746) );
  AND2_X1 U816 ( .A1(G286), .A2(G8), .ZN(n732) );
  NAND2_X1 U817 ( .A1(n746), .A2(n732), .ZN(n740) );
  INV_X1 U818 ( .A(G8), .ZN(n738) );
  NOR2_X1 U819 ( .A1(n733), .A2(G2090), .ZN(n735) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n779), .ZN(n734) );
  NOR2_X1 U821 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U822 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U823 ( .A1(n738), .A2(n737), .ZN(n739) );
  AND2_X1 U824 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X2 U825 ( .A(n741), .B(KEYINPUT32), .ZN(n769) );
  INV_X1 U826 ( .A(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n954) );
  INV_X1 U828 ( .A(n779), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n954), .A2(n742), .ZN(n743) );
  AND2_X1 U830 ( .A1(n754), .A2(n743), .ZN(n756) );
  INV_X1 U831 ( .A(n756), .ZN(n744) );
  AND2_X1 U832 ( .A1(n769), .A2(n744), .ZN(n752) );
  NAND2_X1 U833 ( .A1(G8), .A2(n745), .ZN(n751) );
  INV_X1 U834 ( .A(n746), .ZN(n748) );
  NOR2_X2 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U836 ( .A(KEYINPUT97), .B(n749), .Z(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n770) );
  NAND2_X1 U838 ( .A1(n752), .A2(n770), .ZN(n758) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U841 ( .A1(n760), .A2(n753), .ZN(n944) );
  AND2_X1 U842 ( .A1(n944), .A2(n754), .ZN(n755) );
  OR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U845 ( .A(n759), .B(KEYINPUT98), .ZN(n765) );
  NAND2_X1 U846 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  NOR2_X1 U847 ( .A1(n779), .A2(n761), .ZN(n763) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n937) );
  INV_X1 U849 ( .A(n937), .ZN(n762) );
  NOR2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n775) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n766) );
  XOR2_X1 U853 ( .A(KEYINPUT99), .B(n766), .Z(n767) );
  NAND2_X1 U854 ( .A1(G8), .A2(n767), .ZN(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT100), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U858 ( .A1(n773), .A2(n779), .ZN(n774) );
  NAND2_X1 U859 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U860 ( .A(n776), .B(KEYINPUT101), .ZN(n782) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XOR2_X1 U862 ( .A(n777), .B(KEYINPUT24), .Z(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U864 ( .A(KEYINPUT90), .B(n780), .Z(n781) );
  NAND2_X1 U865 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U866 ( .A(n783), .B(KEYINPUT102), .ZN(n822) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n833) );
  NAND2_X1 U868 ( .A1(n560), .A2(G140), .ZN(n784) );
  XOR2_X1 U869 ( .A(KEYINPUT85), .B(n784), .Z(n786) );
  NAND2_X1 U870 ( .A1(n905), .A2(G104), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U872 ( .A(KEYINPUT34), .B(n787), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G128), .A2(n901), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G116), .A2(n902), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U876 ( .A(KEYINPUT35), .B(n790), .Z(n791) );
  XNOR2_X1 U877 ( .A(KEYINPUT86), .B(n791), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(n794) );
  XNOR2_X1 U879 ( .A(KEYINPUT36), .B(n794), .ZN(n879) );
  NOR2_X1 U880 ( .A1(n833), .A2(n879), .ZN(n1034) );
  INV_X1 U881 ( .A(n795), .ZN(n797) );
  NOR2_X1 U882 ( .A1(n797), .A2(n796), .ZN(n836) );
  NAND2_X1 U883 ( .A1(n1034), .A2(n836), .ZN(n830) );
  NAND2_X1 U884 ( .A1(G95), .A2(n905), .ZN(n799) );
  NAND2_X1 U885 ( .A1(G119), .A2(n901), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U887 ( .A1(G131), .A2(n560), .ZN(n800) );
  XNOR2_X1 U888 ( .A(KEYINPUT87), .B(n800), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n902), .A2(G107), .ZN(n803) );
  NAND2_X1 U891 ( .A1(n804), .A2(n803), .ZN(n885) );
  NAND2_X1 U892 ( .A1(G1991), .A2(n885), .ZN(n805) );
  XOR2_X1 U893 ( .A(KEYINPUT88), .B(n805), .Z(n815) );
  NAND2_X1 U894 ( .A1(n902), .A2(G117), .ZN(n812) );
  NAND2_X1 U895 ( .A1(G129), .A2(n901), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G141), .A2(n560), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n810) );
  NAND2_X1 U898 ( .A1(n905), .A2(G105), .ZN(n808) );
  XOR2_X1 U899 ( .A(KEYINPUT38), .B(n808), .Z(n809) );
  NOR2_X1 U900 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U901 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U902 ( .A(KEYINPUT89), .B(n813), .Z(n878) );
  AND2_X1 U903 ( .A1(n878), .A2(G1996), .ZN(n814) );
  NOR2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n1022) );
  INV_X1 U905 ( .A(n836), .ZN(n816) );
  NOR2_X1 U906 ( .A1(n1022), .A2(n816), .ZN(n825) );
  INV_X1 U907 ( .A(n825), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n830), .A2(n817), .ZN(n820) );
  XNOR2_X1 U909 ( .A(G1986), .B(G290), .ZN(n957) );
  NAND2_X1 U910 ( .A1(n957), .A2(n836), .ZN(n818) );
  XOR2_X1 U911 ( .A(KEYINPUT84), .B(n818), .Z(n819) );
  NOR2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n838) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n878), .ZN(n1012) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n885), .ZN(n1015) );
  NOR2_X1 U917 ( .A1(n823), .A2(n1015), .ZN(n824) );
  NOR2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U919 ( .A(KEYINPUT103), .B(n826), .Z(n827) );
  NOR2_X1 U920 ( .A1(n1012), .A2(n827), .ZN(n828) );
  XNOR2_X1 U921 ( .A(KEYINPUT104), .B(n828), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT39), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U924 ( .A(KEYINPUT105), .B(n832), .Z(n834) );
  NAND2_X1 U925 ( .A1(n833), .A2(n879), .ZN(n1031) );
  NAND2_X1 U926 ( .A1(n834), .A2(n1031), .ZN(n835) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U928 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U929 ( .A(n839), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U932 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U934 ( .A1(n843), .A2(n842), .ZN(G188) );
  XNOR2_X1 U936 ( .A(KEYINPUT77), .B(n844), .ZN(n845) );
  NOR2_X1 U937 ( .A1(G860), .A2(n845), .ZN(n847) );
  XOR2_X1 U938 ( .A(n847), .B(n846), .Z(G145) );
  INV_X1 U939 ( .A(G132), .ZN(G219) );
  INV_X1 U940 ( .A(G120), .ZN(G236) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  INV_X1 U942 ( .A(G82), .ZN(G220) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n849), .A2(n848), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  INV_X1 U946 ( .A(n850), .ZN(G319) );
  XNOR2_X1 U947 ( .A(G1996), .B(G2474), .ZN(n860) );
  XOR2_X1 U948 ( .A(G1986), .B(G1991), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1956), .B(G1961), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U951 ( .A(G1976), .B(G1981), .Z(n854) );
  XNOR2_X1 U952 ( .A(G1966), .B(G1971), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U954 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U955 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n860), .B(n859), .ZN(G229) );
  XOR2_X1 U958 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n862) );
  XNOR2_X1 U959 ( .A(G2678), .B(KEYINPUT43), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2090), .Z(n864) );
  XNOR2_X1 U962 ( .A(G2072), .B(G2067), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U964 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U965 ( .A(G2096), .B(G2100), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n870) );
  XOR2_X1 U967 ( .A(G2084), .B(G2078), .Z(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(G227) );
  NAND2_X1 U969 ( .A1(G124), .A2(n901), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n871), .B(KEYINPUT44), .ZN(n873) );
  NAND2_X1 U971 ( .A1(n905), .A2(G100), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n877) );
  NAND2_X1 U973 ( .A1(G136), .A2(n560), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G112), .A2(n902), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U976 ( .A1(n877), .A2(n876), .ZN(G162) );
  XNOR2_X1 U977 ( .A(G162), .B(n1014), .ZN(n881) );
  XOR2_X1 U978 ( .A(n879), .B(n878), .Z(n880) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(n889) );
  XOR2_X1 U980 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n883) );
  XNOR2_X1 U981 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(KEYINPUT116), .B(n884), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n885), .B(KEYINPUT48), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U986 ( .A(n889), .B(n888), .Z(n900) );
  NAND2_X1 U987 ( .A1(n901), .A2(G127), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n890), .B(KEYINPUT114), .ZN(n892) );
  NAND2_X1 U989 ( .A1(G115), .A2(n902), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n893), .B(KEYINPUT47), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G139), .A2(n560), .ZN(n894) );
  NAND2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n898) );
  NAND2_X1 U994 ( .A1(G103), .A2(n905), .ZN(n896) );
  XNOR2_X1 U995 ( .A(KEYINPUT113), .B(n896), .ZN(n897) );
  NOR2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n1023) );
  XNOR2_X1 U997 ( .A(G164), .B(n1023), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n913) );
  NAND2_X1 U999 ( .A1(G130), .A2(n901), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G118), .A2(n902), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(G106), .A2(n905), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n560), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(KEYINPUT45), .B(n908), .Z(n909) );
  NOR2_X1 U1006 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1007 ( .A(G160), .B(n911), .Z(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n914), .ZN(G395) );
  XNOR2_X1 U1010 ( .A(G286), .B(n915), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n942), .B(G171), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(n918), .B(n949), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n919), .ZN(G397) );
  XNOR2_X1 U1015 ( .A(G2451), .B(G2427), .ZN(n929) );
  XOR2_X1 U1016 ( .A(KEYINPUT107), .B(G2443), .Z(n921) );
  XNOR2_X1 U1017 ( .A(G2435), .B(G2438), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n921), .B(n920), .ZN(n925) );
  XOR2_X1 U1019 ( .A(G2454), .B(G2430), .Z(n923) );
  XNOR2_X1 U1020 ( .A(G1348), .B(G1341), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  XOR2_X1 U1022 ( .A(n925), .B(n924), .Z(n927) );
  XNOR2_X1 U1023 ( .A(G2446), .B(KEYINPUT106), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(n927), .B(n926), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(n929), .B(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n930), .A2(G14), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(G319), .A2(n936), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(G229), .A2(G227), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(KEYINPUT49), .B(n931), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1033 ( .A(G225), .ZN(G308) );
  INV_X1 U1034 ( .A(G108), .ZN(G238) );
  INV_X1 U1035 ( .A(n936), .ZN(G401) );
  XNOR2_X1 U1036 ( .A(KEYINPUT56), .B(G16), .ZN(n961) );
  XNOR2_X1 U1037 ( .A(G1966), .B(G168), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(n939), .B(KEYINPUT57), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT124), .B(n940), .ZN(n948) );
  XOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT125), .Z(n941) );
  XNOR2_X1 U1042 ( .A(n942), .B(n941), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(G1971), .A2(G303), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G1341), .B(n949), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G299), .B(G1956), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(G301), .B(G1961), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n1044) );
  XNOR2_X1 U1056 ( .A(G20), .B(n962), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(G1341), .B(G19), .ZN(n964) );
  XNOR2_X1 U1058 ( .A(G6), .B(G1981), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1061 ( .A(KEYINPUT59), .B(G1348), .Z(n967) );
  XNOR2_X1 U1062 ( .A(G4), .B(n967), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT60), .B(n970), .ZN(n981) );
  XOR2_X1 U1065 ( .A(KEYINPUT126), .B(G5), .Z(n971) );
  XNOR2_X1 U1066 ( .A(n972), .B(n971), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G22), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G24), .B(G1986), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1070 ( .A(G1976), .B(G23), .Z(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(KEYINPUT58), .B(n977), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G21), .B(G1966), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n984), .Z(n985) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n985), .ZN(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT127), .B(n986), .Z(n1042) );
  XOR2_X1 U1080 ( .A(G2090), .B(G35), .Z(n1002) );
  XNOR2_X1 U1081 ( .A(G2072), .B(G33), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G1991), .B(G25), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n994) );
  XOR2_X1 U1084 ( .A(G2067), .B(G26), .Z(n989) );
  NAND2_X1 U1085 ( .A1(n989), .A2(G28), .ZN(n992) );
  XNOR2_X1 U1086 ( .A(KEYINPUT120), .B(G1996), .ZN(n990) );
  XNOR2_X1 U1087 ( .A(G32), .B(n990), .ZN(n991) );
  NOR2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n997) );
  XOR2_X1 U1090 ( .A(G27), .B(n995), .Z(n996) );
  NOR2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1092 ( .A(n998), .B(KEYINPUT122), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(n999), .B(KEYINPUT121), .ZN(n1000) );
  XNOR2_X1 U1094 ( .A(n1000), .B(KEYINPUT53), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(G34), .B(G2084), .ZN(n1003) );
  XNOR2_X1 U1097 ( .A(KEYINPUT54), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1099 ( .A(KEYINPUT55), .B(n1006), .ZN(n1008) );
  INV_X1 U1100 ( .A(G29), .ZN(n1007) );
  NAND2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1009), .A2(G11), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(KEYINPUT123), .B(n1010), .ZN(n1040) );
  XOR2_X1 U1104 ( .A(G2090), .B(G162), .Z(n1011) );
  NOR2_X1 U1105 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1106 ( .A(KEYINPUT51), .B(n1013), .Z(n1018) );
  NOR2_X1 U1107 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1108 ( .A(KEYINPUT117), .B(n1016), .Z(n1017) );
  NAND2_X1 U1109 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1110 ( .A(G160), .B(G2084), .Z(n1019) );
  NOR2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1030) );
  XNOR2_X1 U1113 ( .A(G164), .B(G2078), .ZN(n1026) );
  XNOR2_X1 U1114 ( .A(G2072), .B(n1023), .ZN(n1024) );
  XNOR2_X1 U1115 ( .A(n1024), .B(KEYINPUT118), .ZN(n1025) );
  NAND2_X1 U1116 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1117 ( .A(n1027), .B(KEYINPUT119), .ZN(n1028) );
  XOR2_X1 U1118 ( .A(KEYINPUT50), .B(n1028), .Z(n1029) );
  NOR2_X1 U1119 ( .A1(n1030), .A2(n1029), .ZN(n1032) );
  NAND2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1122 ( .A(KEYINPUT52), .B(n1035), .ZN(n1037) );
  INV_X1 U1123 ( .A(KEYINPUT55), .ZN(n1036) );
  NAND2_X1 U1124 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NAND2_X1 U1125 ( .A1(n1038), .A2(G29), .ZN(n1039) );
  NAND2_X1 U1126 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  NOR2_X1 U1127 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1128 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XOR2_X1 U1129 ( .A(KEYINPUT62), .B(n1045), .Z(G311) );
  INV_X1 U1130 ( .A(G311), .ZN(G150) );
endmodule

