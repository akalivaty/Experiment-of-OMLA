//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT79), .Z(new_n189));
  OAI21_X1  g003(.A(G214), .B1(G237), .B2(G902), .ZN(new_n190));
  XOR2_X1   g004(.A(G110), .B(G122), .Z(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G116), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(KEYINPUT5), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G113), .B1(new_n194), .B2(KEYINPUT5), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n194), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT2), .B(G113), .ZN(new_n199));
  OAI22_X1  g013(.A1(new_n196), .A2(new_n197), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT85), .B1(new_n202), .B2(G104), .ZN(new_n203));
  INV_X1    g017(.A(G104), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(KEYINPUT85), .A3(G104), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n201), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT82), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n202), .B2(G104), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(KEYINPUT82), .A3(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(KEYINPUT81), .A3(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT3), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(new_n202), .A3(KEYINPUT81), .A4(G104), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n201), .A4(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT84), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(new_n218), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n208), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT86), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n214), .A2(new_n216), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n224), .A2(KEYINPUT84), .A3(new_n201), .A4(new_n212), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n218), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n207), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT86), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n200), .B1(new_n223), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n226), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT83), .A4(new_n216), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(G101), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(KEYINPUT4), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n198), .B(new_n199), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n238), .A3(G101), .A4(new_n234), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n191), .B1(new_n229), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n200), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT86), .B1(new_n230), .B2(new_n208), .ZN(new_n243));
  AOI211_X1 g057(.A(new_n222), .B(new_n207), .C1(new_n225), .C2(new_n226), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n246));
  INV_X1    g060(.A(new_n191), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n248), .A3(KEYINPUT6), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n250), .B(new_n191), .C1(new_n229), .C2(new_n240), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT65), .B1(new_n257), .B2(G146), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(G146), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n254), .B(new_n256), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n252), .B1(new_n253), .B2(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n253), .A2(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n265), .A2(KEYINPUT66), .A3(new_n254), .A4(new_n256), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n255), .B(KEYINPUT64), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n257), .A2(G146), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n262), .A2(new_n266), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n264), .A2(new_n269), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT68), .B(KEYINPUT1), .C1(new_n257), .C2(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G128), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT68), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G125), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n265), .A2(new_n280), .A3(G128), .A4(new_n254), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G224), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G953), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT89), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n283), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n249), .A2(new_n251), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n273), .A2(new_n282), .A3(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT91), .ZN(new_n292));
  AOI22_X1  g106(.A1(KEYINPUT90), .A2(new_n282), .B1(new_n272), .B2(G125), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n282), .A2(KEYINPUT90), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n191), .B(KEYINPUT8), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n221), .A2(new_n200), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n227), .A2(new_n242), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n292), .A2(new_n295), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n300), .B2(new_n248), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n288), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n288), .B2(new_n301), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n190), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G469), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  INV_X1    g122(.A(G953), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G227), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT80), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G140), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n262), .A2(new_n266), .A3(new_n271), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n236), .A2(new_n314), .A3(new_n239), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n265), .A2(new_n254), .ZN(new_n316));
  INV_X1    g130(.A(G128), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n317), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n281), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n230), .A2(new_n208), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT10), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n278), .A2(new_n281), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT10), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n243), .B2(new_n244), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(KEYINPUT87), .B(new_n326), .C1(new_n243), .C2(new_n244), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n323), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G137), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(KEYINPUT11), .A3(G134), .ZN(new_n333));
  INV_X1    g147(.A(G134), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G137), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT11), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n337), .B1(new_n334), .B2(G137), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G131), .ZN(new_n340));
  INV_X1    g154(.A(G131), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n338), .A2(new_n333), .A3(new_n341), .A4(new_n335), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT67), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n313), .B1(new_n331), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n324), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n221), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n347), .B1(new_n350), .B2(new_n320), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(KEYINPUT12), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n313), .ZN(new_n354));
  INV_X1    g168(.A(new_n323), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n223), .A2(new_n228), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT87), .B1(new_n356), .B2(new_n326), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n328), .B(new_n325), .C1(new_n223), .C2(new_n228), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n346), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n355), .B(new_n347), .C1(new_n357), .C2(new_n358), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n354), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n362), .B2(KEYINPUT88), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n329), .A2(new_n330), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n347), .B1(new_n364), .B2(new_n355), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n346), .B(new_n323), .C1(new_n329), .C2(new_n330), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT88), .B(new_n313), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n307), .B(new_n308), .C1(new_n363), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n361), .A2(new_n352), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n313), .A2(new_n370), .B1(new_n348), .B2(new_n360), .ZN(new_n371));
  OAI21_X1  g185(.A(G469), .B1(new_n371), .B2(G902), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n189), .B(new_n306), .C1(new_n369), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n332), .A2(G134), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n341), .B1(new_n374), .B2(new_n335), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n278), .B2(new_n281), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n342), .B(new_n343), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n346), .A2(new_n314), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT70), .B1(new_n378), .B2(KEYINPUT30), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n377), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT69), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT69), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n346), .A2(new_n314), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n382), .A2(KEYINPUT30), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n384), .A2(new_n383), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n387), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n382), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n388), .A3(new_n237), .ZN(new_n389));
  INV_X1    g203(.A(new_n237), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n382), .A2(new_n390), .A3(new_n383), .A4(new_n384), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT26), .B(G101), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n309), .A3(G210), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n392), .B(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n396));
  XNOR2_X1  g210(.A(new_n395), .B(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n389), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT28), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n384), .A2(new_n380), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n399), .B1(new_n400), .B2(new_n237), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n237), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n401), .B(new_n402), .C1(new_n399), .C2(new_n391), .ZN(new_n403));
  INV_X1    g217(.A(new_n397), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n398), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n384), .A2(new_n383), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT69), .B1(new_n376), .B2(new_n377), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n237), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n391), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT28), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n401), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(KEYINPUT29), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n308), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G472), .B1(new_n406), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT73), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT73), .B(G472), .C1(new_n406), .C2(new_n414), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n389), .A2(new_n391), .A3(new_n404), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT31), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n403), .A2(new_n397), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT31), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n389), .A2(new_n423), .A3(new_n391), .A4(new_n404), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G472), .A2(G902), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(KEYINPUT32), .B1(new_n427), .B2(KEYINPUT72), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT72), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT32), .ZN(new_n430));
  AOI211_X1 g244(.A(new_n429), .B(new_n430), .C1(new_n425), .C2(new_n426), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n419), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G217), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(G234), .B2(new_n308), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT25), .ZN(new_n436));
  INV_X1    g250(.A(G110), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n317), .A2(G119), .ZN(new_n438));
  OR2_X1    g252(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n192), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI211_X1 g256(.A(KEYINPUT23), .B(new_n438), .C1(new_n442), .C2(KEYINPUT75), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT75), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n442), .A2(new_n444), .B1(G119), .B2(new_n317), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n437), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT76), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g262(.A(KEYINPUT76), .B(new_n437), .C1(new_n443), .C2(new_n445), .ZN(new_n449));
  XOR2_X1   g263(.A(KEYINPUT24), .B(G110), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n438), .A2(new_n440), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G125), .B(G140), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT16), .ZN(new_n456));
  OR3_X1    g270(.A1(new_n279), .A2(KEYINPUT16), .A3(G140), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(G146), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n253), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n458), .ZN(new_n461));
  AOI21_X1  g275(.A(G146), .B1(new_n456), .B2(new_n457), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n461), .A2(new_n462), .B1(new_n452), .B2(new_n451), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n443), .A2(new_n437), .A3(new_n445), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n467));
  NAND3_X1  g281(.A1(new_n309), .A2(G221), .A3(G234), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT22), .B(G137), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n471), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n458), .A2(new_n459), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n446), .A2(new_n447), .B1(new_n452), .B2(new_n451), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n475), .B2(new_n449), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n473), .B1(new_n476), .B2(new_n465), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n436), .B1(new_n479), .B2(G902), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(KEYINPUT25), .A3(new_n308), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n435), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n434), .A2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n461), .A2(new_n462), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n393), .A2(new_n309), .A3(G214), .ZN(new_n488));
  OR2_X1    g302(.A1(KEYINPUT92), .A2(G143), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(new_n341), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT17), .ZN(new_n492));
  NOR2_X1   g306(.A1(KEYINPUT92), .A2(G143), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n488), .B(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G131), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n341), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n487), .B(new_n492), .C1(new_n497), .C2(KEYINPUT17), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(KEYINPUT18), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n490), .B1(new_n500), .B2(new_n341), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n455), .B(new_n253), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(G113), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n204), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n498), .A2(new_n503), .A3(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n308), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G475), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n507), .B1(new_n498), .B2(new_n503), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n455), .B(KEYINPUT19), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n253), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n497), .A2(new_n458), .A3(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n503), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n521), .ZN(new_n523));
  NOR4_X1   g337(.A1(new_n515), .A2(new_n519), .A3(KEYINPUT20), .A4(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n513), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(KEYINPUT94), .B(new_n513), .C1(new_n522), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(KEYINPUT96), .A2(G952), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(KEYINPUT96), .A2(G952), .ZN(new_n532));
  AOI21_X1  g346(.A(G953), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G234), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n393), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(KEYINPUT21), .B(G898), .Z(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI211_X1 g352(.A(new_n308), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT95), .ZN(new_n541));
  XNOR2_X1  g355(.A(G116), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n202), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n317), .A2(G143), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n334), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n257), .A2(G128), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n544), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n548), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n542), .B(G107), .ZN(new_n552));
  NAND2_X1  g366(.A1(KEYINPUT14), .A2(G107), .ZN(new_n553));
  INV_X1    g367(.A(G122), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(G116), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n548), .B(G134), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n542), .A2(KEYINPUT14), .A3(G107), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n551), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n187), .A2(new_n433), .A3(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n551), .B(new_n561), .C1(new_n556), .C2(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n308), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n568), .B1(new_n565), .B2(new_n308), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n541), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n569), .A3(KEYINPUT95), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n529), .A2(new_n540), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n373), .A2(new_n432), .A3(new_n486), .A4(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  NAND2_X1  g392(.A1(new_n370), .A2(new_n313), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n348), .A2(new_n360), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n307), .B1(new_n581), .B2(new_n308), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n361), .A2(new_n354), .A3(new_n352), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n313), .B1(new_n365), .B2(new_n366), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT88), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(G902), .B1(new_n586), .B2(new_n367), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n582), .B1(new_n587), .B2(new_n307), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n425), .A2(new_n308), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G472), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n486), .A3(new_n427), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n588), .A2(new_n189), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n565), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n562), .B2(KEYINPUT97), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n595), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(G478), .A3(new_n308), .A4(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n566), .B1(new_n593), .B2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n529), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT98), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n529), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n305), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n303), .ZN(new_n608));
  INV_X1    g422(.A(new_n540), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n190), .A3(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n592), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT99), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n612), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n306), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n520), .A2(new_n514), .A3(new_n521), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT101), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n524), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n621), .B1(new_n622), .B2(new_n522), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n540), .B1(new_n572), .B2(new_n574), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n522), .A2(new_n622), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n620), .A3(new_n618), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n623), .A2(new_n513), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT102), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n626), .A2(new_n513), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n623), .A4(new_n624), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n616), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n592), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT103), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND2_X1  g450(.A1(new_n590), .A2(new_n427), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n482), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n460), .A2(new_n466), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n640), .B(new_n641), .Z(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n483), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n639), .A2(KEYINPUT104), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n645));
  INV_X1    g459(.A(new_n643), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n645), .B1(new_n482), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n373), .A2(new_n576), .A3(new_n638), .A4(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT37), .B(G110), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G12));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n536), .B1(new_n652), .B2(new_n539), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n629), .A2(new_n623), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n575), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n373), .A2(new_n432), .A3(new_n648), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT105), .B(G128), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G30));
  AOI21_X1  g474(.A(new_n189), .B1(new_n369), .B2(new_n372), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n653), .B(KEYINPUT39), .Z(new_n662));
  AND2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n661), .A2(new_n664), .A3(new_n662), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n304), .A2(new_n305), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n429), .B1(new_n425), .B2(new_n426), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT32), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n389), .A2(new_n391), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n404), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n308), .B1(new_n410), .B2(new_n404), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n482), .A2(new_n646), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n529), .A2(new_n575), .ZN(new_n683));
  INV_X1    g497(.A(new_n190), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n666), .A2(new_n672), .A3(new_n680), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n665), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(new_n257), .ZN(G45));
  NOR2_X1   g502(.A1(new_n601), .A2(new_n653), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n373), .A2(new_n432), .A3(new_n648), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  AOI211_X1 g505(.A(G469), .B(G902), .C1(new_n586), .C2(new_n367), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n584), .A2(new_n585), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n367), .A3(new_n353), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n307), .B1(new_n694), .B2(new_n308), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n692), .A2(new_n695), .A3(new_n189), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n605), .A2(new_n610), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n432), .A3(new_n697), .A4(new_n486), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT41), .B(G113), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT107), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n698), .B(new_n700), .ZN(G15));
  NAND4_X1  g515(.A1(new_n696), .A2(new_n432), .A3(new_n486), .A4(new_n632), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  OAI21_X1  g517(.A(new_n308), .B1(new_n363), .B2(new_n368), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  INV_X1    g519(.A(new_n189), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n616), .A3(new_n706), .A4(new_n369), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AND2_X1   g522(.A1(new_n432), .A2(new_n648), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n576), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NAND2_X1  g525(.A1(new_n412), .A2(new_n397), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n421), .A2(new_n424), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n426), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n590), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n486), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n529), .A2(new_n609), .A3(new_n575), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n696), .A2(new_n616), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G122), .ZN(G24));
  NAND4_X1  g534(.A1(new_n689), .A2(new_n682), .A3(new_n590), .A4(new_n714), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n707), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n279), .ZN(G27));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n427), .B(KEYINPUT32), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n716), .B1(new_n725), .B2(new_n419), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n601), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n654), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n608), .A2(new_n684), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n661), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n724), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n661), .A2(new_n432), .A3(new_n486), .A4(new_n732), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n730), .B1(new_n735), .B2(new_n729), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n706), .B(new_n732), .C1(new_n692), .C2(new_n582), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n726), .A4(new_n731), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n734), .A2(new_n736), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G131), .ZN(G33));
  INV_X1    g555(.A(new_n657), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n735), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n334), .ZN(G36));
  INV_X1    g558(.A(new_n732), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n527), .A2(new_n528), .A3(new_n600), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n527), .A2(new_n600), .A3(KEYINPUT43), .A4(new_n528), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n637), .A2(new_n750), .A3(new_n682), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT44), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n745), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n637), .A2(new_n750), .A3(new_n682), .A4(KEYINPUT44), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT45), .B1(new_n579), .B2(new_n580), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n756), .B1(new_n757), .B2(new_n307), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT109), .B(G469), .C1(new_n371), .C2(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n371), .A2(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(G469), .A2(G902), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n369), .A3(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n755), .A2(new_n767), .A3(new_n706), .A4(new_n662), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n369), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT46), .B1(new_n761), .B2(new_n762), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n706), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT47), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n767), .A2(new_n774), .A3(new_n706), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n432), .A2(new_n745), .A3(new_n729), .A4(new_n486), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n773), .A2(new_n775), .A3(new_n779), .A4(new_n776), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n432), .A2(new_n661), .A3(new_n616), .A4(new_n648), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n722), .B1(new_n784), .B2(new_n657), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n786));
  NOR4_X1   g600(.A1(new_n682), .A2(new_n306), .A3(new_n683), .A4(new_n653), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n680), .A2(new_n787), .A3(new_n661), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(new_n786), .A3(new_n690), .A4(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n729), .A2(new_n715), .A3(new_n681), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n696), .A2(new_n790), .A3(new_n616), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n658), .A2(new_n690), .A3(new_n791), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT114), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n570), .A2(new_n571), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n655), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n432), .A2(new_n648), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n737), .B1(new_n799), .B2(new_n721), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n743), .A2(new_n800), .A3(KEYINPUT113), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n529), .A2(new_n796), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT112), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n592), .B(new_n611), .C1(new_n728), .C2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n710), .A3(new_n649), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n698), .A2(new_n702), .A3(new_n577), .A4(new_n719), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n801), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT113), .B1(new_n743), .B2(new_n800), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n740), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n795), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n794), .B1(new_n789), .B2(new_n793), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n783), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n813));
  INV_X1    g627(.A(new_n805), .ZN(new_n814));
  INV_X1    g628(.A(new_n806), .ZN(new_n815));
  INV_X1    g629(.A(new_n743), .ZN(new_n816));
  INV_X1    g630(.A(new_n800), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n814), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n740), .A2(new_n808), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(KEYINPUT53), .A3(new_n795), .A4(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n812), .A2(new_n813), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n812), .A2(new_n824), .A3(new_n827), .A4(new_n813), .ZN(new_n828));
  INV_X1    g642(.A(new_n823), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n820), .A2(new_n821), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n830), .B2(new_n795), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n810), .A2(new_n783), .A3(new_n811), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT54), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n715), .A2(new_n716), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n535), .B1(new_n748), .B2(new_n749), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n773), .A2(new_n775), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n705), .A2(new_n369), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n706), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n732), .B(new_n837), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n696), .A2(new_n684), .A3(new_n671), .ZN(new_n842));
  NOR2_X1   g656(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n842), .A2(new_n836), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n842), .B2(new_n836), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n839), .A2(new_n189), .A3(new_n745), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n715), .A2(new_n681), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n835), .ZN(new_n849));
  INV_X1    g663(.A(new_n680), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n486), .A3(new_n536), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n529), .A2(new_n600), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n846), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n841), .A2(KEYINPUT51), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n852), .A2(new_n606), .A3(new_n847), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n533), .B(KEYINPUT117), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n857), .B(new_n858), .C1(new_n707), .C2(new_n836), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n726), .A3(new_n835), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n856), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT51), .B1(new_n841), .B2(new_n855), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n826), .A2(new_n828), .A3(new_n833), .A4(new_n866), .ZN(new_n867));
  OR2_X1    g681(.A1(G952), .A2(G953), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n746), .A2(new_n684), .A3(new_n189), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n716), .B(new_n870), .C1(new_n839), .C2(KEYINPUT49), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT111), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n850), .B(new_n671), .C1(KEYINPUT49), .C2(new_n839), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT118), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n869), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(G75));
  NOR2_X1   g695(.A1(new_n309), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n308), .B1(new_n812), .B2(new_n824), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(G210), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n249), .A2(new_n251), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n287), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT55), .Z(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n883), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n885), .A2(new_n889), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  INV_X1    g708(.A(new_n892), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n894), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(G51));
  NAND2_X1  g711(.A1(new_n812), .A2(new_n824), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(KEYINPUT120), .A3(new_n825), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n901), .A3(KEYINPUT54), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n762), .B(KEYINPUT57), .Z(new_n903));
  NAND3_X1  g717(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n694), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n884), .A2(new_n759), .A3(new_n760), .A4(new_n758), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n882), .B1(new_n905), .B2(new_n906), .ZN(G54));
  AND3_X1   g721(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n883), .B1(new_n908), .B2(new_n520), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n520), .B2(new_n908), .ZN(G60));
  AND2_X1   g724(.A1(new_n596), .A2(new_n597), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT59), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n911), .A2(new_n900), .A3(new_n902), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n826), .A2(new_n828), .A3(new_n833), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(new_n913), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n914), .A2(new_n916), .A3(new_n882), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n898), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n882), .B1(new_n920), .B2(new_n479), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n642), .A2(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n642), .A2(KEYINPUT122), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(KEYINPUT121), .A3(new_n924), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n921), .A2(new_n922), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(G66));
  OAI21_X1  g742(.A(G953), .B1(new_n538), .B2(new_n284), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n805), .A2(new_n806), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n886), .B1(G898), .B2(new_n309), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(G69));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n432), .A2(new_n486), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n663), .B(new_n732), .C1(new_n728), .C2(new_n803), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n768), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n778), .B2(new_n780), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n658), .A2(new_n690), .A3(new_n791), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n687), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n940), .B(KEYINPUT62), .C1(new_n665), .C2(new_n686), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n938), .A2(new_n947), .A3(new_n944), .ZN(new_n948));
  AOI21_X1  g762(.A(G953), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n386), .A2(new_n388), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n516), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT123), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n934), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n938), .A2(new_n947), .A3(new_n944), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n947), .B1(new_n938), .B2(new_n944), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(KEYINPUT125), .B(new_n952), .C1(new_n957), .C2(G953), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n652), .A2(G953), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n740), .A2(new_n816), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n767), .A2(new_n706), .A3(new_n662), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n726), .A2(new_n616), .A3(new_n529), .A4(new_n575), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n768), .B(new_n940), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  AOI211_X1 g778(.A(new_n961), .B(new_n964), .C1(new_n780), .C2(new_n778), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n960), .B1(new_n965), .B2(G953), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n951), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(KEYINPUT127), .B(new_n960), .C1(new_n965), .C2(G953), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT126), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n309), .B1(G227), .B2(G900), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n959), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n959), .B2(new_n970), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(new_n957), .A2(new_n930), .ZN(new_n975));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  AOI21_X1  g791(.A(new_n676), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n831), .A2(new_n832), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n676), .A2(new_n398), .A3(new_n977), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n965), .A2(new_n930), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n398), .B1(new_n982), .B2(new_n977), .ZN(new_n983));
  NOR4_X1   g797(.A1(new_n978), .A2(new_n882), .A3(new_n981), .A4(new_n983), .ZN(G57));
endmodule


