//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G227), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G107), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(new_n194), .B2(G107), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n200));
  INV_X1    g014(.A(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G104), .ZN(new_n202));
  INV_X1    g016(.A(G101), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n202), .A3(new_n203), .A4(new_n195), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n198), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT66), .A3(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n208), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT64), .A2(G146), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(G143), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT64), .A2(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(KEYINPUT64), .A2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT65), .A3(G143), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n212), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(KEYINPUT84), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n212), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT65), .B1(new_n221), .B2(G143), .ZN(new_n228));
  NOR4_X1   g042(.A1(new_n219), .A2(new_n220), .A3(new_n217), .A4(new_n210), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n227), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT84), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n210), .A2(G146), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n224), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n218), .A2(new_n222), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(new_n227), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n206), .B(new_n226), .C1(new_n232), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n224), .B1(new_n216), .B2(KEYINPUT1), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT64), .B(G146), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n233), .B1(new_n241), .B2(new_n210), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n234), .B1(new_n221), .B2(G143), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(new_n221), .B2(G143), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT69), .B(new_n244), .C1(new_n246), .C2(new_n224), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n230), .A3(new_n205), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n238), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G134), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT11), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT11), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n252), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(G131), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n260), .ZN(new_n263));
  INV_X1    g077(.A(new_n252), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G131), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n265), .A2(new_n266), .A3(new_n257), .A4(new_n255), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT12), .B1(new_n250), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  INV_X1    g084(.A(new_n268), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n270), .B(new_n271), .C1(new_n238), .C2(new_n249), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT10), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n199), .A2(new_n202), .A3(new_n195), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G101), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n204), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(KEYINPUT0), .A2(G128), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n236), .A2(new_n227), .A3(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(KEYINPUT0), .A2(G128), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n244), .A2(new_n284), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n282), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n238), .A2(new_n274), .B1(new_n279), .B2(new_n287), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n243), .A2(new_n247), .B1(new_n223), .B2(new_n225), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n205), .A2(new_n274), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT85), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n219), .A2(new_n220), .A3(new_n210), .ZN(new_n293));
  OAI21_X1  g107(.A(G128), .B1(new_n293), .B2(new_n245), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT69), .B1(new_n294), .B2(new_n244), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n240), .A2(new_n242), .A3(new_n239), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n230), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT85), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n290), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n292), .A2(new_n299), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n288), .A2(new_n300), .A3(new_n271), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n193), .B1(new_n273), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n238), .A2(new_n274), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n279), .A2(new_n287), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n289), .A2(KEYINPUT85), .A3(new_n291), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n297), .B2(new_n290), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n303), .B(new_n304), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n268), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n288), .A2(new_n300), .A3(new_n271), .ZN(new_n309));
  INV_X1    g123(.A(new_n193), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n187), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n309), .B(new_n310), .C1(new_n272), .C2(new_n269), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n308), .B2(new_n309), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n187), .B(new_n313), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT86), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n271), .B1(new_n288), .B2(new_n300), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n193), .B1(new_n301), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(G902), .B1(new_n322), .B2(new_n315), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(KEYINPUT86), .A3(new_n187), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n314), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G221), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT9), .B(G234), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n328), .B2(new_n313), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n329), .B(KEYINPUT80), .Z(new_n330));
  OAI21_X1  g144(.A(KEYINPUT87), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n312), .A2(new_n313), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G469), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n322), .A2(new_n315), .ZN(new_n334));
  AND4_X1   g148(.A1(KEYINPUT86), .A2(new_n334), .A3(new_n187), .A4(new_n313), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT86), .B1(new_n323), .B2(new_n187), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n338));
  INV_X1    g152(.A(new_n330), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT16), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT76), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(G125), .ZN(new_n346));
  INV_X1    g160(.A(G125), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G140), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n348), .A3(KEYINPUT16), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n350), .A2(new_n342), .A3(new_n343), .A4(G125), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n345), .A2(new_n349), .A3(G146), .A4(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n352), .B(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n214), .A2(new_n346), .A3(new_n348), .A4(new_n215), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n356));
  OAI211_X1 g170(.A(G119), .B(new_n224), .C1(new_n356), .C2(KEYINPUT23), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT23), .ZN(new_n358));
  INV_X1    g172(.A(G119), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(G128), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT74), .B1(new_n359), .B2(G128), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n362), .A2(G110), .ZN(new_n363));
  XNOR2_X1  g177(.A(G119), .B(G128), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT24), .B(G110), .Z(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n354), .A2(new_n355), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n364), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G110), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n371), .B1(new_n362), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n373), .B1(new_n372), .B2(new_n362), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n345), .A2(new_n349), .A3(new_n351), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n208), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n352), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(new_n374), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT77), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n367), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT22), .B(G137), .ZN(new_n383));
  INV_X1    g197(.A(G234), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n326), .A2(new_n384), .A3(G953), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n383), .B(new_n385), .Z(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n367), .B(new_n386), .C1(new_n380), .C2(new_n381), .ZN(new_n389));
  AOI21_X1  g203(.A(G902), .B1(new_n384), .B2(G217), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT79), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT79), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n389), .A3(new_n393), .A4(new_n390), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n313), .A3(new_n389), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n396), .A2(KEYINPUT25), .ZN(new_n397));
  OAI21_X1  g211(.A(G217), .B1(new_n384), .B2(G902), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n396), .B2(KEYINPUT25), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n395), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n257), .B1(new_n264), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n404));
  OAI21_X1  g218(.A(G131), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n267), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT72), .B1(new_n289), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT72), .ZN(new_n408));
  INV_X1    g222(.A(new_n406), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n297), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n282), .A2(new_n268), .A3(new_n285), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n407), .A2(new_n410), .A3(KEYINPUT30), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT71), .ZN(new_n413));
  XOR2_X1   g227(.A(KEYINPUT2), .B(G113), .Z(new_n414));
  INV_X1    g228(.A(KEYINPUT70), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n359), .B2(G116), .ZN(new_n416));
  INV_X1    g230(.A(G116), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT70), .A3(G119), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n359), .A2(G116), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n414), .B1(new_n420), .B2(new_n419), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n413), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n420), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT2), .B(G113), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT71), .A3(new_n421), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n411), .B1(new_n289), .B2(new_n406), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n412), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n407), .A2(new_n410), .A3(new_n429), .A4(new_n411), .ZN(new_n434));
  NOR2_X1   g248(.A1(G237), .A2(G953), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G210), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(KEYINPUT27), .Z(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT26), .B(G101), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n437), .B(new_n438), .Z(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT31), .B1(new_n433), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n439), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT28), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n434), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n429), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n430), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n430), .A2(new_n445), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n442), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n412), .A2(new_n432), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT31), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n434), .A4(new_n439), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(G472), .A2(G902), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT32), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n406), .B1(new_n248), .B2(new_n230), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n212), .B(new_n280), .C1(new_n218), .C2(new_n222), .ZN(new_n461));
  INV_X1    g275(.A(new_n285), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n460), .A2(new_n408), .B1(new_n268), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n429), .B1(new_n464), .B2(new_n407), .ZN(new_n465));
  INV_X1    g279(.A(new_n434), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT28), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n439), .A2(KEYINPUT29), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n446), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n313), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n439), .B1(new_n444), .B2(new_n448), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n450), .A2(new_n434), .A3(new_n442), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT29), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G472), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n401), .B1(new_n459), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(G475), .A2(G902), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n347), .A2(G140), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n343), .A2(G125), .ZN(new_n479));
  OAI21_X1  g293(.A(G146), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n477), .B1(new_n480), .B2(new_n355), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n355), .A3(new_n477), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n435), .A2(G143), .A3(G214), .ZN(new_n484));
  AOI21_X1  g298(.A(G143), .B1(new_n435), .B2(G214), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(KEYINPUT18), .A2(G131), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT92), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n482), .A2(new_n483), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n435), .A2(G214), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n210), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n435), .A2(G143), .A3(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT89), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n491), .A2(KEYINPUT89), .A3(new_n492), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT90), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n484), .B2(new_n485), .ZN(new_n498));
  INV_X1    g312(.A(new_n487), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n489), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n484), .B2(new_n485), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n491), .A2(new_n266), .A3(new_n492), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT96), .B1(new_n506), .B2(KEYINPUT17), .ZN(new_n507));
  AND2_X1   g321(.A1(new_n376), .A2(new_n352), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n504), .A2(new_n505), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n493), .A2(KEYINPUT17), .A3(G131), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n507), .A2(new_n508), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  XOR2_X1   g327(.A(G113), .B(G122), .Z(new_n514));
  XOR2_X1   g328(.A(KEYINPUT95), .B(G104), .Z(new_n515));
  XOR2_X1   g329(.A(new_n514), .B(new_n515), .Z(new_n516));
  AND3_X1   g330(.A1(new_n503), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G125), .B(G140), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT94), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT19), .B1(new_n478), .B2(new_n479), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n521), .A2(new_n523), .A3(new_n221), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n354), .A2(new_n506), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n516), .B1(new_n503), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n476), .B1(new_n517), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT97), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT20), .ZN(new_n530));
  INV_X1    g344(.A(new_n476), .ZN(new_n531));
  INV_X1    g345(.A(new_n516), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n486), .A2(new_n488), .ZN(new_n533));
  INV_X1    g347(.A(new_n483), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n481), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n495), .A2(KEYINPUT90), .A3(new_n496), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n500), .A2(new_n501), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n352), .A2(KEYINPUT78), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n349), .A2(new_n351), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(new_n353), .A3(G146), .A4(new_n345), .ZN(new_n541));
  AND4_X1   g355(.A1(new_n539), .A2(new_n525), .A3(new_n541), .A4(new_n506), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n532), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n503), .A2(new_n513), .A3(new_n516), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n531), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT97), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n530), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n516), .B1(new_n503), .B2(new_n513), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n313), .B1(new_n517), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G475), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n328), .A2(G217), .A3(new_n189), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n210), .A2(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n224), .A2(G143), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n256), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT99), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n256), .B1(new_n555), .B2(new_n556), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n556), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G134), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT99), .B1(new_n563), .B2(new_n557), .ZN(new_n564));
  INV_X1    g378(.A(G122), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G116), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n417), .A2(G122), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(KEYINPUT14), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(G107), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(new_n567), .C1(KEYINPUT14), .C2(new_n201), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g386(.A1(new_n561), .A2(new_n564), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n201), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n566), .A2(new_n567), .A3(G107), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n557), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT13), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n224), .B2(G143), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n210), .A2(KEYINPUT13), .A3(G128), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n556), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT98), .B1(new_n580), .B2(G134), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(KEYINPUT98), .A3(G134), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n576), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n554), .B1(new_n573), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n559), .B1(new_n558), .B2(new_n560), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n563), .A2(KEYINPUT99), .A3(new_n557), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n571), .A4(new_n570), .ZN(new_n588));
  INV_X1    g402(.A(new_n554), .ZN(new_n589));
  INV_X1    g403(.A(new_n583), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n581), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n588), .B(new_n589), .C1(new_n591), .C2(new_n576), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n585), .A2(new_n592), .A3(KEYINPUT100), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT100), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n594), .B(new_n554), .C1(new_n573), .C2(new_n584), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n313), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT101), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n598), .A3(new_n313), .A4(new_n595), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G478), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(KEYINPUT15), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n597), .B1(KEYINPUT15), .B2(new_n601), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(G234), .A2(G237), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(G952), .A3(new_n189), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(G902), .A3(G953), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT21), .B(G898), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n608), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n553), .A2(new_n605), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G214), .B1(G237), .B2(G902), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G210), .B1(G237), .B2(G902), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(G113), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT5), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n359), .A3(G116), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n620), .B2(KEYINPUT88), .ZN(new_n621));
  OAI221_X1 g435(.A(new_n621), .B1(KEYINPUT88), .B2(new_n620), .C1(new_n425), .C2(new_n619), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n421), .A3(new_n206), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n277), .B(KEYINPUT83), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n424), .A2(new_n428), .A3(new_n286), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(G110), .B(G122), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n627), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(KEYINPUT6), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(G224), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(G953), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n347), .B(new_n230), .C1(new_n295), .C2(new_n296), .ZN(new_n635));
  OAI21_X1  g449(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n635), .A2(new_n636), .A3(new_n634), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT6), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n626), .A2(new_n641), .A3(new_n628), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n631), .A2(new_n640), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n633), .A2(KEYINPUT7), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n638), .B2(new_n639), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n635), .A2(new_n636), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n644), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n627), .B(KEYINPUT8), .ZN(new_n648));
  INV_X1    g462(.A(new_n623), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n206), .B1(new_n622), .B2(new_n421), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n647), .A2(new_n630), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n313), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n617), .B1(new_n643), .B2(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n647), .A2(new_n630), .A3(new_n651), .ZN(new_n655));
  INV_X1    g469(.A(new_n639), .ZN(new_n656));
  OAI22_X1  g470(.A1(new_n656), .A2(new_n637), .B1(KEYINPUT7), .B2(new_n633), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n631), .A2(new_n640), .A3(new_n642), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n616), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n615), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n341), .A2(new_n475), .A3(new_n613), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G101), .ZN(G3));
  NAND2_X1  g477(.A1(new_n654), .A2(new_n660), .ZN(new_n664));
  INV_X1    g478(.A(new_n612), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n665), .A3(new_n614), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT33), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n593), .A2(new_n667), .A3(new_n595), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n585), .A2(new_n592), .A3(KEYINPUT33), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n668), .A2(G478), .A3(new_n313), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT102), .B(G478), .Z(new_n671));
  NAND2_X1  g485(.A1(new_n596), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n553), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n453), .A2(new_n313), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n455), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n401), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n341), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n194), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT103), .B(KEYINPUT34), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  OR2_X1    g497(.A1(new_n548), .A2(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n548), .A2(KEYINPUT104), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n530), .A4(new_n547), .ZN(new_n686));
  AND2_X1   g500(.A1(new_n686), .A2(new_n605), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(new_n552), .A3(new_n665), .A4(new_n661), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n341), .A2(new_n679), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT35), .B(G107), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G9));
  NAND2_X1  g506(.A1(new_n397), .A2(new_n399), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n387), .A2(KEYINPUT36), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n382), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n382), .A2(new_n695), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n390), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n693), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n678), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n341), .A2(new_n613), .A3(new_n661), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT37), .B(G110), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  AND3_X1   g519(.A1(new_n453), .A2(new_n457), .A3(new_n454), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n457), .B1(new_n453), .B2(new_n454), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n474), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n693), .A2(new_n699), .A3(new_n700), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT106), .B(G900), .Z(new_n710));
  AOI21_X1  g524(.A(new_n608), .B1(new_n710), .B2(new_n610), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n711), .B1(new_n551), .B2(G475), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n686), .A2(new_n605), .A3(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n708), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n325), .A2(KEYINPUT87), .A3(new_n330), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n338), .B1(new_n337), .B2(new_n339), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n714), .B(new_n661), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  XNOR2_X1  g532(.A(new_n664), .B(KEYINPUT38), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n549), .A2(new_n552), .B1(new_n603), .B2(new_n604), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(new_n614), .A3(new_n701), .A4(new_n720), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n465), .A2(new_n466), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n313), .B1(new_n722), .B2(new_n439), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n442), .B1(new_n450), .B2(new_n434), .ZN(new_n724));
  OAI21_X1  g538(.A(G472), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n459), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n711), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n341), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT40), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n730), .A2(KEYINPUT40), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n210), .ZN(G45));
  INV_X1    g550(.A(new_n711), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n553), .A2(new_n673), .A3(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n658), .A2(new_n616), .A3(new_n659), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n616), .B1(new_n658), .B2(new_n659), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n614), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT108), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n743));
  AOI22_X1  g557(.A1(new_n549), .A2(new_n552), .B1(new_n672), .B2(new_n670), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n661), .A2(new_n743), .A3(new_n744), .A4(new_n737), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n708), .A2(new_n742), .A3(new_n709), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n341), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G146), .ZN(G48));
  NAND2_X1  g562(.A1(new_n320), .A2(new_n324), .ZN(new_n749));
  INV_X1    g563(.A(new_n329), .ZN(new_n750));
  INV_X1    g564(.A(new_n323), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n475), .A3(new_n675), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  AOI22_X1  g571(.A1(new_n320), .A2(new_n324), .B1(G469), .B2(new_n751), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n708), .A3(new_n400), .A4(new_n750), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT109), .B1(new_n759), .B2(new_n688), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n754), .A2(new_n689), .A3(new_n475), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G116), .ZN(G18));
  AND4_X1   g578(.A1(new_n749), .A2(new_n750), .A3(new_n661), .A4(new_n752), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n701), .B1(new_n459), .B2(new_n474), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT110), .A4(new_n613), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n708), .A2(new_n613), .A3(new_n709), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n749), .A2(new_n750), .A3(new_n661), .A4(new_n752), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G119), .ZN(G21));
  NAND2_X1  g587(.A1(new_n441), .A2(new_n452), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n439), .B1(new_n467), .B2(new_n446), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n454), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n400), .A2(new_n677), .A3(new_n776), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n753), .A2(new_n777), .A3(new_n612), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT111), .B1(new_n553), .B2(new_n605), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n741), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n553), .A2(KEYINPUT111), .A3(new_n605), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n614), .B(new_n664), .C1(new_n720), .C2(KEYINPUT111), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT112), .B1(new_n785), .B2(new_n781), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n778), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G122), .ZN(G24));
  INV_X1    g603(.A(new_n738), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n677), .A3(new_n709), .A4(new_n776), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n770), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n347), .ZN(G27));
  INV_X1    g607(.A(KEYINPUT113), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n706), .B2(new_n707), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n456), .A2(KEYINPUT113), .A3(new_n458), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n474), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n400), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n654), .A2(new_n614), .A3(new_n660), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n337), .A2(new_n750), .A3(new_n790), .A4(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(KEYINPUT42), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n325), .A2(new_n329), .A3(new_n799), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n738), .A2(KEYINPUT42), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n475), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n266), .ZN(G33));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n475), .A3(new_n713), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n187), .B1(new_n312), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n810), .B2(new_n312), .ZN(new_n812));
  NAND2_X1  g626(.A1(G469), .A2(G902), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT46), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n320), .B2(new_n324), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(KEYINPUT46), .A3(new_n813), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n329), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n817), .A2(new_n729), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n549), .A2(new_n552), .A3(new_n673), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT43), .Z(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n678), .A3(new_n709), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT44), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n799), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n818), .B(new_n823), .C1(new_n822), .C2(new_n821), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G137), .ZN(G39));
  NOR4_X1   g639(.A1(new_n708), .A2(new_n400), .A3(new_n738), .A4(new_n799), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n817), .A2(KEYINPUT47), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n817), .A2(KEYINPUT47), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(KEYINPUT114), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G140), .ZN(G42));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n820), .A2(new_n608), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n777), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n719), .A2(new_n614), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n754), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n835), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n754), .A4(new_n839), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n754), .A2(new_n800), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n836), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n677), .A3(new_n709), .A4(new_n776), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n726), .A2(new_n400), .A3(new_n608), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n844), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n553), .A2(new_n673), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n843), .A2(KEYINPUT51), .A3(new_n846), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n827), .A2(new_n828), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n758), .A2(new_n330), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT120), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n838), .A2(new_n799), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n854), .B2(KEYINPUT120), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n851), .B1(new_n855), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n846), .A2(new_n850), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n853), .B(KEYINPUT118), .Z(new_n861));
  NAND2_X1  g675(.A1(new_n852), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n860), .B1(new_n862), .B2(new_n856), .ZN(new_n863));
  XOR2_X1   g677(.A(new_n843), .B(KEYINPUT119), .Z(new_n864));
  AOI21_X1  g678(.A(KEYINPUT51), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n798), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n845), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT48), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n848), .A2(new_n744), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n189), .A2(G952), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n837), .B2(new_n765), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n859), .A2(new_n865), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n325), .A2(new_n329), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n693), .A2(new_n700), .A3(new_n699), .A4(new_n737), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n875), .B1(new_n459), .B2(new_n725), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n783), .B1(new_n780), .B2(new_n782), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n785), .A2(KEYINPUT112), .A3(new_n781), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n874), .B(new_n876), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n792), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n717), .A2(new_n747), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n792), .B1(new_n341), .B2(new_n746), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT52), .A3(new_n717), .A4(new_n879), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n763), .A2(new_n662), .A3(new_n772), .A4(new_n703), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n605), .A2(new_n549), .A3(new_n552), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT116), .B1(new_n666), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n888), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n890), .A2(new_n661), .A3(new_n891), .A4(new_n665), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n341), .A2(new_n893), .A3(new_n679), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n680), .A2(new_n894), .A3(new_n755), .A4(new_n788), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n603), .A2(new_n686), .A3(new_n604), .A4(new_n712), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n708), .A2(new_n897), .A3(new_n709), .A4(new_n800), .ZN(new_n898));
  INV_X1    g712(.A(new_n791), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n341), .A2(new_n898), .B1(new_n899), .B2(new_n803), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n802), .A3(new_n805), .A4(new_n808), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n886), .A2(new_n896), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT53), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n887), .A2(new_n901), .A3(new_n895), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n882), .A2(KEYINPUT117), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n881), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g723(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n910));
  NAND4_X1  g724(.A1(new_n884), .A2(new_n717), .A3(new_n879), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n907), .A2(KEYINPUT53), .A3(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n905), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n907), .A2(new_n904), .A3(new_n912), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n904), .B1(new_n907), .B2(new_n886), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n917), .B2(new_n906), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n873), .A2(new_n918), .B1(G952), .B2(G953), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n758), .B(KEYINPUT49), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n400), .A2(new_n339), .A3(new_n614), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT115), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n719), .A2(new_n819), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n920), .A2(new_n922), .A3(new_n726), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n189), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n313), .B1(new_n905), .B2(new_n913), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(G210), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n631), .A2(new_n642), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(new_n640), .Z(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT55), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT122), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n927), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n933), .ZN(new_n936));
  OR3_X1    g750(.A1(new_n929), .A2(KEYINPUT121), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT121), .B1(new_n929), .B2(new_n936), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G51));
  AOI211_X1 g753(.A(new_n313), .B(new_n812), .C1(new_n905), .C2(new_n913), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n813), .B(KEYINPUT57), .Z(new_n941));
  AND3_X1   g755(.A1(new_n907), .A2(KEYINPUT53), .A3(new_n912), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT53), .B1(new_n907), .B2(new_n886), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT54), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n906), .B1(new_n905), .B2(new_n913), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n941), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n940), .B1(new_n946), .B2(new_n334), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT123), .B1(new_n947), .B2(new_n926), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT54), .B1(new_n942), .B2(new_n943), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n914), .ZN(new_n951));
  AOI22_X1  g765(.A1(new_n951), .A2(new_n941), .B1(new_n322), .B2(new_n315), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n949), .B(new_n927), .C1(new_n952), .C2(new_n940), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(new_n953), .ZN(G54));
  NAND3_X1  g768(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n543), .A2(new_n544), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n955), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n958), .A2(new_n959), .A3(new_n926), .ZN(G60));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT59), .Z(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI22_X1  g777(.A1(new_n918), .A2(new_n963), .B1(new_n668), .B2(new_n669), .ZN(new_n964));
  INV_X1    g778(.A(new_n951), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n668), .A2(new_n669), .A3(new_n963), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n927), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n964), .A2(new_n967), .ZN(G63));
  NAND2_X1  g782(.A1(new_n905), .A2(new_n913), .ZN(new_n969));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT60), .Z(new_n971));
  NAND2_X1  g785(.A1(new_n696), .A2(new_n697), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT124), .Z(new_n973));
  NAND3_X1  g787(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n969), .A2(new_n971), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n388), .A2(new_n389), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n927), .B(new_n974), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT61), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G66));
  OAI21_X1  g793(.A(G953), .B1(new_n611), .B2(new_n632), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n896), .B(KEYINPUT125), .Z(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(G953), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n931), .B1(G898), .B2(new_n189), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT126), .Z(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  NAND3_X1  g799(.A1(new_n818), .A2(new_n787), .A3(new_n866), .ZN(new_n986));
  AND4_X1   g800(.A1(new_n717), .A2(new_n824), .A3(new_n986), .A4(new_n884), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n802), .A2(new_n805), .A3(new_n808), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n987), .A2(new_n833), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n189), .ZN(new_n990));
  INV_X1    g804(.A(new_n430), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n412), .B1(KEYINPUT30), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n521), .A2(new_n524), .A3(new_n523), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n992), .B(new_n993), .Z(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(G900), .B2(G953), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n884), .A2(new_n717), .ZN(new_n996));
  OR3_X1    g810(.A1(new_n735), .A2(KEYINPUT62), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT62), .B1(new_n735), .B2(new_n996), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n799), .B1(new_n674), .B2(new_n888), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n731), .A2(new_n475), .A3(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n824), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n833), .A2(new_n997), .A3(new_n998), .A4(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n189), .ZN(new_n1003));
  AOI22_X1  g817(.A1(new_n990), .A2(new_n995), .B1(new_n1003), .B2(new_n994), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n987), .A2(new_n833), .A3(new_n988), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n995), .B1(new_n1006), .B2(G953), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1005), .B1(new_n1007), .B2(KEYINPUT127), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1004), .B(new_n1008), .ZN(G72));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n989), .B2(new_n981), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n927), .B1(new_n1013), .B2(new_n472), .ZN(new_n1014));
  INV_X1    g828(.A(new_n724), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1002), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n981), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1015), .B1(new_n1017), .B2(new_n1011), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n472), .A3(new_n1011), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n917), .A2(new_n1019), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1014), .A2(new_n1018), .A3(new_n1020), .ZN(G57));
endmodule


