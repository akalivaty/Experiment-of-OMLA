//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT67), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n191), .A2(KEYINPUT67), .A3(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G131), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT69), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT69), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(G143), .B2(new_n196), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n200), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n197), .A2(new_n199), .A3(new_n206), .A4(G128), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n188), .A2(new_n195), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n195), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT68), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n213), .B1(new_n189), .B2(G137), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT11), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n213), .B(new_n217), .C1(new_n189), .C2(G137), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n190), .A4(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n210), .B(new_n212), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n217), .B1(new_n192), .B2(new_n213), .ZN(new_n223));
  AOI211_X1 g037(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n191), .C2(G134), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n216), .A4(new_n190), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n219), .A2(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n190), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n227), .A2(new_n228), .B1(new_n229), .B2(G131), .ZN(new_n230));
  XNOR2_X1  g044(.A(G143), .B(G146), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT0), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(new_n201), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n201), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n200), .A2(new_n233), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n222), .B(KEYINPUT30), .C1(new_n230), .C2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(KEYINPUT2), .B(G113), .Z(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT70), .B(G119), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n240), .B(new_n243), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n241), .A2(KEYINPUT70), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G119), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n244), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n247), .B1(new_n251), .B2(new_n242), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n227), .A2(new_n228), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n229), .A2(G131), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT64), .B1(new_n236), .B2(new_n237), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n200), .B1(new_n233), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT64), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n260), .B(new_n261), .C1(new_n200), .C2(new_n233), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n227), .A2(new_n228), .B1(KEYINPUT68), .B2(new_n211), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n257), .A2(new_n264), .B1(new_n265), .B2(new_n210), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n239), .B(new_n254), .C1(new_n266), .C2(KEYINPUT30), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n222), .B(new_n253), .C1(new_n230), .C2(new_n238), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n238), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n257), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n272), .A2(KEYINPUT71), .A3(new_n253), .A4(new_n222), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(G101), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G953), .ZN(new_n279));
  AOI21_X1  g093(.A(G237), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G210), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n275), .B(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n267), .A2(new_n270), .A3(new_n273), .A4(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT31), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n270), .A2(new_n273), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n267), .A4(new_n282), .ZN(new_n287));
  INV_X1    g101(.A(new_n268), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(KEYINPUT28), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n222), .B1(new_n230), .B2(new_n263), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n254), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n270), .A2(new_n291), .A3(new_n273), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n284), .B(new_n287), .C1(new_n282), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n295), .B1(new_n294), .B2(new_n296), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n187), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n284), .A2(new_n287), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n293), .A2(new_n282), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT32), .B(new_n296), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n294), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n296), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT29), .B1(new_n293), .B2(new_n282), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n285), .A2(new_n267), .ZN(new_n308));
  INV_X1    g122(.A(new_n282), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n272), .A2(new_n222), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n270), .B(new_n273), .C1(new_n313), .C2(new_n253), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT28), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(KEYINPUT28), .B2(new_n288), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n282), .A2(KEYINPUT29), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n311), .B(new_n312), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G472), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n299), .A2(new_n306), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n278), .A2(G953), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n276), .A2(KEYINPUT72), .ZN(new_n324));
  OAI211_X1 g138(.A(G214), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n198), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n280), .A2(G143), .A3(G214), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n216), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT92), .B1(new_n329), .B2(G131), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n331));
  AOI211_X1 g145(.A(new_n331), .B(new_n216), .C1(new_n326), .C2(new_n327), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n321), .B(new_n328), .C1(new_n330), .C2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n335));
  INV_X1    g149(.A(G140), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G125), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n335), .B1(KEYINPUT16), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(G146), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n277), .A2(new_n279), .ZN(new_n340));
  AND4_X1   g154(.A1(G143), .A2(new_n340), .A3(G214), .A4(new_n322), .ZN(new_n341));
  AOI21_X1  g155(.A(G143), .B1(new_n280), .B2(G214), .ZN(new_n342));
  OAI21_X1  g156(.A(G131), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n331), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n329), .A2(KEYINPUT92), .A3(G131), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(KEYINPUT17), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n333), .A2(new_n339), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  INV_X1    g162(.A(G104), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n348), .B(new_n349), .ZN(new_n350));
  OAI211_X1 g164(.A(KEYINPUT18), .B(G131), .C1(new_n341), .C2(new_n342), .ZN(new_n351));
  NAND2_X1  g165(.A1(KEYINPUT18), .A2(G131), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n326), .A2(new_n327), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT76), .B1(new_n334), .B2(new_n196), .ZN(new_n354));
  AND2_X1   g168(.A1(G125), .A2(G140), .ZN(new_n355));
  NOR2_X1   g169(.A1(G125), .A2(G140), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT76), .B(new_n196), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI22_X1  g172(.A1(new_n354), .A2(new_n358), .B1(new_n196), .B2(new_n334), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n351), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT91), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n353), .A2(new_n359), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT91), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n351), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n347), .A2(new_n350), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n350), .B1(new_n347), .B2(new_n365), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n312), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G475), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n276), .A2(G952), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(G234), .B2(G237), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n312), .B(new_n340), .C1(G234), .C2(G237), .ZN(new_n373));
  XOR2_X1   g187(.A(KEYINPUT21), .B(G898), .Z(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n372), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n363), .B1(new_n362), .B2(new_n351), .ZN(new_n379));
  AND4_X1   g193(.A1(new_n363), .A2(new_n351), .A3(new_n353), .A4(new_n359), .ZN(new_n380));
  INV_X1    g194(.A(new_n328), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n344), .B2(new_n345), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n338), .A2(new_n196), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n334), .B(KEYINPUT19), .Z(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(G146), .ZN(new_n385));
  OAI22_X1  g199(.A1(new_n379), .A2(new_n380), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n350), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n366), .ZN(new_n389));
  INV_X1    g203(.A(G475), .ZN(new_n390));
  AND4_X1   g204(.A1(new_n378), .A2(new_n389), .A3(new_n390), .A4(new_n312), .ZN(new_n391));
  AOI21_X1  g205(.A(G475), .B1(new_n388), .B2(new_n366), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n378), .B1(new_n392), .B2(new_n312), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n370), .B(new_n377), .C1(new_n391), .C2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT69), .B(G128), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(new_n198), .ZN(new_n396));
  OAI21_X1  g210(.A(G134), .B1(new_n396), .B2(KEYINPUT13), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n198), .A2(G128), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n395), .B2(new_n198), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n244), .A2(G122), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n244), .A2(KEYINPUT93), .A3(G122), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT93), .B1(new_n244), .B2(G122), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(G107), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g220(.A(KEYINPUT9), .B(G234), .Z(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(G217), .A3(new_n276), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT94), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G107), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n401), .B2(KEYINPUT14), .ZN(new_n412));
  XOR2_X1   g226(.A(new_n404), .B(new_n412), .Z(new_n413));
  XNOR2_X1  g227(.A(new_n399), .B(G134), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n406), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n410), .B1(new_n406), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n312), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT95), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G478), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT15), .ZN(new_n422));
  OAI211_X1 g236(.A(KEYINPUT95), .B(new_n312), .C1(new_n416), .C2(new_n417), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n422), .B2(new_n418), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n394), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G221), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(new_n407), .B2(new_n312), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT80), .ZN(new_n430));
  INV_X1    g244(.A(new_n340), .ZN(new_n431));
  INV_X1    g245(.A(G227), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n430), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT3), .B1(new_n349), .B2(G107), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT3), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n411), .A3(G104), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n349), .A2(G107), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT82), .A3(G101), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT4), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n440), .A2(KEYINPUT82), .A3(new_n443), .A4(G101), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n436), .A2(new_n438), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT81), .ZN(new_n447));
  INV_X1    g261(.A(G101), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .A4(new_n439), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n436), .A2(new_n438), .A3(new_n448), .A4(new_n439), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n440), .A2(G101), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n445), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n271), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n449), .A2(new_n451), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n201), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT84), .B1(new_n457), .B2(new_n231), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT84), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n200), .B(new_n459), .C1(new_n201), .C2(new_n207), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n209), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n231), .A2(KEYINPUT83), .A3(new_n206), .A4(G128), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n458), .A2(new_n460), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n411), .A2(G104), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n448), .B1(new_n439), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n456), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n208), .A2(new_n209), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT10), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT85), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n466), .B1(new_n449), .B2(new_n451), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n469), .B1(new_n208), .B2(new_n209), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n455), .A2(new_n470), .A3(new_n476), .A4(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(new_n257), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n473), .A2(KEYINPUT85), .A3(new_n475), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n271), .A2(new_n454), .B1(new_n468), .B2(new_n469), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n230), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n435), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT87), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n490), .B(new_n435), .C1(new_n482), .C2(new_n487), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n485), .A2(new_n486), .A3(new_n230), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n473), .A2(new_n208), .A3(new_n209), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n230), .B1(new_n493), .B2(new_n468), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n494), .A2(KEYINPUT12), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(KEYINPUT12), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n492), .B(new_n434), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n489), .A2(new_n491), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT86), .B(G469), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n312), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n482), .A2(new_n435), .ZN(new_n501));
  INV_X1    g315(.A(new_n487), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n435), .ZN(new_n504));
  OAI21_X1  g318(.A(G469), .B1(new_n504), .B2(G902), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n428), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G214), .B1(G237), .B2(G902), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n509));
  XNOR2_X1  g323(.A(G110), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT88), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n253), .B1(new_n445), .B2(new_n453), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT5), .B(new_n243), .C1(new_n245), .C2(new_n244), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n248), .A2(new_n250), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT5), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(G116), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(G113), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n246), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n473), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n509), .B(new_n512), .C1(new_n513), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT89), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n477), .A2(new_n246), .A3(new_n518), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n450), .B(new_n447), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n524), .A2(new_n452), .B1(new_n442), .B2(new_n444), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n523), .B1(new_n525), .B2(new_n253), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT89), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n509), .A4(new_n512), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G125), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n474), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n238), .B2(new_n530), .ZN(new_n532));
  INV_X1    g346(.A(G224), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n534), .B(KEYINPUT90), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n532), .B(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n526), .A2(new_n512), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n523), .B(new_n511), .C1(new_n525), .C2(new_n253), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(KEYINPUT6), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n529), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n511), .B(KEYINPUT8), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n473), .A2(new_n519), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n520), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT7), .B1(new_n533), .B2(G953), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n532), .B(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n540), .A2(new_n549), .A3(new_n547), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n508), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n426), .A2(new_n506), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT23), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n245), .A2(new_n555), .A3(new_n201), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n241), .A2(new_n395), .B1(new_n245), .B2(new_n201), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n555), .ZN(new_n558));
  INV_X1    g372(.A(G110), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT24), .B(G110), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n558), .A2(new_n559), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n354), .A2(new_n358), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n562), .A2(new_n383), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n557), .A2(new_n560), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n339), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n559), .B2(new_n558), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT77), .B(KEYINPUT78), .Z(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT22), .B(G137), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND3_X1  g387(.A1(new_n565), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n565), .B2(new_n568), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT25), .B1(new_n577), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(G217), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(G234), .B2(new_n312), .ZN(new_n580));
  INV_X1    g394(.A(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n574), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT25), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n312), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n578), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT79), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n580), .A2(G902), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n586), .B(new_n587), .C1(new_n575), .C2(new_n576), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n320), .A2(new_n554), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G101), .ZN(G3));
  OAI21_X1  g408(.A(new_n370), .B1(new_n391), .B2(new_n393), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT33), .B1(new_n416), .B2(KEYINPUT97), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n596), .B1(new_n416), .B2(new_n417), .ZN(new_n597));
  INV_X1    g411(.A(new_n416), .ZN(new_n598));
  INV_X1    g412(.A(new_n417), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n598), .A2(KEYINPUT97), .A3(new_n599), .A4(KEYINPUT33), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n597), .A2(G478), .A3(new_n312), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n420), .A2(new_n421), .A3(new_n423), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n551), .A2(KEYINPUT96), .A3(new_n552), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n549), .B1(new_n540), .B2(new_n547), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n508), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n604), .A2(new_n609), .A3(new_n376), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n294), .B2(new_n312), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n294), .A2(new_n296), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT73), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n428), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n585), .A2(new_n591), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n500), .A2(new_n505), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n611), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT98), .B(KEYINPUT99), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT34), .B(G104), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n392), .A2(new_n312), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT20), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n392), .A2(new_n378), .A3(new_n312), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n393), .A2(KEYINPUT100), .ZN(new_n632));
  OAI211_X1 g446(.A(new_n425), .B(new_n370), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n633), .A2(new_n376), .A3(new_n609), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n621), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT35), .B(G107), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  AND3_X1   g452(.A1(new_n620), .A2(new_n618), .A3(new_n553), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n565), .A2(new_n568), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n587), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n585), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n639), .A2(new_n426), .A3(new_n617), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT37), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n559), .ZN(G12));
  INV_X1    g461(.A(G900), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n372), .B1(new_n373), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n651), .A2(new_n633), .A3(new_n609), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n652), .A2(new_n320), .A3(new_n506), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  INV_X1    g468(.A(new_n552), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n606), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT101), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT38), .Z(new_n658));
  INV_X1    g472(.A(new_n425), .ZN(new_n659));
  INV_X1    g473(.A(new_n595), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n308), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n309), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n312), .B1(new_n314), .B2(new_n282), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n299), .A2(new_n306), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n667), .A2(new_n508), .A3(new_n644), .ZN(new_n668));
  INV_X1    g482(.A(new_n506), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n649), .B(KEYINPUT39), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  NAND3_X1  g486(.A1(new_n661), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  INV_X1    g488(.A(new_n644), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n609), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n604), .A2(new_n649), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n320), .A2(new_n676), .A3(new_n506), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  AND2_X1   g493(.A1(new_n498), .A2(new_n312), .ZN(new_n680));
  INV_X1    g494(.A(G469), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n618), .B(new_n500), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n320), .A2(new_n592), .A3(new_n683), .A4(new_n610), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND4_X1  g500(.A1(new_n634), .A2(new_n320), .A3(new_n592), .A4(new_n683), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT102), .B(G116), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G18));
  NAND4_X1  g503(.A1(new_n320), .A2(new_n676), .A3(new_n683), .A4(new_n426), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NAND2_X1  g505(.A1(new_n316), .A2(new_n309), .ZN(new_n692));
  INV_X1    g506(.A(new_n300), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n296), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n294), .A2(new_n312), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT103), .B(G472), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND4_X1   g512(.A1(new_n585), .A2(new_n695), .A3(new_n591), .A4(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n609), .A2(new_n660), .A3(new_n659), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n699), .A2(new_n683), .A3(new_n700), .A4(new_n377), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  INV_X1    g516(.A(new_n604), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n695), .A3(new_n698), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n651), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n682), .A2(new_n609), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT104), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  NAND3_X1  g524(.A1(new_n551), .A2(new_n507), .A3(new_n552), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n551), .A2(KEYINPUT105), .A3(new_n507), .A4(new_n552), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n713), .A2(new_n620), .A3(new_n618), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n506), .A2(KEYINPUT106), .A3(new_n713), .A4(new_n714), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n320), .A3(new_n592), .A4(new_n677), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n614), .A2(new_n187), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n319), .A2(new_n302), .A3(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n592), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n719), .A3(KEYINPUT42), .A4(new_n677), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  NOR2_X1   g542(.A1(new_n633), .A2(new_n649), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n719), .A2(new_n320), .A3(new_n592), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  NAND2_X1  g545(.A1(new_n660), .A2(new_n603), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT43), .Z(new_n733));
  INV_X1    g547(.A(new_n617), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n644), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n504), .B(KEYINPUT45), .Z(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(G902), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n500), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n618), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n670), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n735), .A2(new_n736), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n713), .A2(new_n714), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n746), .B(KEYINPUT108), .Z(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n737), .A2(new_n744), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n743), .B1(new_n751), .B2(KEYINPUT47), .ZN(new_n752));
  INV_X1    g566(.A(new_n746), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n754));
  NAND3_X1  g568(.A1(new_n742), .A2(new_n618), .A3(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n752), .A2(new_n677), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n320), .A2(new_n592), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n336), .ZN(G42));
  NOR2_X1   g573(.A1(new_n680), .A2(new_n681), .ZN(new_n760));
  INV_X1    g574(.A(new_n500), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(KEYINPUT110), .A2(KEYINPUT49), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n732), .B1(KEYINPUT110), .B2(KEYINPUT49), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n507), .A2(new_n658), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n762), .A2(new_n763), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n619), .A3(new_n667), .A4(new_n767), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT111), .Z(new_n769));
  AND2_X1   g583(.A1(new_n733), .A2(new_n372), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n683), .A3(new_n699), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT50), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n658), .A2(new_n508), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(new_n775));
  INV_X1    g589(.A(new_n603), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n746), .A2(new_n682), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n592), .A2(new_n667), .A3(new_n372), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(new_n660), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n774), .A2(new_n775), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n770), .A2(new_n777), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n644), .A3(new_n695), .A4(new_n698), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n752), .A2(new_n755), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n762), .A2(new_n428), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n770), .A2(new_n699), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n748), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n780), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n787), .A4(new_n782), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n781), .A2(new_n725), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT116), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n371), .B1(new_n793), .B2(KEYINPUT48), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n790), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n786), .A2(new_n707), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n377), .B(new_n507), .C1(new_n655), .C2(new_n606), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n425), .B(new_n370), .C1(new_n393), .C2(new_n391), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n797), .B1(new_n604), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n617), .A3(new_n620), .A4(new_n619), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n645), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n730), .A2(new_n593), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n719), .A2(new_n705), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n370), .B1(new_n631), .B2(new_n632), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n746), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n320), .A2(new_n805), .A3(new_n659), .A4(new_n506), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n651), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n687), .A2(new_n690), .A3(new_n684), .A4(new_n701), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n722), .B2(new_n726), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n811), .B1(new_n808), .B2(new_n810), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n669), .B1(new_n815), .B2(new_n649), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n649), .A2(new_n815), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n609), .A2(new_n660), .A3(new_n659), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n816), .A2(new_n818), .A3(new_n666), .A4(new_n675), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n653), .A3(new_n678), .A4(new_n708), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT53), .B1(new_n814), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n593), .A2(new_n645), .A3(new_n800), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n320), .A2(new_n592), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n717), .B2(new_n718), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n824), .B1(new_n826), .B2(new_n729), .ZN(new_n827));
  INV_X1    g641(.A(new_n809), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n320), .A2(new_n805), .A3(new_n659), .A4(new_n506), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n704), .B1(new_n717), .B2(new_n718), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n706), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n727), .A2(new_n827), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT112), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n822), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT54), .B1(new_n823), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT114), .B1(new_n802), .B2(new_n807), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(new_n810), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n836), .B1(new_n808), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n840), .A2(new_n841), .A3(new_n843), .A4(new_n822), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n593), .A2(new_n645), .A3(new_n800), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n831), .A2(new_n842), .A3(new_n730), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n839), .A2(new_n810), .A3(new_n846), .A4(KEYINPUT53), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n820), .B(KEYINPUT52), .ZN(new_n848));
  OAI21_X1  g662(.A(KEYINPUT115), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n835), .A2(new_n836), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n795), .A2(new_n796), .A3(new_n838), .A4(new_n853), .ZN(new_n854));
  AOI211_X1 g668(.A(KEYINPUT116), .B(KEYINPUT48), .C1(new_n781), .C2(new_n725), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n778), .A2(new_n703), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n769), .B1(new_n857), .B2(new_n858), .ZN(G75));
  NOR2_X1   g673(.A1(new_n340), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n312), .B1(new_n850), .B2(new_n851), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT56), .B1(new_n862), .B2(G210), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n529), .A2(new_n539), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(new_n536), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT55), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n861), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT117), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n862), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n550), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(G51));
  NAND2_X1  g687(.A1(new_n850), .A2(new_n851), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(KEYINPUT118), .A3(new_n853), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n877), .A3(KEYINPUT54), .ZN(new_n878));
  NAND2_X1  g692(.A1(G469), .A2(G902), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT57), .Z(new_n880));
  NAND3_X1  g694(.A1(new_n876), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n498), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n738), .A2(G469), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT119), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n869), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n860), .B1(new_n882), .B2(new_n885), .ZN(G54));
  NAND4_X1  g700(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .A4(new_n389), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n874), .A2(G902), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n868), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n862), .A2(KEYINPUT117), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n389), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n887), .A2(new_n893), .A3(new_n861), .ZN(G60));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n597), .A2(new_n600), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(G478), .A2(G902), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT59), .Z(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n876), .A2(new_n878), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n899), .B1(new_n838), .B2(new_n853), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n861), .B1(new_n902), .B2(new_n896), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n895), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n838), .A2(new_n853), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n897), .B1(new_n905), .B2(new_n899), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n876), .A2(new_n878), .A3(new_n900), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT120), .A4(new_n861), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT60), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n874), .A2(new_n642), .A3(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n874), .A2(new_n911), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n582), .B(KEYINPUT121), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n861), .B(new_n912), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT61), .Z(G66));
  NOR2_X1   g730(.A1(new_n809), .A2(new_n824), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n340), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT122), .ZN(new_n920));
  OAI21_X1  g734(.A(G953), .B1(new_n375), .B2(new_n533), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n864), .B1(G898), .B2(new_n340), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(G69));
  AOI21_X1  g738(.A(new_n825), .B1(new_n604), .B2(new_n798), .ZN(new_n925));
  INV_X1    g739(.A(new_n671), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n753), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n749), .B(new_n927), .C1(new_n756), .C2(new_n757), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n653), .A2(new_n678), .A3(new_n708), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n673), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n673), .A2(new_n931), .A3(new_n932), .A4(new_n930), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n929), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n239), .B1(new_n266), .B2(KEYINPUT30), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(new_n384), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n936), .A2(new_n340), .A3(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n744), .A2(new_n700), .A3(new_n725), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n749), .B(new_n940), .C1(new_n756), .C2(new_n757), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n727), .A2(new_n730), .A3(new_n930), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n340), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n648), .B2(new_n431), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT124), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n431), .B1(new_n432), .B2(new_n648), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G72));
  XNOR2_X1  g762(.A(new_n835), .B(new_n836), .ZN(new_n949));
  XNOR2_X1  g763(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n612), .A2(new_n312), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n950), .B(new_n951), .Z(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n310), .B2(new_n283), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT126), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n952), .B1(new_n936), .B2(new_n918), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n860), .B1(new_n958), .B2(new_n663), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n941), .A2(new_n918), .A3(new_n942), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n662), .B(new_n309), .C1(new_n960), .C2(new_n953), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n956), .A2(new_n957), .A3(new_n959), .A4(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n955), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n949), .B2(new_n954), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n959), .B(new_n961), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT127), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n962), .A2(new_n967), .ZN(G57));
endmodule


