//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n206), .B1(new_n207), .B2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G13), .ZN(new_n209));
  NAND4_X1  g0009(.A1(new_n209), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n207), .B1(new_n215), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n213), .B(new_n221), .C1(new_n224), .C2(new_n227), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G351));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n222), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n202), .B1(new_n245), .B2(G20), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n250), .A2(new_n251), .B1(new_n202), .B2(new_n247), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G150), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n223), .A2(G33), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(G20), .B2(new_n203), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n248), .A2(new_n222), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1698), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G222), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n264), .ZN(new_n268));
  INV_X1    g0068(.A(G223), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(G1698), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n266), .B1(new_n267), .B2(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT67), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(new_n222), .ZN(new_n274));
  AND2_X1   g0074(.A1(G1), .A2(G13), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G274), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n275), .B2(new_n276), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n245), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n275), .A2(new_n276), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n285), .B1(G226), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n279), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n260), .B1(new_n291), .B2(G169), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n290), .A2(G179), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G190), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT70), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(G200), .B2(new_n290), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n260), .B(KEYINPUT69), .Z(new_n298));
  AND2_X1   g0098(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n303), .B(new_n297), .C1(new_n299), .C2(new_n300), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n294), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT17), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n255), .B1(new_n245), .B2(G20), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(new_n250), .B1(new_n247), .B2(new_n255), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n263), .A2(new_n223), .A3(new_n264), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT7), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n264), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT73), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT73), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n309), .B2(new_n310), .ZN(new_n315));
  OAI21_X1  g0115(.A(G68), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G58), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(G20), .B1(new_n319), .B2(new_n201), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n253), .A2(G159), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT16), .B1(new_n316), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT3), .A2(G33), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(KEYINPUT7), .B1(new_n327), .B2(new_n223), .ZN(new_n328));
  INV_X1    g0128(.A(new_n312), .ZN(new_n329));
  OAI21_X1  g0129(.A(G68), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n330), .A2(KEYINPUT16), .A3(new_n323), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n249), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n308), .B1(new_n324), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G232), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n284), .B1(new_n287), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G87), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n262), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(G223), .A2(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(G226), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(G1698), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n341), .B2(new_n268), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT74), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n278), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G1698), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(G1698), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n346), .B(new_n347), .C1(new_n325), .C2(new_n326), .ZN(new_n348));
  INV_X1    g0148(.A(new_n338), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(KEYINPUT74), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n295), .B(new_n336), .C1(new_n344), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n274), .A2(new_n277), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n350), .B2(KEYINPUT74), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n342), .A2(new_n343), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n335), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n352), .B1(G200), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n306), .B1(new_n333), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n308), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n314), .B1(new_n328), .B2(new_n329), .ZN(new_n362));
  INV_X1    g0162(.A(new_n315), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n318), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n361), .B1(new_n364), .B2(new_n322), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n311), .A2(new_n312), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n322), .B1(new_n366), .B2(G68), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n259), .B1(new_n367), .B2(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n360), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT17), .A3(new_n357), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n359), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n356), .A2(G179), .ZN(new_n373));
  INV_X1    g0173(.A(G169), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n356), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n333), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(new_n333), .B2(new_n375), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n265), .A2(G232), .ZN(new_n382));
  INV_X1    g0182(.A(G107), .ZN(new_n383));
  INV_X1    g0183(.A(G238), .ZN(new_n384));
  OAI221_X1 g0184(.A(new_n382), .B1(new_n383), .B2(new_n268), .C1(new_n384), .C2(new_n270), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n278), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n285), .B1(G244), .B2(new_n288), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n381), .B1(new_n388), .B2(new_n374), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(G179), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n255), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n253), .B1(G20), .B2(G77), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(new_n256), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n259), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n245), .A2(G20), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n250), .A2(G77), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(G77), .B2(new_n246), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n390), .B2(KEYINPUT68), .ZN(new_n401));
  AOI211_X1 g0201(.A(new_n396), .B(new_n399), .C1(new_n388), .C2(G200), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n386), .A2(G190), .A3(new_n387), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n391), .A2(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n284), .B1(new_n287), .B2(new_n384), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G226), .A2(G1698), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n334), .B2(G1698), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n408), .A2(new_n268), .B1(G33), .B2(G97), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n409), .A2(KEYINPUT71), .A3(new_n353), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT71), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n334), .A2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G226), .B2(G1698), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n414), .B2(new_n327), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n411), .B1(new_n278), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n406), .B1(new_n410), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n406), .C1(new_n410), .C2(new_n416), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT72), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(KEYINPUT72), .A3(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(G200), .A3(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n318), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n425), .B1(new_n267), .B2(new_n256), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n426), .A2(new_n249), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(KEYINPUT11), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n247), .A2(new_n318), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT12), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(KEYINPUT11), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n250), .A2(G68), .A3(new_n397), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n428), .A2(new_n430), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n295), .B1(new_n417), .B2(KEYINPUT13), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n420), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n424), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n305), .A2(new_n380), .A3(new_n404), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n418), .A2(new_n420), .A3(G179), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n422), .A2(G169), .A3(new_n423), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n422), .A2(KEYINPUT14), .A3(G169), .A4(new_n423), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n433), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n223), .B(G87), .C1(new_n325), .C2(new_n326), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT22), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT24), .ZN(new_n451));
  INV_X1    g0251(.A(G116), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n262), .A2(new_n452), .A3(G20), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT23), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n223), .B2(G107), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n383), .A2(KEYINPUT23), .A3(G20), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n450), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n451), .B1(new_n450), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n249), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n245), .A2(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n259), .A2(new_n246), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT25), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n246), .B2(G107), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g0265(.A1(new_n246), .A2(new_n463), .A3(G107), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n383), .A2(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n460), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT79), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n460), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  OAI211_X1 g0272(.A(G250), .B(new_n345), .C1(new_n325), .C2(new_n326), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT80), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G294), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n477), .C1(new_n473), .C2(KEYINPUT80), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n278), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g0279(.A(KEYINPUT5), .B(G41), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n245), .A2(G45), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n281), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n273), .A2(new_n222), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n482), .B2(new_n480), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G264), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n479), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G169), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n268), .A2(new_n490), .A3(G250), .A4(new_n345), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n474), .A2(new_n491), .A3(new_n476), .A4(new_n477), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(new_n278), .B1(G264), .B2(new_n486), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(G179), .A3(new_n484), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n470), .A2(new_n472), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT81), .B1(new_n488), .B2(G190), .ZN(new_n497));
  INV_X1    g0297(.A(G200), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT81), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n493), .A2(new_n500), .A3(new_n295), .A4(new_n484), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n459), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n450), .A2(new_n451), .A3(new_n457), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n467), .B1(new_n505), .B2(new_n249), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n496), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G244), .B(new_n345), .C1(new_n325), .C2(new_n326), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n345), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  OAI211_X1 g0313(.A(G250), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(new_n278), .B1(G257), .B2(new_n486), .ZN(new_n516));
  AOI21_X1  g0316(.A(G169), .B1(new_n516), .B2(new_n484), .ZN(new_n517));
  INV_X1    g0317(.A(G179), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n513), .B(new_n514), .C1(new_n509), .C2(new_n510), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT4), .B1(new_n265), .B2(G244), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n278), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n486), .A2(G257), .ZN(new_n522));
  AND4_X1   g0322(.A1(new_n518), .A2(new_n521), .A3(new_n484), .A4(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  INV_X1    g0325(.A(G97), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n383), .ZN(new_n527));
  NOR2_X1   g0327(.A1(G97), .A2(G107), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n383), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n383), .B1(new_n362), .B2(new_n363), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT75), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(G107), .B1(new_n313), .B2(new_n315), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT75), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n259), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n247), .A2(new_n526), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n462), .B2(new_n526), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n524), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G238), .B(new_n345), .C1(new_n325), .C2(new_n326), .ZN(new_n543));
  OAI211_X1 g0343(.A(G244), .B(G1698), .C1(new_n325), .C2(new_n326), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n543), .B(new_n544), .C1(new_n262), .C2(new_n452), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n278), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT76), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n481), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n245), .A2(KEYINPUT76), .A3(G45), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n548), .A2(new_n286), .A3(G250), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n281), .A2(new_n482), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(new_n552), .A3(new_n518), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(new_n551), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n278), .B2(new_n545), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n555), .B2(G169), .ZN(new_n556));
  INV_X1    g0356(.A(new_n394), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(new_n246), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n462), .A2(new_n394), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n528), .A2(new_n337), .B1(new_n412), .B2(new_n223), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G97), .ZN(new_n562));
  OAI22_X1  g0362(.A1(new_n560), .A2(new_n561), .B1(new_n256), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT77), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n268), .A2(new_n564), .A3(new_n223), .A4(G68), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n223), .B(G68), .C1(new_n325), .C2(new_n326), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT77), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AOI211_X1 g0368(.A(new_n558), .B(new_n559), .C1(new_n568), .C2(new_n249), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n556), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n249), .ZN(new_n571));
  INV_X1    g0371(.A(new_n462), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(G87), .ZN(new_n573));
  INV_X1    g0373(.A(new_n558), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n546), .A2(new_n552), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n295), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n555), .A2(new_n498), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n570), .B1(new_n576), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n532), .B1(new_n537), .B2(KEYINPUT75), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n534), .A2(new_n535), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n249), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n516), .A2(new_n295), .A3(new_n484), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n521), .A2(new_n484), .A3(new_n522), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(G200), .ZN(new_n587));
  INV_X1    g0387(.A(new_n541), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n542), .A2(new_n581), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n268), .A2(G257), .A3(new_n345), .ZN(new_n593));
  INV_X1    g0393(.A(G303), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n268), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n278), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n486), .A2(G270), .B1(new_n483), .B2(new_n281), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n374), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n572), .A2(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n247), .A2(new_n452), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n513), .B(new_n223), .C1(G33), .C2(new_n526), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n452), .A2(G20), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n249), .A2(KEYINPUT78), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT78), .B1(new_n249), .B2(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(KEYINPUT20), .B(new_n603), .C1(new_n605), .C2(new_n606), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n602), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n591), .B1(new_n599), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n613), .A2(KEYINPUT21), .A3(new_n598), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n596), .A2(G179), .A3(new_n597), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n596), .A2(new_n597), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G200), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n618), .B(new_n611), .C1(new_n295), .C2(new_n617), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n612), .A2(new_n614), .A3(new_n616), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n590), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n448), .A2(new_n508), .A3(new_n621), .ZN(G372));
  NAND2_X1  g0422(.A1(new_n575), .A2(KEYINPUT82), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT82), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n571), .A2(new_n624), .A3(new_n574), .A4(new_n573), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n570), .B1(new_n626), .B2(new_n580), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n507), .A2(new_n542), .A3(new_n627), .A4(new_n589), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n614), .A2(new_n612), .A3(new_n616), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n469), .A2(new_n495), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n580), .A2(new_n576), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n556), .A2(new_n569), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT26), .B1(new_n542), .B2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n516), .A2(new_n518), .A3(new_n484), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(G169), .B2(new_n586), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n584), .B2(new_n588), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(new_n640), .A3(new_n627), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n636), .A2(new_n641), .A3(new_n634), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n632), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n447), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(KEYINPUT83), .ZN(new_n645));
  INV_X1    g0445(.A(new_n294), .ZN(new_n646));
  INV_X1    g0446(.A(new_n378), .ZN(new_n647));
  INV_X1    g0447(.A(new_n436), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n391), .A2(new_n401), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n444), .A2(new_n445), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n647), .B1(new_n650), .B2(new_n371), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT84), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n302), .A2(new_n304), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n651), .A2(new_n652), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n645), .A2(new_n646), .A3(new_n656), .ZN(G369));
  XOR2_X1   g0457(.A(KEYINPUT86), .B(G330), .Z(new_n658));
  NAND3_X1  g0458(.A1(new_n245), .A2(new_n223), .A3(G13), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT27), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n663), .A3(G213), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G343), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n620), .B1(new_n611), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n611), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n629), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n658), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n666), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n470), .A2(new_n472), .A3(new_n671), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n508), .A2(new_n672), .B1(new_n496), .B2(new_n666), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n508), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n629), .A2(new_n666), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n675), .A2(new_n677), .B1(new_n630), .B2(new_n666), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n211), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n680), .A2(KEYINPUT87), .A3(G41), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT87), .ZN(new_n682));
  INV_X1    g0482(.A(G41), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n211), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NOR4_X1   g0486(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n226), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n639), .A2(new_n640), .A3(new_n581), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n639), .A2(new_n627), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n634), .B(new_n691), .C1(new_n692), .C2(new_n640), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n614), .A2(new_n612), .A3(new_n616), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n628), .B1(new_n496), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n666), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT29), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n643), .A2(new_n666), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n697), .B1(KEYINPUT29), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n493), .A2(new_n555), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT88), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT88), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n493), .A2(new_n702), .A3(new_n555), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n521), .A2(new_n522), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n615), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n701), .A2(new_n705), .A3(KEYINPUT30), .A4(new_n703), .ZN(new_n709));
  INV_X1    g0509(.A(new_n586), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n555), .A2(G179), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n488), .A3(new_n617), .A4(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n671), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT31), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n713), .A2(new_n716), .A3(new_n671), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n675), .A2(new_n590), .A3(new_n620), .A4(new_n666), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n658), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n699), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n690), .B1(new_n723), .B2(G1), .ZN(G364));
  XOR2_X1   g0524(.A(new_n670), .B(KEYINPUT89), .Z(new_n725));
  NOR2_X1   g0525(.A1(new_n209), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n245), .B1(new_n726), .B2(G45), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n685), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n658), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n667), .A2(new_n669), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n725), .B(new_n730), .C1(new_n731), .C2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n211), .A2(G355), .A3(new_n268), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G116), .B2(new_n211), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n680), .A2(new_n268), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G45), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n738), .B1(new_n739), .B2(new_n227), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n240), .A2(new_n739), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G13), .A2(G33), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n222), .B1(G20), .B2(new_n374), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n729), .B1(new_n742), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n223), .A2(new_n518), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n751), .A2(new_n295), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n295), .A2(new_n498), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n223), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n752), .A2(G322), .B1(G303), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G311), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n750), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n498), .A2(G190), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  OAI221_X1 g0564(.A(new_n757), .B1(new_n758), .B2(new_n760), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G294), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n295), .A2(G179), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n223), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n753), .A2(new_n750), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n327), .B1(new_n766), .B2(new_n768), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n765), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n754), .A2(new_n759), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT92), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n754), .A2(new_n761), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(G329), .B1(G283), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT93), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n777), .A2(G107), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n780), .B(new_n268), .C1(new_n337), .C2(new_n755), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT91), .ZN(new_n782));
  XOR2_X1   g0582(.A(KEYINPUT90), .B(G159), .Z(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n774), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  INV_X1    g0585(.A(new_n760), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G77), .A2(new_n786), .B1(new_n762), .B2(G68), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n752), .A2(G58), .B1(G50), .B2(new_n769), .ZN(new_n788));
  INV_X1    g0588(.A(new_n768), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G97), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n785), .A2(new_n787), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n773), .A2(new_n779), .B1(new_n782), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n749), .B1(new_n792), .B2(new_n746), .ZN(new_n793));
  INV_X1    g0593(.A(new_n745), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n733), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n734), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NOR2_X1   g0597(.A1(new_n666), .A2(new_n400), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n649), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n404), .B2(new_n799), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n404), .A2(new_n666), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n632), .B2(new_n642), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT95), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n802), .B(KEYINPUT95), .C1(new_n632), .C2(new_n642), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n698), .A2(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n730), .B1(new_n807), .B2(new_n722), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n722), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n801), .A2(new_n743), .ZN(new_n811));
  INV_X1    g0611(.A(new_n746), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n744), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n729), .B1(G77), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n752), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n766), .B1(new_n763), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G116), .B2(new_n786), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n755), .A2(new_n383), .B1(new_n776), .B2(new_n337), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n268), .B(new_n819), .C1(G303), .C2(new_n769), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n775), .A2(G311), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n818), .A2(new_n790), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G137), .A2(new_n769), .B1(new_n762), .B2(G150), .ZN(new_n823));
  INV_X1    g0623(.A(G143), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n760), .B2(new_n783), .C1(new_n824), .C2(new_n815), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  NOR2_X1   g0626(.A1(new_n776), .A2(new_n318), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n268), .B1(new_n755), .B2(new_n202), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(G58), .C2(new_n789), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  INV_X1    g0630(.A(new_n775), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n822), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n814), .B1(new_n833), .B2(new_n746), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT94), .Z(new_n835));
  AOI22_X1  g0635(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  NAND2_X1  g0637(.A1(new_n442), .A2(new_n443), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n438), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT97), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n840), .A3(new_n433), .ZN(new_n841));
  OAI21_X1  g0641(.A(KEYINPUT97), .B1(new_n444), .B2(new_n445), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n445), .A2(new_n666), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n648), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n843), .B1(new_n839), .B2(new_n648), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n801), .B1(new_n718), .B2(new_n719), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n333), .A2(new_n375), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n357), .B(new_n308), .C1(new_n324), .C2(new_n332), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT37), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n369), .B2(new_n664), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT98), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT37), .B1(new_n333), .B2(new_n665), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT98), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(new_n851), .A4(new_n852), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n367), .A2(KEYINPUT16), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n308), .B1(new_n332), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n375), .B2(new_n665), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n854), .B1(new_n863), .B2(new_n852), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n665), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n379), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(KEYINPUT38), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n864), .B1(new_n856), .B2(new_n859), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n867), .B1(new_n371), .B2(new_n378), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n870), .A2(KEYINPUT99), .A3(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT99), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n876), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n875), .A2(KEYINPUT100), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT100), .B1(new_n875), .B2(new_n877), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n850), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT40), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT102), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n359), .A2(new_n370), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT101), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT101), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n359), .A2(new_n370), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n378), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n333), .A2(new_n665), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT37), .B1(new_n853), .B2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n887), .A2(new_n889), .B1(new_n860), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n870), .B(new_n882), .C1(new_n891), .C2(KEYINPUT38), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n866), .A2(new_n869), .A3(KEYINPUT102), .A4(KEYINPUT38), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n847), .A2(KEYINPUT40), .A3(new_n848), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n880), .A2(new_n881), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n448), .A2(new_n721), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n731), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n391), .A2(new_n401), .A3(new_n666), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT96), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n805), .B2(new_n806), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n845), .A2(new_n846), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n878), .B2(new_n879), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n875), .A2(new_n877), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT39), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n671), .B1(new_n841), .B2(new_n842), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n892), .A2(new_n911), .A3(new_n893), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n647), .A2(new_n664), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n699), .A2(new_n447), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(new_n646), .A3(new_n656), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n915), .B(new_n917), .Z(new_n918));
  OAI22_X1  g0718(.A1(new_n900), .A2(new_n918), .B1(new_n245), .B2(new_n726), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n918), .B2(new_n900), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n921), .A2(G116), .A3(new_n224), .A4(new_n922), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT36), .Z(new_n924));
  OR3_X1    g0724(.A1(new_n226), .A2(new_n267), .A3(new_n319), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n202), .A2(G68), .ZN(new_n926));
  AOI211_X1 g0726(.A(new_n245), .B(G13), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  OR3_X1    g0727(.A1(new_n920), .A2(new_n924), .A3(new_n927), .ZN(G367));
  NOR2_X1   g0728(.A1(new_n626), .A2(new_n666), .ZN(new_n929));
  MUX2_X1   g0729(.A(new_n627), .B(new_n570), .S(new_n929), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT103), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n671), .B1(new_n539), .B2(new_n541), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n542), .A2(new_n934), .A3(new_n589), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n542), .B2(new_n666), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT104), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n674), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n933), .B(new_n939), .Z(new_n940));
  NAND2_X1  g0740(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n932), .B2(KEYINPUT105), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n938), .A2(new_n496), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n666), .B1(new_n943), .B2(new_n639), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n936), .A2(new_n675), .A3(new_n677), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT42), .Z(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n940), .B(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n685), .B(KEYINPUT41), .Z(new_n949));
  NAND2_X1  g0749(.A1(new_n675), .A2(new_n677), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n673), .B2(new_n677), .ZN(new_n951));
  NOR3_X1   g0751(.A1(new_n951), .A2(new_n658), .A3(new_n732), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n725), .B2(new_n951), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n723), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT106), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT44), .ZN(new_n956));
  OR4_X1    g0756(.A1(new_n955), .A2(new_n678), .A3(new_n956), .A4(new_n936), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n678), .A2(new_n936), .B1(new_n955), .B2(new_n956), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT107), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n674), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n678), .A2(new_n936), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n678), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n966));
  INV_X1    g0766(.A(new_n674), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n965), .A2(new_n966), .B1(new_n967), .B2(KEYINPUT107), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n960), .A2(new_n962), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n962), .B1(new_n960), .B2(new_n968), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n954), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n949), .B1(new_n971), .B2(new_n723), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(KEYINPUT108), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n727), .B1(new_n972), .B2(KEYINPUT108), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n948), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n747), .B1(new_n211), .B2(new_n394), .C1(new_n738), .C2(new_n236), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n730), .B1(KEYINPUT109), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(KEYINPUT109), .B2(new_n976), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n752), .A2(G150), .B1(G143), .B2(new_n769), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n317), .B2(new_n755), .C1(new_n267), .C2(new_n776), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n768), .A2(new_n318), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n268), .B1(new_n763), .B2(new_n783), .ZN(new_n982));
  INV_X1    g0782(.A(G137), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n760), .A2(new_n202), .B1(new_n774), .B2(new_n983), .ZN(new_n984));
  NOR4_X1   g0784(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n774), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G294), .A2(new_n762), .B1(new_n986), .B2(G317), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n758), .B2(new_n770), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n815), .A2(new_n594), .B1(new_n760), .B2(new_n816), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n756), .A2(KEYINPUT46), .A3(G116), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n755), .B2(new_n452), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n992), .C1(new_n383), .C2(new_n768), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n327), .B1(new_n776), .B2(new_n526), .ZN(new_n994));
  NOR4_X1   g0794(.A1(new_n988), .A2(new_n989), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n985), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT47), .Z(new_n997));
  AOI21_X1  g0797(.A(new_n978), .B1(new_n997), .B2(new_n746), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n930), .B2(new_n794), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n975), .A2(new_n999), .ZN(G387));
  NOR2_X1   g0800(.A1(new_n954), .A2(new_n686), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n723), .B2(new_n953), .ZN(new_n1002));
  OR3_X1    g0802(.A1(new_n233), .A2(new_n739), .A3(new_n268), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n255), .A2(G50), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n739), .B1(new_n318), .B2(new_n267), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n327), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n687), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n680), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n747), .B1(new_n383), .B2(new_n211), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n729), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n763), .A2(new_n255), .B1(new_n755), .B2(new_n267), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n327), .B(new_n1013), .C1(G97), .C2(new_n777), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n786), .A2(G68), .B1(new_n769), .B2(G159), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(KEYINPUT111), .B(G150), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n752), .A2(G50), .B1(new_n986), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n789), .A2(new_n557), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1014), .A2(new_n1015), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n789), .A2(G283), .B1(new_n756), .B2(G294), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n752), .A2(G317), .B1(G303), .B2(new_n786), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G322), .A2(new_n769), .B1(new_n762), .B2(G311), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT112), .Z(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1021), .B1(new_n1026), .B2(KEYINPUT48), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT48), .B2(new_n1026), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT49), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n327), .B1(new_n774), .B2(new_n771), .C1(new_n452), .C2(new_n776), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1020), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1012), .B1(new_n1031), .B2(new_n746), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n673), .A2(new_n794), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n953), .A2(new_n728), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1002), .A2(new_n1034), .ZN(G393));
  INV_X1    g0835(.A(new_n970), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n960), .A2(new_n962), .A3(new_n968), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n686), .B1(new_n1038), .B2(new_n954), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n954), .B2(new_n1038), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n728), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n747), .B1(new_n526), .B2(new_n211), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n243), .B2(new_n737), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n789), .A2(G116), .B1(new_n762), .B2(G303), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1044), .A2(KEYINPUT114), .B1(G294), .B2(new_n786), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(KEYINPUT114), .B2(new_n1044), .ZN(new_n1046));
  XOR2_X1   g0846(.A(new_n1046), .B(KEYINPUT115), .Z(new_n1047));
  AOI22_X1  g0847(.A1(new_n752), .A2(G311), .B1(G317), .B2(new_n769), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT52), .Z(new_n1049));
  AOI22_X1  g0849(.A1(G283), .A2(new_n756), .B1(new_n986), .B2(G322), .ZN(new_n1050));
  NAND4_X1  g0850(.A1(new_n1049), .A2(new_n327), .A3(new_n780), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n755), .A2(new_n318), .B1(new_n774), .B2(new_n824), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n327), .B(new_n1052), .C1(G87), .C2(new_n777), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT113), .Z(new_n1054));
  AOI22_X1  g0854(.A1(new_n752), .A2(G159), .B1(G150), .B2(new_n769), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT51), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n789), .A2(G77), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n392), .A2(new_n786), .B1(new_n762), .B2(G50), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n1047), .A2(new_n1051), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n730), .B(new_n1043), .C1(new_n1060), .C2(new_n746), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n937), .B2(new_n794), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1040), .A2(new_n1041), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(G390));
  INV_X1    g0864(.A(KEYINPUT116), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n801), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n717), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n716), .B1(new_n713), .B2(new_n671), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n621), .A2(new_n508), .A3(new_n671), .ZN(new_n1070));
  OAI211_X1 g0870(.A(G330), .B(new_n1066), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(KEYINPUT117), .B1(new_n905), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(G330), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1073), .B(new_n801), .C1(new_n718), .C2(new_n719), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT117), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n1075), .A3(new_n847), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1065), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n803), .A2(new_n804), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n806), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n902), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n847), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n910), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1081), .A2(new_n1082), .B1(new_n909), .B2(new_n912), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n696), .A2(new_n801), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n901), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n847), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n894), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1077), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1082), .B1(new_n904), .B2(new_n905), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n892), .A2(new_n911), .A3(new_n893), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n911), .B1(new_n875), .B2(new_n877), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n894), .A2(new_n1086), .A3(new_n1082), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT116), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n847), .A2(new_n731), .A3(new_n720), .A4(new_n1066), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1092), .B(new_n1093), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1088), .A2(new_n1096), .A3(new_n728), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n743), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n815), .A2(new_n452), .B1(new_n760), .B2(new_n526), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G283), .B2(new_n769), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n327), .B1(new_n755), .B2(new_n337), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n827), .B(new_n1101), .C1(G107), .C2(new_n762), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n775), .A2(G294), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n1057), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n755), .A2(new_n1016), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT53), .ZN(new_n1106));
  INV_X1    g0906(.A(G128), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n268), .B1(new_n770), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G159), .B2(new_n789), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n815), .A2(new_n830), .B1(new_n776), .B2(new_n202), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n763), .A2(new_n983), .B1(new_n760), .B2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n775), .A2(G125), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1106), .A2(new_n1109), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n812), .B1(new_n1104), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT118), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n729), .B1(new_n392), .B2(new_n813), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1098), .B(new_n1119), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1097), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT119), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1097), .A2(KEYINPUT119), .A3(new_n1120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1088), .A2(new_n1096), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n447), .A2(G330), .A3(new_n720), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n916), .A2(new_n1126), .A3(new_n656), .A4(new_n646), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n720), .A2(new_n731), .A3(new_n1066), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n905), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1072), .A2(new_n1076), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n1080), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n905), .A2(new_n1071), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1095), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1127), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n686), .B1(new_n1125), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1088), .A3(new_n1096), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1123), .A2(new_n1124), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(new_n1127), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n298), .A2(new_n665), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT55), .Z(new_n1144));
  XOR2_X1   g0944(.A(new_n305), .B(new_n1144), .Z(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1146));
  XNOR2_X1  g0946(.A(new_n1145), .B(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n892), .A2(new_n893), .ZN(new_n1149));
  OAI21_X1  g0949(.A(G330), .B1(new_n1149), .B2(new_n895), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n880), .B2(new_n881), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1151), .A2(new_n915), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n915), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1148), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1073), .B1(new_n894), .B2(new_n896), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT100), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n908), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n875), .A2(KEYINPUT100), .A3(new_n877), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n849), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1155), .B1(new_n1159), .B2(KEYINPUT40), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n913), .A2(new_n914), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1161), .A3(new_n907), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1151), .A2(new_n915), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1162), .A2(new_n1163), .A3(new_n1147), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1142), .A2(new_n1154), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n686), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1142), .A2(new_n1154), .A3(KEYINPUT57), .A4(new_n1164), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1154), .A2(new_n728), .A3(new_n1164), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n729), .B1(G50), .B2(new_n813), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(G33), .A2(G41), .ZN(new_n1172));
  AOI211_X1 g0972(.A(G50), .B(new_n1172), .C1(new_n327), .C2(new_n683), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n752), .A2(G107), .B1(G58), .B2(new_n777), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n452), .B2(new_n770), .C1(new_n831), .C2(new_n816), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n683), .B(new_n327), .C1(new_n755), .C2(new_n267), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n763), .A2(new_n526), .B1(new_n760), .B2(new_n394), .ZN(new_n1177));
  OR4_X1    g0977(.A1(new_n981), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1173), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n789), .A2(G150), .B1(G125), .B2(new_n769), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT120), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n815), .A2(new_n1107), .B1(new_n760), .B2(new_n983), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n763), .A2(new_n830), .B1(new_n755), .B2(new_n1111), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(G124), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1172), .B1(new_n774), .B2(new_n1189), .C1(new_n783), .C2(new_n776), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1192));
  OAI221_X1 g0992(.A(new_n1180), .B1(new_n1179), .B2(new_n1178), .C1(new_n1188), .C2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1171), .B1(new_n1193), .B2(new_n746), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1147), .B2(new_n744), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1170), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1169), .A2(new_n1197), .ZN(G375));
  OAI21_X1  g0998(.A(new_n729), .B1(G68), .B2(new_n813), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n752), .A2(G137), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n763), .B2(new_n1111), .C1(new_n830), .C2(new_n770), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT123), .Z(new_n1202));
  AOI22_X1  g1002(.A1(G150), .A2(new_n786), .B1(new_n756), .B2(G159), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n327), .B1(new_n777), .B2(G58), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(new_n202), .B2(new_n768), .C1(new_n1107), .C2(new_n831), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G107), .A2(new_n786), .B1(new_n762), .B2(G116), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT122), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n815), .A2(new_n816), .B1(new_n755), .B2(new_n526), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G294), .B2(new_n769), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n775), .A2(G303), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n268), .B1(new_n777), .B2(G77), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1210), .A2(new_n1019), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1202), .A2(new_n1206), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1199), .B1(new_n1214), .B2(new_n746), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n847), .B2(new_n744), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1095), .A2(new_n1133), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1130), .A2(new_n1080), .B1(new_n1217), .B2(new_n1132), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1218), .B2(new_n727), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT124), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OAI211_X1 g1021(.A(KEYINPUT124), .B(new_n1216), .C1(new_n1218), .C2(new_n727), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n949), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1218), .A2(new_n1127), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1136), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(G381));
  AOI21_X1  g1027(.A(new_n1196), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1139), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n975), .A2(new_n1063), .A3(new_n999), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT125), .Z(new_n1232));
  OR4_X1    g1032(.A1(G381), .A2(new_n1229), .A3(new_n1230), .A4(new_n1232), .ZN(G407));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(G343), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT126), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1162), .A2(new_n1163), .A3(new_n1147), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1147), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1238), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1154), .A2(KEYINPUT126), .A3(new_n1164), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1241), .A2(new_n728), .A3(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1142), .A2(new_n1154), .A3(new_n1224), .A4(new_n1164), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1243), .A2(new_n1139), .A3(new_n1195), .A4(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1237), .B(new_n1245), .C1(new_n1228), .C2(new_n1139), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1225), .B1(new_n1135), .B2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1218), .A2(KEYINPUT60), .A3(new_n1127), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1248), .A2(new_n685), .A3(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(new_n1223), .A3(G384), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(G384), .B1(new_n1250), .B2(new_n1223), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT62), .B1(new_n1246), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1250), .A2(new_n1223), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n836), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1236), .A2(G2897), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1258), .A2(new_n1251), .A3(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1258), .B2(new_n1251), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT61), .B1(new_n1246), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G375), .A2(G378), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1139), .A2(new_n1195), .A3(new_n1244), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1236), .B1(new_n1265), .B2(new_n1243), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1266), .A3(new_n1267), .A4(new_n1254), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1256), .A2(new_n1263), .A3(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(new_n796), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1230), .A2(KEYINPUT127), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1063), .B1(new_n975), .B2(new_n999), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1270), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G387), .A2(G390), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1270), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1274), .A2(KEYINPUT127), .A3(new_n1230), .A4(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1269), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1246), .B2(new_n1255), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1264), .A2(new_n1266), .A3(KEYINPUT63), .A4(new_n1254), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1277), .A3(new_n1263), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(new_n1283), .ZN(G405));
  NAND2_X1  g1084(.A1(new_n1264), .A2(new_n1229), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1254), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1264), .A2(new_n1229), .A3(new_n1255), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1286), .A2(new_n1277), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1277), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(G402));
endmodule


