//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n968;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G57gat), .ZN(new_n204));
  INV_X1    g003(.A(G85gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G141gat), .B(G148gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n210), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  INV_X1    g015(.A(G148gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G155gat), .B(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT2), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n214), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G134gat), .ZN(new_n230));
  INV_X1    g029(.A(G120gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G113gat), .ZN(new_n232));
  INV_X1    g031(.A(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n230), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  AOI211_X1 g036(.A(KEYINPUT1), .B(G134gat), .C1(new_n232), .C2(new_n234), .ZN(new_n238));
  OAI21_X1  g037(.A(G127gat), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G134gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G127gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT1), .B1(new_n232), .B2(new_n234), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n241), .B(new_n242), .C1(new_n243), .C2(new_n230), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n228), .A2(new_n239), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n244), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n226), .ZN(new_n249));
  AOI211_X1 g048(.A(KEYINPUT4), .B(new_n225), .C1(new_n239), .C2(new_n244), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n207), .B(new_n246), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n207), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n239), .A2(new_n225), .A3(new_n244), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n225), .B1(new_n239), .B2(new_n244), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n251), .A2(new_n256), .A3(KEYINPUT76), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(KEYINPUT76), .B2(new_n251), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n206), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n251), .A2(KEYINPUT76), .ZN(new_n260));
  INV_X1    g059(.A(new_n256), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n251), .A2(new_n256), .A3(KEYINPUT76), .ZN(new_n263));
  INV_X1    g062(.A(new_n206), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT6), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n259), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n262), .A2(KEYINPUT6), .A3(new_n263), .A4(new_n264), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT35), .ZN(new_n270));
  NAND2_X1  g069(.A1(G211gat), .A2(G218gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT22), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274));
  AND2_X1   g073(.A1(G197gat), .A2(G204gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n273), .B(KEYINPUT73), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT74), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G211gat), .A2(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n271), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT74), .B1(new_n280), .B2(new_n271), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G226gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n292));
  OR2_X1    g091(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n294));
  AOI21_X1  g093(.A(G190gat), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI211_X1 g099(.A(KEYINPUT67), .B(KEYINPUT28), .C1(new_n300), .C2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(G169gat), .ZN(new_n307));
  INV_X1    g106(.A(G176gat), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n305), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n297), .A2(new_n301), .A3(new_n302), .A4(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n302), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT64), .B(KEYINPUT24), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT64), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n302), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(KEYINPUT65), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI22_X1  g119(.A1(KEYINPUT65), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n318), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n323), .A2(new_n321), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n316), .A2(KEYINPUT66), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n328), .A2(new_n302), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n328), .A3(new_n302), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n327), .A2(new_n329), .A3(new_n319), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT25), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n310), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n291), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT25), .B1(new_n314), .B2(new_n317), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n336), .A2(new_n324), .B1(new_n331), .B2(KEYINPUT25), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n290), .B1(new_n337), .B2(new_n310), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n289), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(new_n291), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT29), .B1(new_n337), .B2(new_n310), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n288), .B(new_n340), .C1(new_n341), .C2(new_n291), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G8gat), .B(G36gat), .Z(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G64gat), .ZN(new_n345));
  INV_X1    g144(.A(G92gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(KEYINPUT75), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n339), .A2(new_n342), .A3(new_n347), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n347), .B1(new_n339), .B2(new_n342), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT30), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n269), .A2(new_n270), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT82), .ZN(new_n359));
  XOR2_X1   g158(.A(G78gat), .B(G106gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT31), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(G50gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G228gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n288), .B1(new_n366), .B2(KEYINPUT29), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n283), .A2(new_n334), .A3(new_n225), .A4(new_n287), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n368), .A2(KEYINPUT78), .A3(new_n245), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT78), .B1(new_n368), .B2(new_n245), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n365), .B(new_n367), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT29), .B1(new_n284), .B2(new_n281), .ZN(new_n373));
  INV_X1    g172(.A(new_n274), .ZN(new_n374));
  NAND2_X1  g173(.A1(G197gat), .A2(G204gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n376), .A2(KEYINPUT22), .A3(new_n271), .A4(new_n280), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n372), .B(new_n225), .C1(new_n378), .C2(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT3), .B1(new_n373), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT77), .B1(new_n380), .B2(new_n226), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n367), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n364), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n371), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  INV_X1    g184(.A(G22gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n385), .A2(new_n386), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n384), .A2(KEYINPUT79), .A3(G22gat), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n363), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n386), .A2(KEYINPUT80), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n371), .B2(new_n383), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n371), .A2(new_n383), .A3(new_n394), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n362), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT81), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n389), .B1(new_n384), .B2(new_n387), .ZN(new_n400));
  AOI211_X1 g199(.A(new_n385), .B(new_n386), .C1(new_n371), .C2(new_n383), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n362), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  INV_X1    g202(.A(new_n397), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n363), .B1(new_n404), .B2(new_n395), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n356), .B1(new_n268), .B2(new_n267), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n337), .A2(new_n239), .A3(new_n244), .A4(new_n310), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n333), .A2(new_n248), .ZN(new_n412));
  INV_X1    g211(.A(G227gat), .ZN(new_n413));
  INV_X1    g212(.A(G233gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT69), .ZN(new_n418));
  XNOR2_X1  g217(.A(G15gat), .B(G43gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT70), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(G71gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G99gat), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n416), .A2(new_n425), .A3(KEYINPUT32), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n418), .A2(new_n422), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(KEYINPUT33), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT32), .A3(new_n416), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n411), .A2(new_n412), .ZN(new_n431));
  INV_X1    g230(.A(new_n415), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n427), .A3(new_n429), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n436), .A2(new_n427), .A3(KEYINPUT72), .A4(new_n429), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n359), .A2(new_n407), .A3(new_n410), .A4(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n440), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n436), .B1(new_n427), .B2(new_n429), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n406), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n403), .B1(new_n402), .B2(new_n405), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n447), .B(new_n408), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n444), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n441), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n447), .A2(KEYINPUT36), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n269), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n399), .B(new_n406), .C1(new_n457), .C2(new_n356), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n253), .A2(new_n254), .A3(new_n252), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n246), .B1(new_n249), .B2(new_n250), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n252), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT39), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n463), .A3(new_n252), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n206), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT40), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n466), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n467), .A2(new_n265), .A3(new_n356), .A4(new_n468), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n343), .A2(KEYINPUT37), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n343), .A2(KEYINPUT37), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n347), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n472), .A2(KEYINPUT38), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(KEYINPUT38), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n475), .A2(new_n268), .A3(new_n267), .A4(new_n349), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n469), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n407), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n456), .B(new_n458), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n452), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT83), .ZN(new_n481));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(G197gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT11), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(new_n307), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n485), .B(KEYINPUT12), .Z(new_n486));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT13), .Z(new_n488));
  XOR2_X1   g287(.A(G15gat), .B(G22gat), .Z(new_n489));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n490));
  INV_X1    g289(.A(G1gat), .ZN(new_n491));
  OR3_X1    g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n489), .B2(new_n490), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n492), .B(new_n493), .C1(KEYINPUT16), .C2(new_n489), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(G50gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G43gat), .ZN(new_n498));
  INV_X1    g297(.A(G43gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(G50gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT15), .ZN(new_n501));
  INV_X1    g300(.A(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n503), .A3(KEYINPUT14), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT14), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n505), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G29gat), .A2(G36gat), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n498), .A2(new_n500), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n509), .B(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n508), .A2(new_n513), .A3(new_n501), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT85), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT15), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n518), .A2(new_n507), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT85), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n519), .A2(new_n520), .A3(new_n513), .A4(new_n515), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n510), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n496), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n494), .B(G8gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n517), .A2(new_n521), .ZN(new_n525));
  INV_X1    g324(.A(new_n510), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n488), .B1(new_n523), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT17), .B1(new_n527), .B2(KEYINPUT86), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT86), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n522), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n496), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n524), .A2(new_n527), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(new_n487), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(KEYINPUT88), .A3(KEYINPUT18), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n536), .A2(new_n537), .A3(new_n487), .A4(new_n540), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n486), .B(new_n531), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n486), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n541), .ZN(new_n544));
  INV_X1    g343(.A(new_n531), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n452), .A2(new_n479), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n481), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT89), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT97), .ZN(new_n553));
  INV_X1    g352(.A(G99gat), .ZN(new_n554));
  INV_X1    g353(.A(G106gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n560), .A2(KEYINPUT101), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT7), .ZN(new_n563));
  AOI22_X1  g362(.A1(KEYINPUT8), .A2(new_n558), .B1(new_n205), .B2(new_n346), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(KEYINPUT101), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n561), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT98), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(new_n560), .B2(new_n565), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n559), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT98), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT92), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT9), .ZN(new_n576));
  OR2_X1    g375(.A1(G71gat), .A2(G78gat), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G57gat), .B(G64gat), .Z(new_n579));
  INV_X1    g378(.A(KEYINPUT9), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n575), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT93), .A4(new_n582), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT90), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n574), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(KEYINPUT90), .A2(G71gat), .A3(G78gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n579), .A2(new_n581), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n577), .B(KEYINPUT91), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n585), .A2(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n567), .A2(new_n573), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n570), .A2(new_n571), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n573), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n585), .A2(new_n586), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n591), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT100), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n594), .B1(new_n569), .B2(new_n572), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n601), .A2(new_n602), .A3(new_n592), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n593), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT102), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n610), .B(new_n593), .C1(new_n600), .C2(new_n603), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n599), .B(KEYINPUT96), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n601), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n605), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(new_n308), .ZN(new_n617));
  INV_X1    g416(.A(G204gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n607), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n609), .A2(new_n615), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n606), .B1(new_n611), .B2(new_n613), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n619), .B1(new_n608), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT89), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n481), .A2(new_n628), .A3(new_n547), .A4(new_n549), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n551), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n612), .A2(KEYINPUT21), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n496), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(new_n242), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n634), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n636), .A3(new_n496), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n639));
  XNOR2_X1  g438(.A(G183gat), .B(G211gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n639), .B(new_n640), .Z(new_n641));
  OR2_X1    g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n638), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n645));
  NOR2_X1   g444(.A1(new_n592), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT95), .B(G155gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n648), .A3(new_n643), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n532), .A2(new_n535), .ZN(new_n653));
  AND2_X1   g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n653), .A2(new_n596), .B1(KEYINPUT41), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n527), .A2(new_n601), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(G190gat), .B(G218gat), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n655), .A2(new_n658), .A3(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n654), .A2(KEYINPUT41), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G134gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(new_n222), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n666), .B2(KEYINPUT99), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n660), .A2(KEYINPUT99), .A3(new_n661), .A4(new_n665), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n652), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n630), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n269), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(new_n491), .ZN(G1324gat));
  NOR2_X1   g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n672), .A2(new_n357), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n679));
  INV_X1    g478(.A(new_n672), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n495), .B1(new_n680), .B2(new_n356), .ZN(new_n681));
  OAI21_X1  g480(.A(KEYINPUT42), .B1(new_n681), .B2(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(G1325gat));
  INV_X1    g482(.A(new_n456), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n680), .A2(G15gat), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(G15gat), .B1(new_n680), .B2(new_n443), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(G1326gat));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n407), .ZN(new_n688));
  XOR2_X1   g487(.A(KEYINPUT43), .B(G22gat), .Z(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  NAND3_X1  g489(.A1(new_n481), .A2(new_n670), .A3(new_n549), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT44), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n480), .A2(new_n670), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(KEYINPUT44), .B2(new_n691), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n694), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n626), .B(KEYINPUT103), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n652), .A3(new_n547), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  OR3_X1    g501(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n269), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT106), .B1(new_n702), .B2(new_n269), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(G29gat), .A3(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n551), .A2(new_n670), .A3(new_n627), .A4(new_n629), .ZN(new_n706));
  INV_X1    g505(.A(new_n652), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n502), .A3(new_n457), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(new_n710), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n503), .A3(new_n356), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT46), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n702), .B2(new_n357), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(KEYINPUT46), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(G1329gat));
  INV_X1    g515(.A(new_n696), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n693), .B1(new_n692), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT105), .B1(new_n691), .B2(KEYINPUT44), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n684), .B(new_n701), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G43gat), .ZN(new_n721));
  INV_X1    g520(.A(new_n443), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(G43gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT47), .B1(new_n725), .B2(KEYINPUT107), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n720), .A2(G43gat), .B1(new_n708), .B2(new_n723), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n726), .A2(new_n730), .ZN(G1330gat));
  NAND3_X1  g530(.A1(new_n698), .A2(new_n478), .A3(new_n701), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G50gat), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n708), .A2(new_n497), .A3(new_n478), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n698), .A2(KEYINPUT108), .A3(new_n478), .A4(new_n701), .ZN(new_n740));
  AND3_X1   g539(.A1(new_n739), .A2(G50gat), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n734), .A2(KEYINPUT48), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n737), .B1(new_n741), .B2(new_n742), .ZN(G1331gat));
  INV_X1    g542(.A(new_n699), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n652), .A2(new_n670), .A3(new_n547), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n480), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n457), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n356), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  NAND2_X1  g552(.A1(new_n746), .A2(new_n443), .ZN(new_n754));
  INV_X1    g553(.A(G71gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n746), .A2(G71gat), .A3(new_n684), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(KEYINPUT110), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(new_n760), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(KEYINPUT109), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n759), .A2(new_n764), .A3(new_n761), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n763), .A2(KEYINPUT50), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT50), .B1(new_n763), .B2(new_n765), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n746), .A2(new_n478), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g569(.A1(new_n707), .A2(new_n547), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n698), .A2(new_n626), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n269), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n480), .A2(new_n670), .A3(new_n771), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT51), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n627), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(new_n205), .A3(new_n457), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n773), .A2(new_n777), .ZN(G1336gat));
  NAND4_X1  g577(.A1(new_n698), .A2(new_n626), .A3(new_n356), .A4(new_n771), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G92gat), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n775), .A2(new_n699), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n346), .A3(new_n356), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n780), .A2(new_n785), .A3(new_n782), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(G1337gat));
  NAND4_X1  g586(.A1(new_n698), .A2(new_n626), .A3(new_n684), .A4(new_n771), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G99gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n776), .A2(new_n554), .A3(new_n443), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(KEYINPUT111), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(G1338gat));
  NAND4_X1  g594(.A1(new_n698), .A2(new_n626), .A3(new_n478), .A4(new_n771), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT112), .B(G106gat), .Z(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n555), .A3(new_n478), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT53), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n802), .A3(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n801), .A2(new_n803), .ZN(G1339gat));
  NAND3_X1  g603(.A1(new_n611), .A2(new_n606), .A3(new_n613), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n615), .A2(KEYINPUT54), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n620), .B1(new_n624), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(KEYINPUT55), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n623), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n614), .A2(new_n807), .A3(new_n605), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n805), .A2(KEYINPUT54), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n619), .B(new_n812), .C1(new_n813), .C2(new_n624), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n547), .A2(new_n811), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n544), .A2(new_n543), .A3(new_n545), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n487), .B1(new_n536), .B2(new_n537), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n523), .A2(new_n528), .A3(new_n488), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n485), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n626), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n670), .B1(new_n817), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n811), .A2(new_n823), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n668), .A2(new_n669), .A3(new_n816), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n652), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n745), .A2(new_n627), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n407), .A2(new_n447), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n269), .A2(new_n356), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n233), .A3(new_n547), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n831), .B2(new_n407), .ZN(new_n838));
  AOI211_X1 g637(.A(KEYINPUT113), .B(new_n478), .C1(new_n829), .C2(new_n830), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n722), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n834), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n829), .A2(new_n830), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT113), .B1(new_n843), .B2(new_n478), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n831), .A2(new_n837), .A3(new_n407), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n844), .A2(new_n443), .A3(new_n834), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT114), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n842), .A2(new_n847), .A3(new_n547), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n836), .B1(new_n848), .B2(new_n233), .ZN(G1340gat));
  NAND3_X1  g648(.A1(new_n835), .A2(new_n231), .A3(new_n626), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n842), .A2(new_n847), .A3(new_n744), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n231), .ZN(G1341gat));
  XOR2_X1   g651(.A(KEYINPUT68), .B(G127gat), .Z(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n835), .A2(new_n707), .A3(new_n854), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n842), .A2(new_n847), .A3(new_n707), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n854), .ZN(G1342gat));
  NAND2_X1  g656(.A1(new_n670), .A2(new_n357), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n858), .B(KEYINPUT115), .Z(new_n859));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n269), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n240), .A3(new_n832), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT56), .Z(new_n862));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n847), .A3(new_n670), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(KEYINPUT116), .A3(G134gat), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT116), .B1(new_n863), .B2(G134gat), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(G1343gat));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n831), .A2(new_n867), .A3(new_n478), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n456), .A2(new_n834), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  XOR2_X1   g669(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n806), .B2(new_n808), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT118), .B1(new_n810), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n814), .A2(new_n871), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n623), .A4(new_n809), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n874), .A2(new_n547), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n670), .B1(new_n878), .B2(new_n824), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n652), .B1(new_n879), .B2(new_n828), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n407), .B1(new_n880), .B2(new_n830), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n868), .B(new_n870), .C1(new_n881), .C2(new_n867), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n542), .A2(new_n546), .ZN(new_n883));
  OAI21_X1  g682(.A(G141gat), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT58), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n843), .A2(new_n407), .A3(new_n869), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n215), .A3(new_n547), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n886), .B(new_n889), .Z(G1344gat));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n217), .A3(new_n626), .ZN(new_n891));
  XOR2_X1   g690(.A(new_n891), .B(KEYINPUT120), .Z(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT122), .B1(new_n881), .B2(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n745), .A2(new_n627), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n627), .A2(new_n822), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n875), .A2(new_n623), .A3(new_n809), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n883), .B1(new_n898), .B2(KEYINPUT118), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n899), .B2(new_n877), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n900), .A2(new_n670), .B1(new_n827), .B2(new_n826), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(new_n652), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n895), .B(new_n867), .C1(new_n902), .C2(new_n407), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n831), .A2(KEYINPUT57), .A3(new_n478), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n894), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n870), .A2(KEYINPUT121), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n870), .A2(KEYINPUT121), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n627), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n217), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n905), .A2(KEYINPUT123), .A3(new_n908), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n893), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n893), .B(G148gat), .C1(new_n882), .C2(new_n627), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n892), .B1(new_n913), .B2(new_n915), .ZN(G1345gat));
  OAI21_X1  g715(.A(G155gat), .B1(new_n882), .B2(new_n652), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n887), .A2(new_n221), .A3(new_n707), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(G1346gat));
  INV_X1    g718(.A(new_n670), .ZN(new_n920));
  OAI21_X1  g719(.A(G162gat), .B1(new_n882), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n684), .A2(new_n407), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n860), .A2(new_n222), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n457), .A2(new_n357), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n833), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n307), .A3(new_n547), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n840), .A2(new_n547), .A3(new_n925), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT124), .B1(new_n929), .B2(G169gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  NAND4_X1  g732(.A1(new_n844), .A2(new_n443), .A3(new_n845), .A4(new_n925), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n934), .A2(new_n308), .A3(new_n699), .ZN(new_n935));
  AOI21_X1  g734(.A(G176gat), .B1(new_n927), .B2(new_n626), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  NOR2_X1   g736(.A1(new_n926), .A2(new_n300), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT125), .B1(new_n938), .B2(new_n707), .ZN(new_n939));
  OAI21_X1  g738(.A(G183gat), .B1(new_n934), .B2(new_n652), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  OR3_X1    g741(.A1(new_n926), .A2(G190gat), .A3(new_n920), .ZN(new_n943));
  OAI21_X1  g742(.A(G190gat), .B1(new_n934), .B2(new_n920), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1351gat));
  AND3_X1   g747(.A1(new_n831), .A2(new_n922), .A3(new_n925), .ZN(new_n949));
  INV_X1    g748(.A(G197gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n950), .A3(new_n547), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT126), .Z(new_n952));
  AND4_X1   g751(.A1(new_n547), .A2(new_n905), .A3(new_n456), .A4(new_n925), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n950), .ZN(G1352gat));
  NAND3_X1  g753(.A1(new_n949), .A2(new_n618), .A3(new_n626), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT62), .Z(new_n956));
  AND4_X1   g755(.A1(new_n456), .A2(new_n905), .A3(new_n744), .A4(new_n925), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n618), .ZN(G1353gat));
  INV_X1    g757(.A(G211gat), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n949), .A2(new_n959), .A3(new_n707), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n905), .A2(new_n707), .A3(new_n456), .A4(new_n925), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  AOI21_X1  g763(.A(G218gat), .B1(new_n949), .B2(new_n670), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n905), .A2(new_n456), .A3(new_n925), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n670), .A2(G218gat), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1355gat));
endmodule


