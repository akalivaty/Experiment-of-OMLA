//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT5), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT5), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n188), .A2(G113), .A3(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT2), .B(G113), .Z(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(new_n187), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT83), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT3), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n196), .A2(G104), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n202), .A2(new_n196), .A3(KEYINPUT83), .A4(G104), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n198), .A2(new_n200), .A3(new_n201), .A4(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  OAI21_X1  g020(.A(G101), .B1(new_n199), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n195), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n209), .B(KEYINPUT88), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n195), .A2(new_n208), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g026(.A(G110), .B(G122), .Z(new_n213));
  XOR2_X1   g027(.A(new_n213), .B(KEYINPUT8), .Z(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n223), .A2(KEYINPUT64), .A3(G146), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT64), .B1(new_n223), .B2(G146), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n222), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n223), .A2(G146), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n231));
  OAI21_X1  g045(.A(G128), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n220), .A2(new_n226), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G125), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  OR2_X1    g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n216), .A2(KEYINPUT0), .A3(G128), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n235), .B1(new_n240), .B2(new_n234), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G224), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT7), .ZN(new_n244));
  XOR2_X1   g058(.A(new_n241), .B(new_n244), .Z(new_n245));
  NAND3_X1  g059(.A1(new_n198), .A2(new_n200), .A3(new_n203), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G101), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT4), .A4(new_n204), .ZN(new_n249));
  OR2_X1    g063(.A1(new_n193), .A2(new_n187), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n194), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(G101), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n249), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n213), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n211), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n215), .A2(new_n245), .A3(new_n256), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n241), .B(new_n243), .Z(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n211), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n213), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT6), .A3(new_n256), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n259), .A2(new_n262), .A3(new_n213), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n258), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n257), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(G210), .B1(G237), .B2(G902), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT89), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n268), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n257), .A2(new_n264), .A3(new_n265), .A4(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(KEYINPUT90), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G214), .B1(G237), .B2(G902), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT90), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n266), .A2(new_n274), .A3(new_n268), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT13), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n218), .B2(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT93), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n223), .A2(G128), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(new_n277), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n279), .B(new_n282), .C1(G128), .C2(new_n223), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n280), .A2(new_n277), .ZN(new_n286));
  OAI21_X1  g100(.A(G134), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G122), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(G116), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n288), .A2(G116), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(new_n196), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n218), .A2(G143), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n280), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT95), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n296), .A2(G134), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n287), .A2(new_n293), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT14), .B1(new_n288), .B2(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT96), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT96), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n301), .B(KEYINPUT14), .C1(new_n288), .C2(G116), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n291), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT97), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g119(.A1(new_n290), .A2(KEYINPUT14), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n300), .A2(KEYINPUT97), .A3(new_n291), .A4(new_n302), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G107), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT98), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n296), .B(G134), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n292), .A2(new_n196), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT98), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(new_n313), .A3(G107), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n310), .A2(new_n311), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n298), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT9), .B(G234), .Z(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G217), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n318), .A2(new_n319), .A3(G953), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT99), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n298), .A2(new_n315), .A3(new_n320), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n316), .A2(KEYINPUT99), .A3(new_n321), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n265), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G478), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT15), .ZN(new_n329));
  XOR2_X1   g143(.A(new_n327), .B(new_n329), .Z(new_n330));
  NAND2_X1  g144(.A1(new_n242), .A2(G952), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(G234), .B2(G237), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT21), .B(G898), .Z(new_n334));
  NAND2_X1  g148(.A1(G234), .A2(G237), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(G902), .A3(G953), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G237), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n242), .A3(G214), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(new_n223), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G131), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n339), .B(G143), .ZN(new_n342));
  INV_X1    g156(.A(G131), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G125), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT16), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n234), .A2(KEYINPUT77), .A3(G140), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n234), .A2(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n346), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n350), .B2(KEYINPUT77), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n347), .B1(new_n351), .B2(KEYINPUT16), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n341), .A2(new_n344), .B1(new_n352), .B2(G146), .ZN(new_n353));
  INV_X1    g167(.A(new_n351), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT19), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n350), .B2(KEYINPUT19), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT19), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n351), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n359), .A3(new_n221), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n349), .A2(new_n346), .A3(new_n221), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n351), .B2(new_n221), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT18), .A2(G131), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n342), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n342), .A2(new_n343), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT18), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n353), .A2(new_n360), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(G113), .B(G122), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(new_n205), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT92), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n362), .A3(new_n364), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n356), .A2(new_n359), .A3(new_n221), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n341), .A2(new_n344), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n352), .A2(G146), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n372), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n378));
  INV_X1    g192(.A(new_n370), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n352), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT78), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(new_n221), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT78), .B1(new_n352), .B2(G146), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n375), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT17), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n341), .A2(new_n344), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n366), .A2(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n370), .B(new_n372), .C1(new_n385), .C2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n371), .A2(new_n380), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G475), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n265), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n387), .A2(new_n388), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n396), .A2(new_n375), .A3(new_n384), .A4(new_n383), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n370), .B1(new_n397), .B2(new_n372), .ZN(new_n398));
  INV_X1    g212(.A(new_n390), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n265), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G475), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n391), .A2(KEYINPUT20), .A3(new_n392), .A4(new_n265), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n395), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n330), .A2(new_n337), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT100), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n327), .B(new_n329), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n403), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT100), .A3(new_n337), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n276), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n240), .A2(new_n249), .A3(new_n253), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n217), .B1(new_n216), .B2(new_n219), .ZN(new_n414));
  AND4_X1   g228(.A1(new_n217), .A2(new_n219), .A3(new_n222), .A4(new_n224), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT64), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n221), .B2(G143), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n223), .A2(KEYINPUT64), .A3(G146), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n230), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n218), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n420));
  OAI22_X1  g234(.A1(new_n414), .A2(new_n415), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n421), .A2(KEYINPUT10), .A3(new_n204), .A4(new_n207), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT11), .A2(G134), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(KEYINPUT65), .A2(G137), .ZN(new_n425));
  NOR2_X1   g239(.A1(KEYINPUT65), .A2(G137), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(KEYINPUT11), .A2(G134), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n423), .B1(new_n428), .B2(G137), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n343), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n343), .B1(new_n427), .B2(new_n429), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n434));
  INV_X1    g248(.A(new_n216), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n226), .A2(new_n220), .B1(new_n435), .B2(new_n232), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n436), .B2(new_n208), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n413), .A2(new_n422), .A3(new_n433), .A4(new_n437), .ZN(new_n438));
  XOR2_X1   g252(.A(G110), .B(G140), .Z(new_n439));
  AND2_X1   g253(.A1(new_n242), .A2(G227), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT85), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n233), .A2(new_n208), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n436), .A2(new_n208), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n233), .A2(new_n208), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n449), .B(KEYINPUT85), .C1(new_n208), .C2(new_n436), .ZN(new_n450));
  INV_X1    g264(.A(new_n433), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT12), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(KEYINPUT86), .A3(new_n453), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT12), .B(new_n451), .C1(new_n446), .C2(new_n447), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n444), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n413), .A2(new_n437), .A3(new_n422), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n451), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n441), .B1(new_n462), .B2(new_n438), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n412), .B(new_n265), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(G469), .A2(G902), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n438), .A3(new_n441), .ZN(new_n466));
  INV_X1    g280(.A(new_n438), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n458), .B2(new_n459), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n468), .B2(new_n441), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n464), .B(new_n465), .C1(new_n469), .C2(new_n412), .ZN(new_n470));
  OAI21_X1  g284(.A(G221), .B1(new_n318), .B2(G902), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT82), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n411), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT79), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n478), .B(KEYINPUT22), .Z(new_n479));
  XOR2_X1   g293(.A(new_n479), .B(G137), .Z(new_n480));
  OR3_X1    g294(.A1(new_n218), .A2(KEYINPUT75), .A3(G119), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT75), .B1(new_n218), .B2(G119), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n190), .B2(G128), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n218), .A2(KEYINPUT74), .A3(G119), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n481), .A2(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g300(.A(KEYINPUT24), .B(G110), .Z(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT23), .B1(new_n218), .B2(G119), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT76), .B1(new_n218), .B2(G119), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G110), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n385), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  OAI22_X1  g307(.A1(new_n491), .A2(G110), .B1(new_n486), .B2(new_n487), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n375), .A2(new_n494), .A3(new_n361), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n493), .A2(KEYINPUT80), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT80), .B1(new_n493), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n480), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n497), .A2(new_n480), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n319), .B1(G234), .B2(new_n265), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g317(.A1(new_n503), .A2(KEYINPUT81), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n499), .A3(new_n265), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT25), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n498), .A2(new_n499), .A3(new_n507), .A4(new_n265), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n503), .A2(KEYINPUT81), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(G134), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n425), .B2(new_n426), .ZN(new_n513));
  NAND2_X1  g327(.A1(G134), .A2(G137), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(G131), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n430), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT67), .B1(new_n233), .B2(new_n516), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n430), .A2(new_n515), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n421), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n238), .B(new_n239), .C1(new_n431), .C2(new_n432), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT68), .ZN(new_n525));
  OR3_X1    g339(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n516), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n518), .A2(new_n421), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT69), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT30), .A4(new_n521), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT68), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n530), .A3(new_n523), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n525), .A2(new_n251), .A3(new_n529), .A4(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n251), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n526), .A2(new_n528), .A3(new_n533), .A4(new_n521), .ZN(new_n534));
  NOR2_X1   g348(.A1(G237), .A2(G953), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G210), .ZN(new_n536));
  XOR2_X1   g350(.A(new_n536), .B(KEYINPUT27), .Z(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT26), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(new_n201), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n532), .A2(new_n534), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT31), .ZN(new_n541));
  INV_X1    g355(.A(new_n539), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n527), .A2(new_n521), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT70), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n527), .A2(new_n521), .A3(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n533), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n522), .A2(new_n251), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n548), .B1(new_n551), .B2(new_n534), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n542), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT31), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n532), .A2(new_n554), .A3(new_n534), .A4(new_n539), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n541), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(G472), .A2(G902), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT71), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(KEYINPUT32), .A3(new_n558), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n550), .A2(new_n552), .A3(new_n542), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n539), .B1(new_n532), .B2(new_n534), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT29), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n549), .A2(KEYINPUT72), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n547), .A2(new_n567), .A3(new_n548), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n526), .A2(new_n528), .A3(new_n521), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n251), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n534), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n566), .B(new_n568), .C1(new_n572), .C2(new_n548), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n539), .A2(KEYINPUT29), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n265), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(G472), .B1(new_n565), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n561), .A2(new_n562), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT73), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n561), .A2(new_n576), .A3(new_n579), .A4(new_n562), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n511), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n476), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(KEYINPUT101), .B(G101), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G3));
  INV_X1    g399(.A(G472), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n556), .B2(new_n265), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n558), .B2(new_n556), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n589), .A2(new_n474), .A3(new_n511), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n325), .A2(new_n591), .A3(new_n326), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n322), .A2(KEYINPUT33), .A3(new_n324), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n328), .A2(G902), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n327), .A2(new_n328), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n403), .ZN(new_n598));
  INV_X1    g412(.A(new_n337), .ZN(new_n599));
  INV_X1    g413(.A(new_n273), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n269), .B2(new_n271), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n590), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT34), .B(G104), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  NAND2_X1  g420(.A1(new_n408), .A2(new_n404), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n607), .A2(new_n599), .A3(new_n602), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n590), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NOR2_X1   g425(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n493), .A2(new_n495), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n502), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n509), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n411), .A2(new_n475), .A3(new_n588), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(KEYINPUT37), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G110), .ZN(G12));
  AOI21_X1  g433(.A(new_n474), .B1(new_n578), .B2(new_n580), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n332), .B(KEYINPUT102), .Z(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(G900), .B2(new_n336), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n607), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n602), .B1(new_n509), .B2(new_n615), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n620), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G128), .ZN(G30));
  NAND2_X1  g442(.A1(new_n272), .A2(new_n275), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT38), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n623), .B(KEYINPUT39), .Z(new_n631));
  OR2_X1    g445(.A1(new_n474), .A2(new_n631), .ZN(new_n632));
  AOI211_X1 g446(.A(new_n600), .B(new_n630), .C1(new_n632), .C2(KEYINPUT40), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n330), .A2(new_n404), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n632), .A2(KEYINPUT40), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n561), .A2(new_n562), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n532), .A2(new_n534), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n539), .ZN(new_n638));
  AOI21_X1  g452(.A(G902), .B1(new_n572), .B2(new_n542), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n586), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n616), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n633), .A2(new_n634), .A3(new_n635), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G143), .ZN(G45));
  NAND3_X1  g459(.A1(new_n597), .A2(new_n403), .A3(new_n623), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT103), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n597), .A2(KEYINPUT103), .A3(new_n403), .A4(new_n623), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n601), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n642), .B1(new_n650), .B2(KEYINPUT104), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n648), .A2(new_n652), .A3(new_n601), .A4(new_n649), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n651), .A2(new_n620), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G146), .ZN(G48));
  NAND2_X1  g469(.A1(new_n578), .A2(new_n580), .ZN(new_n656));
  INV_X1    g470(.A(new_n511), .ZN(new_n657));
  INV_X1    g471(.A(new_n444), .ZN(new_n658));
  INV_X1    g472(.A(new_n457), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT86), .B1(new_n452), .B2(new_n453), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n459), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n463), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G469), .B1(new_n662), .B2(G902), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n663), .A2(new_n464), .A3(new_n473), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n656), .A2(new_n657), .A3(new_n603), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT105), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n581), .A2(new_n667), .A3(new_n603), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT41), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G113), .ZN(G15));
  NAND4_X1  g485(.A1(new_n656), .A2(new_n657), .A3(new_n608), .A4(new_n664), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n581), .A2(KEYINPUT106), .A3(new_n608), .A4(new_n664), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  NAND2_X1  g491(.A1(new_n407), .A2(new_n410), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n626), .A2(new_n664), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n678), .A2(new_n656), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n190), .ZN(G21));
  NAND2_X1  g495(.A1(new_n573), .A2(new_n542), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n541), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT107), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n685), .A3(new_n541), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n684), .A2(new_n555), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n587), .B1(new_n687), .B2(new_n558), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n657), .A2(new_n688), .A3(new_n664), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n634), .A2(new_n601), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n689), .A2(new_n599), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n288), .ZN(G24));
  AND2_X1   g506(.A1(new_n648), .A2(new_n649), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n679), .A3(new_n688), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G125), .ZN(G27));
  NAND2_X1  g509(.A1(new_n636), .A2(KEYINPUT108), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n561), .A2(new_n697), .A3(new_n562), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n576), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n629), .A2(new_n273), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n474), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n699), .A2(new_n693), .A3(new_n701), .A4(new_n657), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT42), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT42), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n581), .A2(new_n704), .A3(new_n693), .A4(new_n701), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n343), .ZN(G33));
  NAND3_X1  g521(.A1(new_n581), .A2(new_n625), .A3(new_n701), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n597), .A2(new_n710), .A3(new_n404), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n403), .B(KEYINPUT109), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(new_n597), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n711), .B1(new_n713), .B2(new_n710), .ZN(new_n714));
  OR3_X1    g528(.A1(new_n714), .A2(new_n588), .A3(new_n642), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n700), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n469), .B(KEYINPUT45), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(KEYINPUT46), .A3(new_n465), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n722), .B(G469), .C1(new_n719), .C2(G902), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n464), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n473), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n631), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n715), .A2(new_n716), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n717), .A2(new_n718), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G137), .ZN(G39));
  OR2_X1    g543(.A1(new_n725), .A2(KEYINPUT47), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n656), .A2(new_n657), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n725), .A2(KEYINPUT47), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n693), .A2(new_n718), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n731), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G140), .ZN(G42));
  NAND4_X1  g549(.A1(new_n713), .A2(new_n657), .A3(new_n473), .A4(new_n273), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT110), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n663), .A2(new_n464), .ZN(new_n738));
  OR2_X1    g552(.A1(new_n738), .A2(KEYINPUT49), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n641), .B1(KEYINPUT49), .B2(new_n738), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n737), .A2(new_n630), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n742));
  INV_X1    g556(.A(new_n276), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n607), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n408), .A2(KEYINPUT112), .A3(new_n404), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n598), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n590), .A2(new_n337), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n617), .B(new_n748), .C1(new_n582), .C2(new_n476), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n703), .A2(new_n705), .A3(new_n708), .ZN(new_n750));
  INV_X1    g564(.A(new_n701), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n656), .A2(new_n409), .A3(new_n623), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n693), .A2(new_n688), .ZN(new_n753));
  AOI211_X1 g567(.A(new_n642), .B(new_n751), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n749), .A2(new_n750), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n691), .B1(new_n666), .B2(new_n668), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n680), .B1(new_n674), .B2(new_n675), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n758), .B1(new_n756), .B2(new_n757), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n690), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n474), .A2(new_n624), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n642), .A3(new_n641), .A4(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n654), .A2(new_n627), .A3(new_n694), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n693), .A2(new_n679), .A3(new_n688), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n656), .A2(new_n475), .A3(new_n653), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n651), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(KEYINPUT52), .A3(new_n627), .A4(new_n764), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n765), .A2(new_n767), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n774), .B2(new_n766), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n742), .B1(new_n761), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT114), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n755), .B(new_n774), .C1(new_n759), .C2(new_n760), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(new_n742), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n780), .B(new_n742), .C1(new_n761), .C2(new_n775), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n777), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT54), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n756), .A2(new_n757), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n755), .A2(KEYINPUT53), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n775), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n778), .A2(KEYINPUT115), .A3(new_n742), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT115), .B1(new_n778), .B2(new_n742), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n783), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n784), .B1(new_n783), .B2(new_n791), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n718), .A2(new_n664), .ZN(new_n794));
  OR4_X1    g608(.A1(new_n511), .A2(new_n641), .A3(new_n794), .A4(new_n333), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(new_n598), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n699), .A2(new_n657), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n714), .A2(new_n622), .ZN(new_n799));
  INV_X1    g613(.A(new_n794), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n714), .A2(KEYINPUT117), .A3(new_n622), .A4(new_n794), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT48), .Z(new_n804));
  NOR3_X1   g618(.A1(new_n714), .A2(new_n689), .A3(new_n622), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n331), .B(new_n804), .C1(new_n601), .C2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n616), .B(new_n688), .C1(new_n801), .C2(new_n802), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n807), .B(KEYINPUT118), .Z(new_n808));
  NAND2_X1  g622(.A1(new_n730), .A2(new_n732), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n809), .B1(new_n473), .B2(new_n738), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n657), .A2(new_n688), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(new_n718), .A4(new_n799), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n805), .A2(new_n600), .A3(new_n630), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT50), .Z(new_n814));
  OR3_X1    g628(.A1(new_n795), .A2(new_n403), .A3(new_n597), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n808), .A2(new_n812), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n812), .A2(new_n817), .A3(new_n814), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n816), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n816), .B1(KEYINPUT51), .B2(new_n818), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n796), .B(new_n806), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n792), .A2(new_n793), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(G952), .A2(G953), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n741), .B1(new_n822), .B2(new_n823), .ZN(G75));
  XNOR2_X1  g638(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n787), .B1(new_n789), .B2(new_n790), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(G902), .A3(new_n268), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n261), .A2(new_n263), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(new_n258), .Z(new_n831));
  AND3_X1   g645(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n831), .B1(new_n828), .B2(new_n829), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n826), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n828), .A2(new_n829), .ZN(new_n835));
  INV_X1    g649(.A(new_n831), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n825), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n242), .A2(G952), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(G51));
  XOR2_X1   g656(.A(new_n465), .B(KEYINPUT57), .Z(new_n843));
  AND2_X1   g657(.A1(new_n827), .A2(KEYINPUT54), .ZN(new_n844));
  INV_X1    g658(.A(new_n791), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n463), .B2(new_n460), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n827), .A2(G902), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n720), .B(KEYINPUT121), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n840), .B1(new_n847), .B2(new_n850), .ZN(G54));
  NAND3_X1  g665(.A1(new_n848), .A2(KEYINPUT58), .A3(G475), .ZN(new_n852));
  INV_X1    g666(.A(new_n391), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n854), .A2(new_n855), .A3(new_n840), .ZN(G60));
  NAND2_X1  g670(.A1(new_n592), .A2(new_n593), .ZN(new_n857));
  NAND2_X1  g671(.A1(G478), .A2(G902), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT59), .Z(new_n859));
  NOR2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n844), .B2(new_n845), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n841), .ZN(new_n862));
  INV_X1    g676(.A(new_n859), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n792), .B2(new_n793), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n862), .B1(new_n864), .B2(new_n857), .ZN(G63));
  NAND2_X1  g679(.A1(G217), .A2(G902), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT122), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT60), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n827), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n614), .B(KEYINPUT123), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n871), .B(new_n841), .C1(new_n500), .C2(new_n869), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n869), .A2(new_n500), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT61), .A3(new_n841), .A4(new_n871), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(G66));
  AOI21_X1  g691(.A(new_n242), .B1(new_n334), .B2(G224), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n759), .A2(new_n760), .ZN(new_n879));
  INV_X1    g693(.A(new_n749), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n878), .B1(new_n882), .B2(new_n242), .ZN(new_n883));
  INV_X1    g697(.A(G898), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n830), .B1(new_n884), .B2(G953), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n883), .B(new_n885), .ZN(G69));
  NAND2_X1  g700(.A1(new_n581), .A2(new_n747), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n632), .A3(new_n700), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n728), .A2(new_n734), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n644), .A2(new_n627), .A3(new_n771), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n888), .B(new_n889), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(G953), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n525), .A2(new_n529), .A3(new_n531), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n356), .A2(new_n359), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n897), .B(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n771), .A2(new_n627), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n726), .A2(new_n762), .A3(new_n797), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n889), .A2(new_n750), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n242), .ZN(new_n904));
  NAND2_X1  g718(.A1(G900), .A2(G953), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n899), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n242), .B1(G227), .B2(G900), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT125), .Z(new_n909));
  OR3_X1    g723(.A1(new_n907), .A2(KEYINPUT126), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT126), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n907), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G72));
  NAND2_X1  g727(.A1(G472), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT63), .Z(new_n915));
  NAND3_X1  g729(.A1(new_n532), .A2(new_n534), .A3(new_n542), .ZN(new_n916));
  AND4_X1   g730(.A1(new_n638), .A2(new_n782), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n894), .A2(new_n881), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n915), .B(KEYINPUT127), .Z(new_n919));
  AOI21_X1  g733(.A(new_n638), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n881), .A2(new_n903), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n921), .B2(new_n919), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n917), .A2(new_n920), .A3(new_n840), .A4(new_n922), .ZN(G57));
endmodule


