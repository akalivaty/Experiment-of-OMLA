//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  INV_X1    g034(.A(new_n456), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT68), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n471), .A3(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n472), .B2(KEYINPUT70), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n469), .A2(new_n471), .A3(new_n474), .A4(G125), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n465), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n468), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n465), .A2(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT71), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(new_n470), .A3(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n482), .A3(new_n469), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n478), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n476), .A2(new_n484), .ZN(G160));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n465), .C2(G112), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n483), .A2(new_n465), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G124), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n480), .A2(new_n482), .A3(new_n469), .ZN(new_n491));
  INV_X1    g066(.A(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(G136), .B2(new_n494), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n492), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(G138), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n469), .A2(new_n471), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G114), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT4), .A2(G138), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n465), .A2(new_n507), .B1(G126), .B2(G2105), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n502), .B(new_n506), .C1(new_n508), .C2(new_n483), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n512), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT72), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT72), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n513), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n523), .A2(G88), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n524), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G50), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n527), .A2(KEYINPUT73), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(KEYINPUT73), .B1(new_n527), .B2(new_n529), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n516), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G166));
  AND2_X1   g108(.A1(new_n523), .A2(new_n526), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n539), .B1(G51), .B2(new_n528), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n535), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n519), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n528), .B2(G52), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n523), .A2(G90), .A3(new_n526), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n519), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(new_n528), .B2(G43), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n523), .A2(G81), .A3(new_n526), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n524), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n570), .A2(new_n571), .B1(KEYINPUT77), .B2(KEYINPUT9), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT77), .B(KEYINPUT9), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n524), .A2(new_n573), .A3(G53), .A4(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n519), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G651), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n523), .A2(G91), .A3(new_n526), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n575), .A2(new_n579), .A3(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n532), .A2(KEYINPUT78), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n583), .B(new_n516), .C1(new_n530), .C2(new_n531), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n582), .A2(new_n584), .ZN(G303));
  NAND3_X1  g160(.A1(new_n524), .A2(G49), .A3(G543), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n524), .A2(KEYINPUT79), .A3(G49), .A4(G543), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n523), .A2(G87), .A3(new_n526), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(G73), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G61), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n595), .B1(new_n511), .B2(new_n512), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n594), .B1(new_n596), .B2(KEYINPUT80), .ZN(new_n597));
  OAI211_X1 g172(.A(KEYINPUT80), .B(G61), .C1(new_n517), .C2(new_n518), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n523), .A2(G86), .A3(new_n526), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n528), .A2(G48), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(G305));
  XNOR2_X1  g178(.A(KEYINPUT81), .B(G85), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n534), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n519), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(new_n528), .B2(G47), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  NAND3_X1  g185(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n523), .A2(new_n526), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(G79), .A2(G543), .ZN(new_n617));
  INV_X1    g192(.A(G66), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n519), .B2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(new_n528), .B2(G54), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  MUX2_X1   g196(.A(new_n621), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g197(.A(new_n621), .B(G301), .S(G868), .Z(G321));
  INV_X1    g198(.A(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(G299), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G168), .B2(new_n624), .ZN(G280));
  XNOR2_X1  g201(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g202(.A(new_n621), .ZN(new_n628));
  INV_X1    g203(.A(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(G860), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT83), .ZN(G148));
  OAI21_X1  g206(.A(new_n624), .B1(new_n561), .B2(new_n562), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n621), .A2(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(new_n624), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n487), .A2(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n465), .C2(G111), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n493), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n492), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT12), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  INV_X1    g218(.A(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n654), .A2(new_n657), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT85), .Z(new_n662));
  AOI21_X1  g237(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n663));
  INV_X1    g238(.A(G14), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT17), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT87), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n671), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n674), .B(new_n670), .C1(new_n667), .C2(new_n671), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n669), .A2(new_n667), .A3(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n644), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT88), .B(G2096), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n687), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n687), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1986), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT89), .B(KEYINPUT90), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n701), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(G229));
  AND3_X1   g281(.A1(new_n491), .A2(G131), .A3(new_n492), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT91), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(new_n465), .ZN(new_n710));
  INV_X1    g285(.A(G107), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n487), .B2(G119), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n708), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G25), .B2(G29), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  AND2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G24), .ZN(new_n722));
  INV_X1    g297(.A(G290), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n721), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1986), .ZN(new_n725));
  OR3_X1    g300(.A1(new_n719), .A2(new_n720), .A3(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G23), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n721), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT33), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G1976), .ZN(new_n731));
  MUX2_X1   g306(.A(G6), .B(G305), .S(G16), .Z(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT32), .B(G1981), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G22), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G166), .B2(G16), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n734), .B1(new_n736), .B2(G1971), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(G1971), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n731), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n726), .B1(KEYINPUT34), .B2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(KEYINPUT34), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(KEYINPUT36), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n740), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(G168), .A2(G16), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT97), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G16), .B2(G21), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(KEYINPUT97), .B2(new_n747), .ZN(new_n751));
  INV_X1    g326(.A(G1966), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n754), .A2(G33), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n494), .A2(G139), .ZN(new_n756));
  INV_X1    g331(.A(G127), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n501), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G115), .B2(G2104), .ZN(new_n759));
  NAND2_X1  g334(.A1(G103), .A2(G2104), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n710), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(KEYINPUT25), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n710), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  OAI221_X1 g339(.A(new_n756), .B1(new_n465), .B2(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n755), .B1(new_n765), .B2(G29), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(new_n442), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n721), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n721), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n768), .B1(G1961), .B2(new_n770), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n753), .B(new_n771), .C1(G1961), .C2(new_n770), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n754), .A2(G27), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G164), .B2(new_n754), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT98), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(new_n443), .ZN(new_n776));
  NAND2_X1  g351(.A1(G160), .A2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n778), .B2(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT24), .B2(new_n778), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G2084), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n754), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI221_X1 g360(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n465), .C2(G116), .ZN(new_n786));
  INV_X1    g361(.A(G140), .ZN(new_n787));
  INV_X1    g362(.A(G128), .ZN(new_n788));
  OAI221_X1 g363(.A(new_n786), .B1(new_n493), .B2(new_n787), .C1(new_n488), .C2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n785), .B1(new_n790), .B2(new_n754), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT94), .B(G2067), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n776), .A2(new_n782), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n766), .A2(new_n442), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n639), .A2(new_n754), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT30), .B(G28), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT31), .A2(G11), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n797), .A2(new_n754), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n795), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n754), .A2(G32), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n494), .A2(G141), .B1(G105), .B2(new_n477), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n487), .A2(G129), .ZN(new_n804));
  NAND3_X1  g379(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT26), .ZN(new_n807));
  AND3_X1   g382(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n802), .B1(new_n808), .B2(new_n754), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT27), .B(G1996), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n801), .B(new_n811), .C1(G2084), .C2(new_n781), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n754), .A2(G35), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G162), .B2(new_n754), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT29), .B(G2090), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n563), .A2(new_n721), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n721), .B2(G19), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT92), .B(G1341), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n794), .A2(new_n812), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(G4), .A2(G16), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(new_n628), .B2(G16), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1348), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n818), .A2(new_n819), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n721), .A2(G20), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT23), .ZN(new_n827));
  INV_X1    g402(.A(G299), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n721), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1956), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n824), .A2(new_n825), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n772), .A2(new_n821), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n746), .A2(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n519), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(KEYINPUT99), .B(G55), .Z(new_n838));
  AOI22_X1  g413(.A1(new_n837), .A2(G651), .B1(new_n528), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT100), .B(G93), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n523), .A2(new_n526), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n561), .B2(new_n562), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n557), .A2(new_n559), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n842), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT38), .Z(new_n848));
  NOR2_X1   g423(.A1(new_n621), .A2(new_n629), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g426(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n842), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(G145));
  NAND2_X1  g431(.A1(new_n487), .A2(G130), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT101), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n494), .A2(G142), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n465), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n858), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n789), .B(new_n509), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n714), .B(KEYINPUT102), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(new_n642), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n714), .B(KEYINPUT102), .ZN(new_n868));
  INV_X1    g443(.A(new_n642), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n808), .B(new_n765), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n867), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n867), .B2(new_n870), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n865), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n867), .A2(new_n870), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n871), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n867), .A2(new_n870), .A3(new_n872), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n877), .A2(new_n864), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n639), .B(G160), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(G162), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  INV_X1    g459(.A(new_n882), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n875), .A2(new_n879), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g463(.A1(new_n842), .A2(new_n624), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(G305), .B(G288), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n532), .A2(new_n723), .ZN(new_n892));
  OAI211_X1 g467(.A(G290), .B(new_n516), .C1(new_n531), .C2(new_n530), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(new_n893), .B2(new_n892), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(KEYINPUT104), .A3(new_n894), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n895), .B2(new_n896), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n897), .B1(new_n902), .B2(new_n890), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n621), .A2(new_n828), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n616), .A2(G299), .A3(new_n620), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(KEYINPUT41), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  INV_X1    g484(.A(new_n905), .ZN(new_n910));
  AOI21_X1  g485(.A(G299), .B1(new_n616), .B2(new_n620), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n904), .A2(KEYINPUT103), .A3(KEYINPUT41), .A4(new_n905), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n847), .B(new_n633), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n904), .A2(new_n905), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n903), .B(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n889), .B1(new_n919), .B2(new_n624), .ZN(G295));
  OAI21_X1  g495(.A(new_n889), .B1(new_n919), .B2(new_n624), .ZN(G331));
  NAND2_X1  g496(.A1(new_n546), .A2(new_n548), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT74), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n923), .A2(G286), .A3(new_n549), .ZN(new_n924));
  AOI21_X1  g499(.A(G286), .B1(new_n923), .B2(new_n549), .ZN(new_n925));
  INV_X1    g500(.A(new_n842), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n844), .A2(KEYINPUT75), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(new_n560), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n924), .A2(new_n925), .B1(new_n928), .B2(new_n845), .ZN(new_n929));
  OAI21_X1  g504(.A(G168), .B1(new_n550), .B2(new_n551), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(G286), .A3(new_n549), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n930), .A2(new_n843), .A3(new_n846), .A4(new_n931), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n929), .A2(new_n932), .A3(new_n917), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n932), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n902), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n902), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n899), .A2(new_n901), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n910), .A2(new_n911), .A3(new_n909), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n912), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n906), .A2(KEYINPUT105), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n943), .B(new_n935), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n929), .A2(new_n932), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT41), .B1(new_n904), .B2(new_n905), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(KEYINPUT105), .B2(new_n906), .ZN(new_n951));
  INV_X1    g526(.A(new_n947), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n917), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT106), .B1(new_n935), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n942), .B(new_n948), .C1(new_n953), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n938), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n940), .A2(new_n941), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n938), .A2(new_n956), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n938), .A2(new_n956), .A3(KEYINPUT107), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(KEYINPUT43), .A3(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n937), .A2(new_n938), .A3(new_n957), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n966), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g542(.A(new_n808), .B(G1996), .ZN(new_n968));
  INV_X1    g543(.A(G2067), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n789), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n714), .B(new_n718), .Z(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(G290), .B(G1986), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G40), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n476), .A2(new_n976), .A3(new_n484), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT45), .B1(new_n509), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT108), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n975), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G8), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n509), .A2(new_n978), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(new_n977), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n590), .A2(new_n591), .A3(G1976), .A4(new_n592), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(KEYINPUT110), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT52), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n985), .A2(new_n987), .A3(new_n988), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n601), .A2(new_n602), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n995), .A2(KEYINPUT111), .A3(new_n697), .A4(new_n600), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n600), .A2(new_n697), .A3(new_n601), .A4(new_n602), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G305), .A2(G1981), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1000), .A2(KEYINPUT49), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT49), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n994), .B1(new_n1004), .B2(new_n985), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n582), .A2(G8), .A3(new_n584), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n582), .A2(KEYINPUT55), .A3(G8), .A4(new_n584), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n472), .A2(KEYINPUT70), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(new_n475), .A3(new_n466), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n710), .ZN(new_n1014));
  INV_X1    g589(.A(new_n484), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(G40), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1011), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n509), .A2(new_n978), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1971), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n509), .A2(new_n1023), .A3(new_n978), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n509), .B2(new_n978), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n1016), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT109), .B(G2090), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n983), .B1(new_n1022), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1005), .A2(new_n1010), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n728), .A2(new_n991), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT112), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1000), .B1(new_n1004), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n985), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT63), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1010), .A2(new_n1030), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n977), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n1026), .B2(new_n1016), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1025), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1021), .B1(new_n1043), .B2(new_n1028), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1008), .B(new_n1009), .C1(new_n1044), .C2(new_n983), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1005), .A2(new_n1038), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n509), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n977), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n752), .B1(new_n1048), .B2(new_n979), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1020), .A2(new_n1047), .A3(new_n977), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(KEYINPUT114), .A3(new_n752), .ZN(new_n1053));
  INV_X1    g628(.A(G2084), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1027), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(G8), .A3(G168), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1037), .B1(new_n1046), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n1010), .A2(new_n1030), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1057), .A2(new_n1037), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1038), .A4(new_n1005), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1036), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1020), .A2(new_n443), .A3(new_n1047), .A4(new_n977), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1064));
  NAND3_X1  g639(.A1(new_n1039), .A2(new_n977), .A3(new_n1024), .ZN(new_n1065));
  INV_X1    g640(.A(G1961), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1063), .A2(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1063), .A2(KEYINPUT122), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT53), .B1(new_n1063), .B2(KEYINPUT122), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(G171), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT124), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1073), .A3(G171), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1011), .A2(new_n979), .A3(new_n1016), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(KEYINPUT53), .A4(new_n443), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT125), .B1(new_n1063), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(G301), .A3(new_n1067), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT126), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT126), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1080), .A2(new_n1083), .A3(G301), .A4(new_n1067), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1072), .A2(new_n1074), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1070), .A2(G171), .ZN(new_n1088));
  AOI21_X1  g663(.A(G301), .B1(new_n1080), .B2(new_n1067), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1086), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n1046), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1051), .A2(G168), .A3(new_n1055), .A4(new_n1053), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1049), .A2(new_n1050), .B1(new_n1027), .B2(new_n1054), .ZN(new_n1094));
  AOI21_X1  g669(.A(G168), .B1(new_n1094), .B2(new_n1053), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1093), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT51), .B1(new_n1092), .B2(G8), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT121), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1056), .A2(G286), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1100), .A2(KEYINPUT51), .A3(G8), .A4(new_n1092), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1087), .A2(new_n1091), .A3(new_n1099), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(G1348), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1065), .A2(new_n1106), .B1(new_n969), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(new_n621), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT119), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n575), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n572), .A2(KEYINPUT116), .A3(new_n574), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n580), .A2(new_n579), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT117), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1114), .A2(new_n1116), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT115), .B(G1956), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1043), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT56), .B(G2072), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1075), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1118), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1024), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1123), .B1(new_n1126), .B2(new_n1119), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(KEYINPUT118), .A3(new_n1117), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1075), .A2(new_n1122), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1117), .B(new_n1129), .C1(new_n1043), .C2(new_n1120), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1110), .A2(new_n1124), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1127), .B2(new_n1117), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT120), .B(new_n1118), .C1(new_n1121), .C2(new_n1123), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1130), .B(KEYINPUT118), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1124), .A2(KEYINPUT61), .A3(new_n1130), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1108), .A2(new_n621), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT60), .B1(new_n1142), .B2(new_n1109), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT58), .B(G1341), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1052), .A2(G1996), .B1(new_n1107), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n563), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT59), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1148), .A3(new_n563), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n621), .A2(KEYINPUT60), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1147), .A2(new_n1149), .B1(new_n1108), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1141), .A2(new_n1143), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1133), .B1(new_n1140), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1062), .B1(new_n1105), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1102), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1099), .A2(KEYINPUT62), .A3(new_n1104), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1046), .B1(new_n1074), .B2(new_n1072), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n982), .B1(new_n1154), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n715), .A2(new_n718), .ZN(new_n1163));
  OAI22_X1  g738(.A1(new_n971), .A2(new_n1163), .B1(G2067), .B2(new_n789), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n981), .ZN(new_n1165));
  INV_X1    g740(.A(new_n981), .ZN(new_n1166));
  OR3_X1    g741(.A1(new_n1166), .A2(G1986), .A3(G290), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT48), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n1166), .B2(new_n973), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT47), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1166), .A2(G1996), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT46), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n970), .A2(new_n808), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1174), .B1(new_n981), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1174), .B2(new_n1173), .ZN(new_n1177));
  OAI221_X1 g752(.A(new_n1165), .B1(new_n1170), .B2(new_n1171), .C1(new_n1172), .C2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1178), .B1(new_n1172), .B2(new_n1177), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1162), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g755(.A1(new_n940), .A2(new_n958), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n682), .A2(new_n461), .A3(new_n683), .ZN(new_n1183));
  NOR2_X1   g757(.A1(G401), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g758(.A1(new_n887), .A2(new_n1182), .A3(new_n705), .A4(new_n1184), .ZN(G225));
  INV_X1    g759(.A(G225), .ZN(G308));
endmodule


