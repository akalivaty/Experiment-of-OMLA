//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  INV_X1    g047(.A(new_n461), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n473), .B1(new_n470), .B2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n467), .B(new_n472), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OR2_X1    g054(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT65), .A2(G2104), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(KEYINPUT3), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n461), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n483), .A2(new_n475), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  INV_X1    g062(.A(G100), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n488), .A2(new_n475), .A3(KEYINPUT66), .ZN(new_n489));
  AOI21_X1  g064(.A(KEYINPUT66), .B1(new_n488), .B2(new_n475), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G112), .B2(new_n475), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n485), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  AND2_X1   g068(.A1(new_n461), .A2(new_n463), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n495), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n482), .A2(new_n461), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(KEYINPUT4), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n474), .A2(G126), .A3(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT67), .B(G114), .ZN(new_n503));
  OAI211_X1 g078(.A(G2104), .B(new_n502), .C1(new_n503), .C2(new_n475), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n500), .A2(new_n505), .ZN(G164));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT70), .A3(G62), .ZN(new_n508));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT71), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT70), .B1(new_n507), .B2(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(G651), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT72), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n515), .B(G651), .C1(new_n511), .C2(new_n512), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT6), .B1(new_n517), .B2(new_n519), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g097(.A(new_n517), .B(KEYINPUT6), .C1(new_n518), .C2(new_n519), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n522), .A2(G88), .A3(new_n507), .A4(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n522), .A2(G50), .A3(G543), .A4(new_n523), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n514), .A2(new_n516), .A3(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(new_n522), .A2(G543), .A3(new_n523), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT73), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n522), .A2(new_n531), .A3(G543), .A4(new_n523), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n522), .A2(new_n523), .ZN(new_n538));
  INV_X1    g113(.A(new_n507), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  XOR2_X1   g116(.A(KEYINPUT74), .B(G89), .Z(new_n542));
  OAI211_X1 g117(.A(new_n536), .B(new_n537), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n534), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n519), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(G52), .B2(new_n533), .ZN(G171));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n533), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n540), .A2(G81), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n519), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n550), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NOR3_X1   g131(.A1(new_n551), .A2(new_n554), .A3(new_n550), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  AOI22_X1  g138(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n564), .A2(new_n519), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n540), .B2(G91), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(new_n529), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n567), .B1(new_n568), .B2(G53), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  NOR3_X1   g145(.A1(new_n529), .A2(KEYINPUT9), .A3(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n566), .B1(new_n569), .B2(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n533), .A2(G52), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n573), .B(new_n546), .C1(new_n547), .C2(new_n541), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  NAND2_X1  g150(.A1(new_n540), .A2(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n568), .A2(G49), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n539), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n568), .A2(G48), .B1(G651), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n522), .A2(G86), .A3(new_n507), .A4(new_n523), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(KEYINPUT76), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(KEYINPUT76), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n583), .B1(new_n586), .B2(new_n587), .ZN(G305));
  AND2_X1   g163(.A1(new_n533), .A2(G47), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n540), .A2(G85), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n519), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G301), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n530), .A2(KEYINPUT77), .A3(new_n532), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT77), .B1(new_n530), .B2(new_n532), .ZN(new_n599));
  OAI21_X1  g174(.A(G54), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n519), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n522), .A2(G92), .A3(new_n507), .A4(new_n523), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g182(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n600), .A2(KEYINPUT78), .A3(new_n607), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n596), .B1(new_n611), .B2(new_n595), .ZN(G284));
  XOR2_X1   g187(.A(G284), .B(KEYINPUT79), .Z(G321));
  NOR2_X1   g188(.A1(G286), .A2(new_n595), .ZN(new_n614));
  XOR2_X1   g189(.A(G299), .B(KEYINPUT80), .Z(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n595), .ZN(G297));
  AOI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n595), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NOR2_X1   g194(.A1(new_n558), .A2(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n611), .A2(new_n618), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G868), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n471), .A2(new_n494), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT13), .B(G2100), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n484), .A2(G135), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n486), .A2(G123), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(G14), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(KEYINPUT14), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT84), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n643), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n649), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n653), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n638), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n654), .A2(new_n658), .ZN(new_n662));
  INV_X1    g237(.A(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT86), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n665), .A3(new_n660), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT88), .Z(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n672), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT17), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n672), .A2(new_n669), .A3(new_n676), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n676), .B(KEYINPUT89), .Z(new_n682));
  OAI211_X1 g257(.A(new_n678), .B(new_n681), .C1(new_n674), .C2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n692), .B(new_n695), .C1(new_n687), .C2(new_n691), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(G229));
  NOR2_X1   g277(.A1(G29), .A2(G33), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT97), .B(KEYINPUT25), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n494), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(new_n475), .ZN(new_n708));
  AOI211_X1 g283(.A(new_n706), .B(new_n708), .C1(G139), .C2(new_n484), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(G29), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G2072), .Z(new_n711));
  INV_X1    g286(.A(G2084), .ZN(new_n712));
  INV_X1    g287(.A(G34), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n713), .A2(KEYINPUT24), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(KEYINPUT24), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(KEYINPUT98), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(KEYINPUT98), .B2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n478), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n711), .B1(new_n712), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G1961), .ZN(new_n721));
  NOR2_X1   g296(.A1(G5), .A2(G16), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT103), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(G301), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n720), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(G19), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n558), .B2(new_n724), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n726), .B1(G1341), .B2(new_n728), .C1(new_n721), .C2(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n718), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n484), .A2(G140), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n486), .A2(G128), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n475), .A2(G116), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT96), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n731), .B1(new_n738), .B2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G2067), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n728), .A2(G1341), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n729), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G4), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n611), .B2(G16), .ZN(new_n745));
  INV_X1    g320(.A(G1348), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT26), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n484), .A2(G141), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n749), .B(new_n750), .C1(G105), .C2(new_n471), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n486), .A2(G129), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT99), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(new_n718), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT100), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G29), .B2(G32), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(KEYINPUT100), .B2(new_n755), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT101), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n718), .A2(G35), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G162), .B2(new_n718), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT29), .ZN(new_n765));
  INV_X1    g340(.A(G2090), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT31), .B(G11), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n769), .A2(G28), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n718), .B1(new_n769), .B2(G28), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n768), .B1(new_n770), .B2(new_n771), .C1(new_n634), .C2(new_n718), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n712), .B2(new_n719), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n718), .A2(G27), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G164), .B2(new_n718), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT104), .B(G2078), .Z(new_n776));
  OAI21_X1  g351(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n767), .B(new_n778), .C1(new_n759), .C2(new_n760), .ZN(new_n779));
  NOR2_X1   g354(.A1(G286), .A2(new_n724), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT102), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(KEYINPUT102), .B1(G16), .B2(G21), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(G1966), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n724), .A2(G20), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT23), .Z(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G299), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n784), .A2(G1966), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n779), .A2(new_n785), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n743), .A2(new_n747), .A3(new_n762), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n718), .A2(G25), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n486), .A2(G119), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT92), .Z(new_n796));
  OR2_X1    g371(.A1(G95), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n484), .A2(G131), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n794), .B1(new_n803), .B2(new_n718), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  XOR2_X1   g380(.A(new_n804), .B(new_n805), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n724), .A2(G24), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n593), .B2(new_n724), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT93), .B(G1986), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n724), .A2(G23), .ZN(new_n812));
  INV_X1    g387(.A(G288), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n724), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT33), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1976), .ZN(new_n816));
  NOR2_X1   g391(.A1(G16), .A2(G22), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G166), .B2(G16), .ZN(new_n818));
  INV_X1    g393(.A(G1971), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  MUX2_X1   g395(.A(G6), .B(G305), .S(G16), .Z(new_n821));
  XOR2_X1   g396(.A(KEYINPUT32), .B(G1981), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n816), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT95), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT95), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n811), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n828), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n825), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n834), .A3(new_n831), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n793), .B1(new_n833), .B2(new_n835), .ZN(G311));
  INV_X1    g411(.A(new_n793), .ZN(new_n837));
  INV_X1    g412(.A(new_n835), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n834), .B1(new_n829), .B2(new_n831), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(G150));
  AND2_X1   g415(.A1(new_n533), .A2(G55), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n540), .A2(G93), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n519), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n557), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n555), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n551), .A2(new_n554), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT38), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n611), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n855));
  AOI21_X1  g430(.A(G860), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g432(.A(G860), .B1(new_n841), .B2(new_n844), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT37), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(G145));
  XNOR2_X1  g435(.A(new_n634), .B(new_n478), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n492), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n802), .B(new_n627), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n754), .B(new_n709), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n501), .A2(new_n504), .ZN(new_n866));
  AOI221_X4 g441(.A(KEYINPUT105), .B1(new_n494), .B2(new_n496), .C1(new_n499), .C2(KEYINPUT4), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n494), .A2(new_n496), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n866), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n738), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n486), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n475), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n877), .B1(G142), .B2(new_n484), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT106), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n873), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n865), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n865), .A2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n862), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(new_n862), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n881), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g465(.A(new_n621), .B(new_n851), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n600), .A2(new_n607), .ZN(new_n892));
  INV_X1    g467(.A(G299), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT107), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n895));
  AOI211_X1 g470(.A(new_n895), .B(G299), .C1(new_n600), .C2(new_n607), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n608), .A2(G299), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G288), .B(KEYINPUT111), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(G305), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n593), .B(G303), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n902), .B(new_n903), .Z(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT42), .Z(new_n905));
  XOR2_X1   g480(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n899), .A2(KEYINPUT110), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n895), .B1(new_n608), .B2(G299), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT107), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT108), .B1(new_n894), .B2(new_n896), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n898), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n897), .A2(new_n898), .A3(new_n907), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT110), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n908), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n891), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n900), .A2(new_n905), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n905), .B1(new_n900), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G868), .B2(new_n845), .ZN(G295));
  OAI21_X1  g500(.A(new_n924), .B1(G868), .B2(new_n845), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n928));
  NOR3_X1   g503(.A1(G171), .A2(G168), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(new_n928), .ZN(new_n931));
  NAND2_X1  g506(.A1(G301), .A2(KEYINPUT112), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(G168), .A3(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n848), .A2(new_n930), .A3(new_n850), .A4(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  INV_X1    g510(.A(new_n850), .ZN(new_n936));
  OAI22_X1  g511(.A1(new_n935), .A2(new_n929), .B1(new_n847), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n908), .A2(new_n916), .A3(new_n919), .A4(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n899), .A2(new_n934), .A3(new_n937), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n904), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n888), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n904), .B1(new_n939), .B2(new_n940), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n927), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n943), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n906), .B1(new_n934), .B2(new_n937), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n946), .A2(new_n914), .B1(new_n947), .B2(new_n899), .ZN(new_n948));
  AOI21_X1  g523(.A(G37), .B1(new_n948), .B2(new_n904), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n949), .A3(KEYINPUT43), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n944), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT44), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n942), .B2(new_n943), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n945), .A2(new_n949), .A3(new_n927), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n952), .A2(new_n957), .ZN(G397));
  XOR2_X1   g533(.A(new_n802), .B(new_n805), .Z(new_n959));
  XOR2_X1   g534(.A(new_n754), .B(G1996), .Z(new_n960));
  XNOR2_X1  g535(.A(new_n738), .B(new_n740), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n593), .B(G1986), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT4), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n474), .B2(new_n498), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT105), .B1(new_n968), .B2(new_n497), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n869), .A2(new_n868), .A3(new_n870), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n505), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n971), .B2(G1384), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n872), .A2(KEYINPUT113), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n484), .A2(G137), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(new_n467), .A3(G40), .A4(new_n472), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n965), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n981));
  AND3_X1   g556(.A1(G303), .A2(G8), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(G303), .B2(G8), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT116), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  INV_X1    g560(.A(new_n981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n988));
  NAND3_X1  g563(.A1(G303), .A2(G8), .A3(new_n981), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n974), .B1(new_n500), .B2(new_n505), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n978), .B1(new_n993), .B2(new_n973), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT114), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n995), .B1(new_n992), .B2(new_n994), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n996), .A2(new_n997), .A3(G1971), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n872), .A2(new_n999), .A3(new_n974), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n978), .B1(new_n993), .B2(KEYINPUT50), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(G2090), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n991), .B(G8), .C1(new_n998), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT63), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1000), .A2(new_n1001), .A3(new_n712), .ZN(new_n1007));
  INV_X1    g582(.A(new_n978), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT45), .B(new_n974), .C1(new_n500), .C2(new_n505), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n872), .A2(new_n974), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n973), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1007), .B1(new_n1012), .B2(G1966), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(G8), .A3(G168), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1005), .A2(new_n1006), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(G8), .B1(new_n998), .B2(new_n1003), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n982), .A2(new_n983), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n969), .A2(new_n970), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n1019), .B2(new_n866), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n1008), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n813), .A2(G1976), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(G8), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT52), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1021), .A2(new_n1022), .A3(G8), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n583), .A2(new_n584), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(new_n583), .C1(new_n587), .C2(new_n586), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT49), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(new_n1031), .A3(KEYINPUT49), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1034), .A2(G8), .A3(new_n1021), .A4(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1024), .A2(new_n1027), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT121), .B1(new_n1018), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n992), .A2(new_n994), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(KEYINPUT114), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n819), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1003), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1017), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1037), .B(KEYINPUT121), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1015), .B1(new_n1038), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n999), .B1(new_n872), .B2(new_n974), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n978), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT118), .B(new_n1008), .C1(new_n1020), .C2(new_n999), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n993), .A2(KEYINPUT50), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n766), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1043), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1039), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(new_n1043), .A3(KEYINPUT119), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1046), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1004), .A2(new_n1037), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1014), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1049), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1021), .A2(G8), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT117), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1036), .A2(new_n1025), .A3(new_n813), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1031), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(new_n1005), .B2(new_n1037), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n992), .A2(new_n994), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1074), .B2(new_n789), .ZN(new_n1075));
  XNOR2_X1  g650(.A(G299), .B(KEYINPUT57), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1070), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1079), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1054), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n978), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(KEYINPUT118), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1956), .B1(new_n1083), .B2(new_n1052), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT123), .B(new_n1076), .C1(new_n1084), .C2(new_n1073), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(new_n1080), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1021), .A2(G2067), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1000), .A2(new_n1001), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1091), .B2(new_n746), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n611), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n609), .A2(new_n610), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1002), .A2(KEYINPUT122), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1000), .A2(new_n1001), .A3(new_n1088), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n746), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1087), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT60), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1094), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1093), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1074), .A2(new_n789), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1077), .B1(new_n1104), .B2(new_n1072), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1076), .B(new_n1073), .C1(new_n1074), .C2(new_n789), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1079), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1021), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(G1996), .B2(new_n1040), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n558), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT59), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1086), .A2(new_n1103), .A3(new_n1107), .A4(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1078), .B(new_n1085), .C1(new_n1094), .C2(new_n1092), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1106), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n976), .A2(new_n1008), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(G2078), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n976), .A2(KEYINPUT124), .A3(new_n1008), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1120), .A2(new_n992), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G2078), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1125), .B1(new_n996), .B2(new_n997), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1126), .A2(new_n1121), .B1(new_n1091), .B2(new_n721), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G171), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1012), .A2(new_n1122), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1095), .A2(new_n721), .A3(new_n1096), .ZN(new_n1132));
  AOI21_X1  g707(.A(G2078), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1131), .B(new_n1132), .C1(new_n1133), .C2(KEYINPUT53), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1127), .A2(KEYINPUT125), .A3(G301), .A4(new_n1131), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1129), .A2(KEYINPUT54), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1124), .A2(new_n1127), .A3(G301), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1134), .A2(G171), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(G8), .A3(new_n1059), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1061), .B1(new_n1144), .B2(new_n1017), .ZN(new_n1145));
  OAI211_X1 g720(.A(new_n1007), .B(G168), .C1(new_n1012), .C2(G1966), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT51), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1146), .A2(new_n1147), .A3(G8), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1013), .A2(G286), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(G8), .A3(new_n1146), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1148), .B1(new_n1150), .B2(KEYINPUT51), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1137), .A2(new_n1142), .A3(new_n1145), .A4(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1064), .B(new_n1069), .C1(new_n1117), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1139), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1156), .A2(new_n1145), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1156), .B2(new_n1145), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n980), .B1(new_n1154), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n979), .ZN(new_n1163));
  INV_X1    g738(.A(new_n754), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1163), .B1(new_n961), .B2(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT127), .Z(new_n1166));
  NOR2_X1   g741(.A1(new_n1163), .A2(G1996), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT46), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1169), .B(KEYINPUT47), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n803), .A2(new_n805), .ZN(new_n1171));
  OAI22_X1  g746(.A1(new_n962), .A2(new_n1171), .B1(G2067), .B2(new_n738), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(new_n979), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT48), .ZN(new_n1174));
  OR3_X1    g749(.A1(new_n1163), .A2(G1986), .A3(G290), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n963), .A2(new_n1163), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1175), .A2(new_n1174), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1173), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1170), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1162), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g755(.A1(G229), .A2(new_n457), .A3(G227), .ZN(new_n1182));
  AND4_X1   g756(.A1(new_n667), .A2(new_n955), .A3(new_n889), .A4(new_n1182), .ZN(G308));
  NAND4_X1  g757(.A1(new_n667), .A2(new_n955), .A3(new_n889), .A4(new_n1182), .ZN(G225));
endmodule


