//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AND2_X1   g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n459), .A2(KEYINPUT67), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(KEYINPUT67), .B1(G567), .B2(new_n456), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT3), .B(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(new_n463), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n476), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n483), .A2(G137), .B1(G101), .B2(new_n464), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n474), .A2(new_n487), .ZN(G160));
  NOR2_X1   g063(.A1(new_n477), .A2(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n483), .A2(G136), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n463), .B2(G114), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G102), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n463), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n497), .A2(new_n499), .A3(G2104), .A4(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G126), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n475), .B2(new_n476), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n506), .B(new_n509), .C1(new_n476), .C2(new_n475), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n504), .B1(new_n508), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT70), .A3(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(new_n516), .B1(KEYINPUT5), .B2(new_n513), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n522), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n520), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AND3_X1   g105(.A1(new_n517), .A2(G89), .A3(new_n525), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(new_n523), .ZN(new_n535));
  INV_X1    g110(.A(G51), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR3_X1   g112(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n517), .A2(G64), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n519), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n517), .A2(G90), .A3(new_n525), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n523), .A2(G52), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(G171));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n514), .A2(new_n516), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n547), .A2(G81), .A3(new_n525), .A4(new_n548), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n523), .A2(G43), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n552), .B(KEYINPUT72), .C1(new_n556), .C2(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AOI22_X1  g143(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n569), .A2(new_n519), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n523), .A2(new_n572), .A3(G53), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n572), .B1(new_n523), .B2(G53), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT73), .ZN(new_n576));
  INV_X1    g151(.A(new_n526), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n577), .A2(G91), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n571), .A2(new_n575), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(G91), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n573), .A2(new_n574), .B1(new_n526), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT73), .B1(new_n581), .B2(new_n570), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND2_X1  g161(.A1(new_n577), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n523), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n519), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n523), .A2(G48), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n526), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n523), .A2(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n526), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT74), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n519), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n547), .A2(G66), .A3(new_n548), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n519), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n523), .A2(G54), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n607), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OAI211_X1 g189(.A(KEYINPUT75), .B(new_n611), .C1(new_n614), .C2(new_n519), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n577), .A2(KEYINPUT10), .A3(G92), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n526), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n606), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n606), .B1(new_n623), .B2(G868), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(new_n583), .B2(G868), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(new_n583), .B2(G868), .ZN(G280));
  XNOR2_X1  g203(.A(KEYINPUT76), .B(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n623), .B1(G860), .B2(new_n629), .ZN(G148));
  NAND2_X1  g205(.A1(new_n623), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n466), .A2(new_n464), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  INV_X1    g213(.A(G2100), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n489), .A2(G123), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n483), .A2(G135), .ZN(new_n643));
  OR2_X1    g218(.A1(G99), .A2(G2105), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n644), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(G2096), .Z(new_n647));
  NAND3_X1  g222(.A1(new_n640), .A2(new_n641), .A3(new_n647), .ZN(G156));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(KEYINPUT14), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G1341), .B(G1348), .Z(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G14), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n662), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(G401));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT80), .B(KEYINPUT18), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT81), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(KEYINPUT17), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n676), .A2(new_n671), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n673), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2096), .B(G2100), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n689), .A2(new_n692), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n686), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n698), .B(new_n699), .ZN(new_n703));
  NOR3_X1   g278(.A1(new_n703), .A2(new_n696), .A3(KEYINPUT83), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n685), .B1(new_n702), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(G1991), .B(G1996), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n697), .A2(new_n701), .A3(new_n686), .ZN(new_n708));
  OAI21_X1  g283(.A(KEYINPUT83), .B1(new_n703), .B2(new_n696), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n708), .A2(new_n709), .A3(new_n684), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n705), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n707), .B1(new_n705), .B2(new_n710), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n683), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n705), .A2(new_n710), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(new_n706), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n705), .A2(new_n707), .A3(new_n710), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n716), .A3(new_n682), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n713), .A2(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G23), .ZN(new_n720));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n719), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT33), .B(G1976), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT88), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT85), .B(G16), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G22), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G166), .B2(new_n730), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(G1971), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n719), .A2(G6), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n596), .B2(new_n719), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT32), .B(G1981), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT87), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n735), .B(new_n737), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n727), .A2(new_n728), .A3(new_n733), .A4(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT34), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n489), .A2(G119), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n483), .A2(G131), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n463), .A2(G107), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n742), .B(new_n743), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G25), .B(new_n746), .S(G29), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT35), .B(G1991), .Z(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT84), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n747), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n730), .A2(G24), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n602), .A2(new_n604), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n730), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G1986), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n755), .B2(new_n754), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n741), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT36), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT36), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n741), .A2(new_n760), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g336(.A1(G160), .A2(G29), .ZN(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT24), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT92), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n623), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G4), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G35), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G162), .B2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G2090), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n769), .A2(new_n773), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n772), .B2(new_n771), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n730), .A2(G19), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n563), .B2(new_n730), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  INV_X1    g359(.A(G29), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G33), .ZN(new_n786));
  NAND2_X1  g361(.A1(G115), .A2(G2104), .ZN(new_n787));
  INV_X1    g362(.A(G127), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n477), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G2105), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT25), .Z(new_n792));
  INV_X1    g367(.A(G139), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n792), .C1(new_n793), .C2(new_n467), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n786), .B1(new_n795), .B2(new_n785), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G2072), .Z(new_n797));
  NOR2_X1   g372(.A1(G168), .A2(new_n719), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n719), .B2(G21), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1966), .ZN(new_n800));
  NOR2_X1   g375(.A1(G27), .A2(G29), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G164), .B2(G29), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n797), .B(new_n800), .C1(G2078), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n719), .A2(G5), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G171), .B2(new_n719), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n766), .A2(new_n767), .B1(new_n805), .B2(G1961), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n806), .B1(G1961), .B2(new_n805), .C1(G2090), .C2(new_n777), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n785), .A2(G32), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n464), .ZN(new_n809));
  NAND3_X1  g384(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT26), .Z(new_n811));
  INV_X1    g386(.A(G129), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n466), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n808), .B1(new_n815), .B2(new_n785), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT27), .B(G1996), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n646), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(G29), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT30), .B(G28), .ZN(new_n821));
  OR2_X1    g396(.A1(KEYINPUT31), .A2(G11), .ZN(new_n822));
  NAND2_X1  g397(.A1(KEYINPUT31), .A2(G11), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n821), .A2(new_n785), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G2078), .B2(new_n802), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n785), .A2(G26), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT28), .Z(new_n828));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n829));
  INV_X1    g404(.A(G140), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n467), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n483), .A2(KEYINPUT90), .A3(G140), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n463), .A2(G116), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT91), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n836), .B1(new_n834), .B2(new_n835), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n837), .A2(new_n838), .B1(new_n489), .B2(G128), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n833), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n828), .B1(new_n840), .B2(G29), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G2067), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n818), .A2(new_n826), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n803), .A2(new_n807), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n729), .A2(G20), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT23), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n583), .B2(new_n719), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT95), .B(G1956), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n781), .A2(new_n784), .A3(new_n844), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT96), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n844), .A2(new_n849), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n852), .A2(new_n781), .A3(new_n853), .A4(new_n784), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n759), .A2(new_n761), .B1(new_n851), .B2(new_n854), .ZN(G311));
  NAND2_X1  g430(.A1(new_n759), .A2(new_n761), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n851), .A2(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(G150));
  AOI22_X1  g433(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n519), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT97), .B(G55), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n526), .A2(new_n861), .B1(new_n535), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(KEYINPUT99), .B(G860), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n623), .A2(G559), .ZN(new_n869));
  XOR2_X1   g444(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n864), .A2(new_n558), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(new_n562), .B2(new_n864), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n871), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT39), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n868), .B1(new_n875), .B2(new_n865), .ZN(G145));
  XNOR2_X1  g451(.A(new_n746), .B(new_n637), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n489), .A2(G130), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n483), .A2(G142), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n877), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n510), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n509), .B1(new_n466), .B2(new_n506), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n503), .B(new_n502), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n840), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(G164), .A2(new_n833), .A3(new_n839), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n889), .A2(new_n794), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n794), .B1(new_n889), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n814), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n889), .A2(new_n890), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n795), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n794), .A3(new_n890), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n815), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n485), .A2(new_n486), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n646), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n899), .A2(new_n900), .A3(new_n646), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(G162), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n494), .B1(new_n905), .B2(new_n901), .ZN(new_n906));
  AOI22_X1  g481(.A1(new_n885), .A2(new_n898), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n883), .A2(new_n893), .A3(new_n897), .A4(new_n884), .ZN(new_n908));
  AOI21_X1  g483(.A(G37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n904), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n898), .B2(new_n883), .ZN(new_n911));
  INV_X1    g486(.A(new_n882), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n877), .B(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n893), .A3(new_n897), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n911), .A2(KEYINPUT101), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT101), .B1(new_n911), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n909), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g493(.A(new_n873), .B(new_n631), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n583), .A2(new_n622), .ZN(new_n921));
  AOI22_X1  g496(.A1(new_n579), .A2(new_n582), .B1(new_n616), .B2(new_n621), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n583), .A2(new_n622), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n579), .A2(new_n616), .A3(new_n582), .A4(new_n621), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(KEYINPUT41), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(KEYINPUT103), .ZN(new_n929));
  INV_X1    g504(.A(new_n919), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n924), .A2(new_n925), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(KEYINPUT103), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n752), .A2(G305), .ZN(new_n934));
  NAND2_X1  g509(.A1(G290), .A2(new_n596), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(G303), .B(G288), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n937), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT42), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n932), .A2(new_n933), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n932), .B2(new_n933), .ZN(new_n944));
  OAI21_X1  g519(.A(G868), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n860), .A2(new_n863), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(G868), .B2(new_n946), .ZN(G295));
  OAI21_X1  g522(.A(new_n945), .B1(G868), .B2(new_n946), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n539), .A2(new_n540), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(G651), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n542), .A2(new_n543), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n541), .A2(new_n544), .A3(KEYINPUT104), .ZN(new_n954));
  OAI21_X1  g529(.A(G286), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(new_n952), .A3(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT104), .B1(new_n541), .B2(new_n544), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(G168), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n946), .B1(new_n560), .B2(new_n561), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n872), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n955), .A2(new_n958), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n873), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n959), .B(KEYINPUT105), .C1(new_n960), .C2(new_n872), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n963), .A2(new_n931), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n927), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n969), .A3(new_n941), .ZN(new_n970));
  INV_X1    g545(.A(G37), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n941), .B1(new_n967), .B2(new_n969), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n970), .A2(new_n971), .ZN(new_n976));
  INV_X1    g551(.A(new_n941), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n978), .A2(new_n927), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n965), .A2(new_n931), .A3(new_n961), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n965), .A2(new_n931), .A3(new_n961), .A4(KEYINPUT106), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n977), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n976), .A2(new_n985), .A3(KEYINPUT43), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT44), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n976), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n972), .B2(new_n973), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(KEYINPUT44), .B2(new_n992), .ZN(G397));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G164), .B2(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n480), .A2(new_n484), .A3(G40), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1986), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n752), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT107), .Z(new_n1000));
  OR2_X1    g575(.A1(new_n840), .A2(G2067), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n840), .A2(G2067), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n814), .B(G1996), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n746), .B(new_n748), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1006), .B(new_n1007), .C1(new_n998), .C2(new_n752), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n997), .B1(new_n1000), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n1010));
  INV_X1    g585(.A(G1961), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n508), .A2(new_n510), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n502), .A2(new_n503), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1384), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n996), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n886), .A2(new_n887), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(new_n504), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT111), .B1(new_n1019), .B2(KEYINPUT50), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1014), .A2(new_n1021), .A3(new_n1015), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1016), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n996), .B1(new_n1019), .B2(new_n994), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n1017), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G2078), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n888), .A2(KEYINPUT108), .A3(KEYINPUT45), .A4(new_n1017), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1011), .A2(new_n1023), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1024), .A2(KEYINPUT53), .A3(new_n1028), .A4(new_n1025), .ZN(new_n1033));
  AOI21_X1  g608(.A(G301), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1023), .A2(new_n1011), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n480), .A2(new_n484), .A3(G40), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n995), .A2(new_n1036), .A3(new_n1029), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(KEYINPUT53), .A3(new_n1028), .A4(new_n1027), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1039));
  AND4_X1   g614(.A1(G301), .A2(new_n1035), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1010), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT123), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(KEYINPUT123), .B(new_n1010), .C1(new_n1034), .C2(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n888), .A2(new_n1015), .A3(new_n1017), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1036), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1021), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1019), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1966), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1051), .A2(new_n767), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT121), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1053), .A2(new_n1052), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n767), .B(new_n1016), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1055), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1046), .B1(new_n1061), .B2(G168), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n1063));
  INV_X1    g638(.A(G8), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1063), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT122), .B(new_n1066), .C1(new_n1054), .C2(new_n1064), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(G8), .ZN(new_n1071));
  OAI22_X1  g646(.A1(new_n1062), .A2(new_n1070), .B1(new_n1071), .B2(new_n1061), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1024), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT109), .B(G1971), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT110), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1078));
  INV_X1    g653(.A(G2090), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1051), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G303), .A2(G8), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT55), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1081), .A2(G8), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1981), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n596), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(G1981), .B1(new_n592), .B2(new_n595), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(KEYINPUT49), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1064), .B1(new_n1036), .B2(new_n1014), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT49), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1088), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n592), .A2(new_n595), .A3(G1981), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT113), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT113), .B(new_n1092), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G1976), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT52), .B1(G288), .B2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n587), .A2(G1976), .A3(new_n588), .A4(new_n589), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1101), .A2(new_n1090), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1036), .A2(new_n1014), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(new_n1102), .A3(G8), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1105), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT112), .B1(new_n1105), .B2(KEYINPUT52), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1103), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1099), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1019), .A2(KEYINPUT50), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1016), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G2090), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1083), .B1(new_n1113), .B2(new_n1064), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1085), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(G171), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1032), .A2(G301), .A3(new_n1033), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1117), .A2(KEYINPUT54), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1045), .A2(new_n1072), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1956), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1048), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(KEYINPUT115), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1111), .A2(new_n1126), .A3(new_n1122), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1073), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1125), .A2(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n581), .A2(new_n570), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT57), .B1(new_n1132), .B2(KEYINPUT116), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT116), .B(KEYINPUT57), .C1(new_n581), .C2(new_n570), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1130), .A2(new_n1131), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1037), .A2(new_n1027), .A3(new_n1129), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1124), .A2(KEYINPUT115), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1126), .B1(new_n1111), .B2(new_n1122), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1136), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT119), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1137), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1050), .A2(new_n1049), .ZN(new_n1146));
  AOI21_X1  g721(.A(G1348), .B1(new_n1146), .B2(new_n1016), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1104), .A2(G2067), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1148), .ZN(new_n1150));
  OAI211_X1 g725(.A(KEYINPUT118), .B(new_n1150), .C1(new_n1051), .C2(G1348), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1144), .B1(new_n622), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT117), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1141), .A2(new_n1155), .A3(new_n1142), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1153), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT58), .B(G1341), .Z(new_n1158));
  NAND2_X1  g733(.A1(new_n1104), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1073), .B2(G1996), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n563), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1144), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1167), .B1(new_n1156), .B2(new_n1154), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(new_n1164), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1149), .A2(new_n1170), .A3(new_n1151), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n623), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT120), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1173), .B1(new_n1152), .B2(KEYINPUT60), .ZN(new_n1174));
  AOI211_X1 g749(.A(KEYINPUT120), .B(new_n1170), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1152), .A2(KEYINPUT60), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT120), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1171), .A2(new_n623), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1152), .A2(new_n1173), .A3(KEYINPUT60), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1166), .A2(new_n1169), .A3(new_n1176), .A4(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1121), .B1(new_n1157), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1094), .B(KEYINPUT114), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n721), .A2(new_n1100), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n1099), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1090), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1109), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1187), .B1(new_n1085), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT63), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1065), .A2(G168), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1190), .B1(new_n1115), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1081), .A2(G8), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(new_n1083), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1191), .A2(new_n1190), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1194), .A2(new_n1085), .A3(new_n1109), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1189), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1197));
  AND4_X1   g772(.A1(new_n1034), .A2(new_n1085), .A3(new_n1114), .A4(new_n1109), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1061), .A2(new_n1071), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1070), .ZN(new_n1200));
  AND3_X1   g775(.A1(new_n1056), .A2(new_n1057), .A3(KEYINPUT121), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT121), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1202));
  OAI21_X1  g777(.A(G168), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1203), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1199), .B1(new_n1200), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1198), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1072), .A2(KEYINPUT62), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1197), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1009), .B1(new_n1183), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1000), .A2(new_n997), .ZN(new_n1211));
  XNOR2_X1  g786(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1212));
  AND2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1214));
  INV_X1    g789(.A(new_n997), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT125), .ZN(new_n1217));
  NOR3_X1   g792(.A1(new_n1213), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n997), .B1(new_n1004), .B2(new_n814), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT46), .ZN(new_n1220));
  INV_X1    g795(.A(G1996), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1220), .B1(new_n997), .B2(new_n1221), .ZN(new_n1222));
  NOR3_X1   g797(.A1(new_n1215), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1219), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  XOR2_X1   g799(.A(new_n1224), .B(KEYINPUT47), .Z(new_n1225));
  INV_X1    g800(.A(new_n748), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n746), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1006), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1215), .B1(new_n1228), .B2(new_n1001), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1229), .B(KEYINPUT124), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1218), .A2(new_n1225), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1210), .A2(new_n1231), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g807(.A(new_n680), .B(G319), .C1(new_n664), .C2(new_n665), .ZN(new_n1234));
  AOI21_X1  g808(.A(new_n1234), .B1(new_n713), .B2(new_n717), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n917), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g810(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g811(.A(KEYINPUT127), .B1(new_n991), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1239));
  AOI211_X1 g813(.A(new_n1239), .B(new_n1236), .C1(new_n989), .C2(new_n990), .ZN(new_n1240));
  NOR2_X1   g814(.A1(new_n1238), .A2(new_n1240), .ZN(G308));
  NAND2_X1  g815(.A1(new_n991), .A2(new_n1237), .ZN(G225));
endmodule


