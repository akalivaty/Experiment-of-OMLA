

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  AND2_X1 U324 ( .A1(n534), .A2(n557), .ZN(n438) );
  NOR2_X1 U325 ( .A1(n480), .A2(n590), .ZN(n481) );
  NOR2_X1 U326 ( .A1(n560), .A2(n489), .ZN(n586) );
  XOR2_X1 U327 ( .A(n447), .B(n446), .Z(n292) );
  XOR2_X1 U328 ( .A(n370), .B(n419), .Z(n293) );
  INV_X1 U329 ( .A(KEYINPUT46), .ZN(n429) );
  INV_X1 U330 ( .A(KEYINPUT75), .ZN(n411) );
  XNOR2_X1 U331 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U332 ( .A(G141GAT), .B(G22GAT), .Z(n442) );
  XNOR2_X1 U333 ( .A(n449), .B(n413), .ZN(n414) );
  XNOR2_X1 U334 ( .A(n421), .B(n420), .ZN(n422) );
  NOR2_X1 U335 ( .A1(n531), .A2(n439), .ZN(n488) );
  NOR2_X1 U336 ( .A1(n478), .A2(n477), .ZN(n496) );
  XNOR2_X1 U337 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U338 ( .A(KEYINPUT36), .B(n577), .Z(n590) );
  XNOR2_X1 U339 ( .A(n468), .B(KEYINPUT26), .ZN(n560) );
  INV_X1 U340 ( .A(G204GAT), .ZN(n490) );
  NOR2_X1 U341 ( .A1(n462), .A2(n457), .ZN(n576) );
  XNOR2_X1 U342 ( .A(n483), .B(KEYINPUT38), .ZN(n514) );
  XNOR2_X1 U343 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U344 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U345 ( .A(n493), .B(n492), .ZN(G1353GAT) );
  XNOR2_X1 U346 ( .A(n487), .B(n486), .ZN(G1328GAT) );
  XOR2_X1 U347 ( .A(G50GAT), .B(KEYINPUT68), .Z(n295) );
  XNOR2_X1 U348 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U350 ( .A(n296), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(G29GAT), .B(G36GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n379) );
  XOR2_X1 U353 ( .A(KEYINPUT29), .B(KEYINPUT65), .Z(n300) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(KEYINPUT67), .ZN(n299) );
  XNOR2_X1 U355 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n379), .B(n301), .ZN(n310) );
  XNOR2_X1 U357 ( .A(G1GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n302), .B(KEYINPUT69), .ZN(n396) );
  XOR2_X1 U359 ( .A(n442), .B(n396), .Z(n304) );
  NAND2_X1 U360 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U362 ( .A(n305), .B(KEYINPUT66), .Z(n308) );
  XNOR2_X1 U363 ( .A(G8GAT), .B(G169GAT), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n306), .B(G197GAT), .ZN(n358) );
  XNOR2_X1 U365 ( .A(n358), .B(KEYINPUT30), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n580) );
  XNOR2_X1 U368 ( .A(n580), .B(KEYINPUT70), .ZN(n547) );
  XOR2_X1 U369 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n312) );
  XNOR2_X1 U370 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n311) );
  XNOR2_X1 U371 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U372 ( .A(G120GAT), .B(G71GAT), .Z(n418) );
  XOR2_X1 U373 ( .A(n313), .B(n418), .Z(n315) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G99GAT), .ZN(n314) );
  XNOR2_X1 U375 ( .A(n315), .B(n314), .ZN(n320) );
  XOR2_X1 U376 ( .A(G134GAT), .B(G190GAT), .Z(n367) );
  XNOR2_X1 U377 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n316), .B(G127GAT), .ZN(n344) );
  XOR2_X1 U379 ( .A(n367), .B(n344), .Z(n318) );
  NAND2_X1 U380 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U382 ( .A(n320), .B(n319), .Z(n328) );
  XOR2_X1 U383 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n322) );
  XNOR2_X1 U384 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U386 ( .A(G183GAT), .B(n323), .Z(n355) );
  XOR2_X1 U387 ( .A(G169GAT), .B(G176GAT), .Z(n325) );
  XNOR2_X1 U388 ( .A(KEYINPUT88), .B(KEYINPUT64), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U390 ( .A(n355), .B(n326), .ZN(n327) );
  XOR2_X1 U391 ( .A(n328), .B(n327), .Z(n462) );
  XOR2_X1 U392 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n330) );
  XNOR2_X1 U393 ( .A(KEYINPUT93), .B(KEYINPUT4), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n330), .B(n329), .ZN(n348) );
  XOR2_X1 U395 ( .A(G148GAT), .B(G120GAT), .Z(n332) );
  XNOR2_X1 U396 ( .A(G162GAT), .B(G134GAT), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U398 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n334) );
  XNOR2_X1 U399 ( .A(G141GAT), .B(G57GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U401 ( .A(n336), .B(n335), .Z(n342) );
  XNOR2_X1 U402 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n337), .B(KEYINPUT3), .ZN(n452) );
  XOR2_X1 U404 ( .A(G85GAT), .B(n452), .Z(n339) );
  NAND2_X1 U405 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U406 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(n340), .ZN(n341) );
  XNOR2_X1 U408 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U409 ( .A(n343), .B(KEYINPUT1), .Z(n346) );
  XNOR2_X1 U410 ( .A(n344), .B(G1GAT), .ZN(n345) );
  XNOR2_X1 U411 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n474) );
  INV_X1 U413 ( .A(n474), .ZN(n531) );
  XOR2_X1 U414 ( .A(KEYINPUT95), .B(KEYINPUT98), .Z(n350) );
  XNOR2_X1 U415 ( .A(KEYINPUT82), .B(KEYINPUT96), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U417 ( .A(KEYINPUT97), .B(n351), .ZN(n353) );
  AND2_X1 U418 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U419 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U420 ( .A(n355), .B(n354), .Z(n357) );
  XNOR2_X1 U421 ( .A(G36GAT), .B(G190GAT), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n366) );
  XNOR2_X1 U424 ( .A(G204GAT), .B(KEYINPUT90), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n360), .B(KEYINPUT21), .ZN(n361) );
  XOR2_X1 U426 ( .A(n361), .B(KEYINPUT89), .Z(n363) );
  XNOR2_X1 U427 ( .A(G218GAT), .B(G211GAT), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n451) );
  XNOR2_X1 U429 ( .A(G92GAT), .B(G64GAT), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n364), .B(G176GAT), .ZN(n416) );
  XNOR2_X1 U431 ( .A(n451), .B(n416), .ZN(n365) );
  XNOR2_X1 U432 ( .A(n366), .B(n365), .ZN(n534) );
  XOR2_X1 U433 ( .A(G162GAT), .B(KEYINPUT79), .Z(n443) );
  XOR2_X1 U434 ( .A(n443), .B(n367), .Z(n369) );
  NAND2_X1 U435 ( .A1(G232GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(G85GAT), .B(G99GAT), .Z(n419) );
  XOR2_X1 U438 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n372) );
  XNOR2_X1 U439 ( .A(G218GAT), .B(G106GAT), .ZN(n371) );
  XNOR2_X1 U440 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U441 ( .A(KEYINPUT81), .B(KEYINPUT9), .Z(n374) );
  XNOR2_X1 U442 ( .A(G92GAT), .B(KEYINPUT80), .ZN(n373) );
  XNOR2_X1 U443 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U444 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n293), .B(n377), .ZN(n378) );
  XOR2_X1 U446 ( .A(n379), .B(n378), .Z(n577) );
  XOR2_X1 U447 ( .A(G78GAT), .B(G183GAT), .Z(n381) );
  XNOR2_X1 U448 ( .A(G127GAT), .B(G71GAT), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U450 ( .A(G64GAT), .B(G211GAT), .Z(n383) );
  XNOR2_X1 U451 ( .A(G155GAT), .B(G22GAT), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U453 ( .A(n385), .B(n384), .Z(n390) );
  XOR2_X1 U454 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n387) );
  NAND2_X1 U455 ( .A1(G231GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U457 ( .A(KEYINPUT15), .B(n388), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U459 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n392) );
  XNOR2_X1 U460 ( .A(G8GAT), .B(KEYINPUT82), .ZN(n391) );
  XNOR2_X1 U461 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U462 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U463 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n395), .B(KEYINPUT13), .ZN(n417) );
  XNOR2_X1 U465 ( .A(n417), .B(n396), .ZN(n397) );
  XOR2_X1 U466 ( .A(n398), .B(n397), .Z(n494) );
  NOR2_X1 U467 ( .A1(n590), .A2(n494), .ZN(n400) );
  XNOR2_X1 U468 ( .A(KEYINPUT45), .B(KEYINPUT116), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n426) );
  XOR2_X1 U470 ( .A(KEYINPUT32), .B(KEYINPUT72), .Z(n402) );
  XNOR2_X1 U471 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n402), .B(n401), .ZN(n425) );
  XOR2_X1 U473 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n404) );
  XNOR2_X1 U474 ( .A(G204GAT), .B(KEYINPUT73), .ZN(n403) );
  XNOR2_X1 U475 ( .A(n404), .B(n403), .ZN(n415) );
  INV_X1 U476 ( .A(KEYINPUT74), .ZN(n405) );
  NAND2_X1 U477 ( .A1(n405), .A2(G78GAT), .ZN(n408) );
  INV_X1 U478 ( .A(G78GAT), .ZN(n406) );
  NAND2_X1 U479 ( .A1(n406), .A2(KEYINPUT74), .ZN(n407) );
  NAND2_X1 U480 ( .A1(n408), .A2(n407), .ZN(n410) );
  XNOR2_X1 U481 ( .A(G148GAT), .B(G106GAT), .ZN(n409) );
  XNOR2_X1 U482 ( .A(n410), .B(n409), .ZN(n449) );
  NAND2_X1 U483 ( .A1(G230GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U484 ( .A(n415), .B(n414), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U486 ( .A(n419), .B(n418), .Z(n420) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n428) );
  NAND2_X1 U488 ( .A1(n426), .A2(n428), .ZN(n427) );
  NOR2_X1 U489 ( .A1(n547), .A2(n427), .ZN(n436) );
  XNOR2_X1 U490 ( .A(KEYINPUT41), .B(n428), .ZN(n572) );
  NAND2_X1 U491 ( .A1(n572), .A2(n580), .ZN(n430) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n433) );
  INV_X1 U493 ( .A(n577), .ZN(n431) );
  NAND2_X1 U494 ( .A1(n431), .A2(n494), .ZN(n432) );
  NOR2_X1 U495 ( .A1(n433), .A2(n432), .ZN(n434) );
  XOR2_X1 U496 ( .A(n434), .B(KEYINPUT47), .Z(n435) );
  NOR2_X1 U497 ( .A1(n436), .A2(n435), .ZN(n437) );
  XOR2_X1 U498 ( .A(n437), .B(KEYINPUT48), .Z(n557) );
  XOR2_X1 U499 ( .A(KEYINPUT54), .B(n438), .Z(n439) );
  XOR2_X1 U500 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n441) );
  XNOR2_X1 U501 ( .A(G197GAT), .B(KEYINPUT23), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n447) );
  XOR2_X1 U503 ( .A(KEYINPUT22), .B(n442), .Z(n445) );
  XNOR2_X1 U504 ( .A(G50GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  NAND2_X1 U506 ( .A1(G228GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n292), .B(n448), .ZN(n450) );
  XOR2_X1 U508 ( .A(n450), .B(n449), .Z(n454) );
  XNOR2_X1 U509 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U510 ( .A(n454), .B(n453), .ZN(n475) );
  NAND2_X1 U511 ( .A1(n488), .A2(n475), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U514 ( .A1(n547), .A2(n576), .ZN(n460) );
  INV_X1 U515 ( .A(G169GAT), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(KEYINPUT121), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n460), .B(n459), .ZN(G1348GAT) );
  NAND2_X1 U518 ( .A1(n547), .A2(n428), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT78), .ZN(n499) );
  INV_X1 U520 ( .A(n462), .ZN(n544) );
  NAND2_X1 U521 ( .A1(n544), .A2(n534), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT100), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n464), .A2(n475), .ZN(n466) );
  XOR2_X1 U524 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n465) );
  XNOR2_X1 U525 ( .A(n466), .B(n465), .ZN(n470) );
  XOR2_X1 U526 ( .A(n534), .B(KEYINPUT27), .Z(n473) );
  NOR2_X1 U527 ( .A1(n544), .A2(n475), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n467), .B(KEYINPUT99), .ZN(n468) );
  NOR2_X1 U529 ( .A1(n473), .A2(n560), .ZN(n469) );
  NOR2_X1 U530 ( .A1(n470), .A2(n469), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n471), .A2(n531), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT102), .ZN(n478) );
  NOR2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n558) );
  XOR2_X1 U534 ( .A(n475), .B(KEYINPUT28), .Z(n537) );
  INV_X1 U535 ( .A(n537), .ZN(n476) );
  NAND2_X1 U536 ( .A1(n558), .A2(n476), .ZN(n543) );
  NOR2_X1 U537 ( .A1(n543), .A2(n544), .ZN(n477) );
  INV_X1 U538 ( .A(n494), .ZN(n585) );
  NOR2_X1 U539 ( .A1(n496), .A2(n585), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT107), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT108), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(KEYINPUT37), .ZN(n530) );
  NOR2_X1 U543 ( .A1(n499), .A2(n530), .ZN(n483) );
  NAND2_X1 U544 ( .A1(n531), .A2(n514), .ZN(n487) );
  XOR2_X1 U545 ( .A(KEYINPUT39), .B(KEYINPUT109), .Z(n485) );
  INV_X1 U546 ( .A(G29GAT), .ZN(n484) );
  INV_X1 U547 ( .A(n488), .ZN(n489) );
  INV_X1 U548 ( .A(n586), .ZN(n589) );
  OR2_X1 U549 ( .A1(n589), .A2(n428), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n491) );
  XOR2_X1 U551 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n501) );
  NOR2_X1 U552 ( .A1(n577), .A2(n494), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(KEYINPUT16), .ZN(n498) );
  INV_X1 U554 ( .A(n496), .ZN(n497) );
  NAND2_X1 U555 ( .A1(n498), .A2(n497), .ZN(n518) );
  NOR2_X1 U556 ( .A1(n499), .A2(n518), .ZN(n507) );
  NAND2_X1 U557 ( .A1(n507), .A2(n531), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U559 ( .A(G1GAT), .B(n502), .ZN(G1324GAT) );
  NAND2_X1 U560 ( .A1(n534), .A2(n507), .ZN(n503) );
  XNOR2_X1 U561 ( .A(n503), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U563 ( .A1(n507), .A2(n544), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G15GAT), .B(n506), .ZN(G1326GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n509) );
  NAND2_X1 U567 ( .A1(n507), .A2(n537), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U569 ( .A(G22GAT), .B(n510), .ZN(G1327GAT) );
  NAND2_X1 U570 ( .A1(n514), .A2(n534), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n511), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n514), .A2(n544), .ZN(n512) );
  XNOR2_X1 U573 ( .A(n512), .B(KEYINPUT40), .ZN(n513) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n513), .ZN(G1330GAT) );
  NAND2_X1 U575 ( .A1(n514), .A2(n537), .ZN(n515) );
  XNOR2_X1 U576 ( .A(n515), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n521) );
  INV_X1 U578 ( .A(n572), .ZN(n516) );
  NOR2_X1 U579 ( .A1(n580), .A2(n516), .ZN(n517) );
  XOR2_X1 U580 ( .A(KEYINPUT110), .B(n517), .Z(n529) );
  NOR2_X1 U581 ( .A1(n529), .A2(n518), .ZN(n519) );
  XOR2_X1 U582 ( .A(KEYINPUT111), .B(n519), .Z(n525) );
  NAND2_X1 U583 ( .A1(n525), .A2(n531), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NAND2_X1 U586 ( .A1(n534), .A2(n525), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n544), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U591 ( .A1(n525), .A2(n537), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(G78GAT), .B(n528), .Z(G1335GAT) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(KEYINPUT114), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n531), .A2(n538), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n538), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n544), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n540) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U605 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  INV_X1 U606 ( .A(n557), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n545) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT117), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n547), .A2(n554), .ZN(n548) );
  XNOR2_X1 U611 ( .A(n548), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n550) );
  NAND2_X1 U613 ( .A1(n554), .A2(n572), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G120GAT), .B(n551), .ZN(G1341GAT) );
  NAND2_X1 U616 ( .A1(n554), .A2(n585), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n552), .B(KEYINPUT50), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(n553), .ZN(G1342GAT) );
  XOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U620 ( .A1(n554), .A2(n577), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(G1343GAT) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U623 ( .A1(n560), .A2(n559), .ZN(n567) );
  NAND2_X1 U624 ( .A1(n580), .A2(n567), .ZN(n561) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n561), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n563) );
  NAND2_X1 U627 ( .A1(n567), .A2(n572), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(G148GAT), .B(KEYINPUT53), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n585), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n577), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n570) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT122), .B(n571), .Z(n574) );
  NAND2_X1 U639 ( .A1(n572), .A2(n576), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n585), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U643 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1351GAT) );
  NAND2_X1 U646 ( .A1(n586), .A2(n580), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n582) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT126), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

