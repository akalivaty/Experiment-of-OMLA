//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G197gat), .B(G204gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n210), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g015(.A1(new_n212), .A2(KEYINPUT73), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n217), .A2(new_n209), .A3(new_n211), .A4(new_n213), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(KEYINPUT74), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n220), .B(new_n210), .C1(new_n214), .C2(new_n215), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n208), .B1(new_n222), .B2(KEYINPUT29), .ZN(new_n223));
  AND2_X1   g022(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT2), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G148gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT78), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G148gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n232), .A3(G141gat), .ZN(new_n233));
  INV_X1    g032(.A(G141gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G148gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G155gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n227), .ZN(new_n238));
  NAND2_X1  g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n228), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n229), .A2(G141gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(KEYINPUT2), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n239), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n237), .A3(new_n227), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT77), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n245), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n249), .ZN(new_n253));
  NOR3_X1   g052(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n239), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT77), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n241), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n207), .B1(new_n223), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(KEYINPUT77), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(new_n251), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n245), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(new_n208), .A3(new_n241), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n222), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT80), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n267), .A3(new_n222), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n258), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n265), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n255), .A2(KEYINPUT77), .B1(new_n244), .B2(new_n243), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n233), .A2(new_n235), .B1(new_n239), .B2(new_n238), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n271), .A2(new_n260), .B1(new_n228), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n216), .A2(new_n218), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n263), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n275), .B2(new_n208), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n207), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G22gat), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n269), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n269), .B2(new_n277), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n206), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n269), .A2(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G22gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n269), .A2(new_n277), .A3(new_n278), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n205), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G190gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(G183gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT27), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G183gat), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n288), .A2(new_n290), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT66), .B(G190gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n297), .A2(new_n298), .A3(new_n302), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n291), .A2(new_n287), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n303), .A2(KEYINPUT23), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G169gat), .B2(G176gat), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT64), .A4(new_n311), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n315), .A2(new_n320), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n291), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n299), .A2(new_n291), .B1(G190gat), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT65), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n298), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n309), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n324), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n308), .B(new_n323), .C1(new_n331), .C2(new_n321), .ZN(new_n332));
  AND2_X1   g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n332), .A2(new_n263), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n222), .B(new_n334), .C1(new_n335), .C2(new_n333), .ZN(new_n336));
  INV_X1    g135(.A(new_n222), .ZN(new_n337));
  INV_X1    g136(.A(new_n334), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n333), .B1(new_n332), .B2(new_n263), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(KEYINPUT75), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n344), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n336), .B2(new_n340), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT30), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n340), .A3(new_n348), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n347), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n354));
  INV_X1    g153(.A(G120gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G113gat), .ZN(new_n356));
  INV_X1    g155(.A(G113gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G120gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT69), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n356), .A2(new_n358), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n361), .ZN(new_n366));
  INV_X1    g165(.A(new_n363), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT68), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT1), .B1(new_n356), .B2(new_n358), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT68), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n369), .A2(new_n370), .A3(new_n363), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n364), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n262), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n257), .B2(new_n372), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n366), .A2(KEYINPUT68), .A3(new_n367), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n370), .B1(new_n369), .B2(new_n363), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n363), .A2(new_n361), .A3(new_n362), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n377), .A2(new_n378), .B1(new_n379), .B2(new_n360), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n273), .A2(KEYINPUT4), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n373), .A2(new_n374), .A3(new_n376), .A4(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n257), .A2(new_n372), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n377), .A2(new_n378), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n261), .A2(new_n385), .A3(new_n241), .A4(new_n364), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n374), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n383), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n376), .A2(new_n381), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(new_n383), .A3(new_n374), .A4(new_n373), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G1gat), .B(G29gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT0), .ZN(new_n395));
  XNOR2_X1  g194(.A(G57gat), .B(G85gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n390), .A2(new_n392), .A3(new_n397), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n202), .A2(new_n286), .A3(new_n353), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n332), .A2(new_n380), .ZN(new_n406));
  AND2_X1   g205(.A1(G227gat), .A2(G233gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n330), .A2(new_n408), .A3(new_n311), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n320), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT25), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n372), .A2(new_n411), .A3(new_n323), .A4(new_n308), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(KEYINPUT32), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT70), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n413), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n413), .A2(new_n417), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n416), .B1(new_n413), .B2(KEYINPUT32), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n421), .A2(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n407), .B1(new_n406), .B2(new_n412), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT34), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT72), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n421), .A2(new_n422), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n424), .A2(new_n423), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n425), .A2(new_n427), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n428), .B1(new_n435), .B2(KEYINPUT72), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n405), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n435), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(new_n286), .A3(new_n353), .A4(new_n404), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT35), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n433), .A2(KEYINPUT36), .A3(new_n434), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT71), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n433), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n434), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n429), .A2(new_n427), .A3(new_n430), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n427), .B1(new_n429), .B2(new_n430), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT72), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n428), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT36), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n281), .A2(new_n285), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n402), .A2(new_n403), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n347), .A2(new_n352), .A3(new_n351), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n336), .A2(new_n340), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n457), .B1(new_n336), .B2(new_n340), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n348), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT38), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT38), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(new_n348), .C1(new_n458), .C2(new_n459), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n463), .A3(new_n345), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n464), .A2(new_n404), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT40), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n354), .A2(new_n262), .A3(new_n372), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n376), .A2(new_n381), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n388), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n384), .A2(new_n386), .A3(new_n374), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT39), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT81), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n473), .A3(KEYINPUT39), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT39), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n476), .B(new_n388), .C1(new_n467), .C2(new_n468), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n397), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n466), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(KEYINPUT40), .A3(new_n397), .A4(new_n477), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n399), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n286), .B1(new_n353), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n456), .B1(new_n465), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n441), .B1(new_n452), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G113gat), .B(G141gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G197gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT11), .B(G169gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G15gat), .B(G22gat), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(G1gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n495), .B2(G1gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(G8gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n494), .B(new_n496), .C1(new_n498), .C2(G8gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n507), .B1(G29gat), .B2(G36gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(G29gat), .A2(G36gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n512));
  INV_X1    g311(.A(G43gat), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n513), .A2(G50gat), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT15), .B1(new_n513), .B2(G50gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n511), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n510), .A2(KEYINPUT83), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT84), .B(G50gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n513), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT85), .B1(new_n513), .B2(G50gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n511), .B1(new_n521), .B2(KEYINPUT85), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n517), .B(new_n518), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n503), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n521), .B(KEYINPUT85), .C1(new_n513), .C2(G50gat), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n519), .A4(new_n511), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(KEYINPUT17), .A3(new_n517), .A4(new_n518), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n527), .B1(new_n534), .B2(new_n503), .ZN(new_n535));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(KEYINPUT18), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n536), .B(KEYINPUT13), .Z(new_n538));
  AND2_X1   g337(.A1(new_n503), .A2(new_n526), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(new_n527), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(new_n535), .B2(new_n536), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n492), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n535), .A2(new_n536), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n542), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n547), .A2(new_n491), .A3(new_n537), .A4(new_n540), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n548), .A3(KEYINPUT88), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT88), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n550), .B(new_n492), .C1(new_n541), .C2(new_n544), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT92), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT41), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(G85gat), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT8), .A2(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n558), .B2(new_n559), .ZN(new_n562));
  NAND3_X1  g361(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G99gat), .B(G106gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n556), .B1(new_n526), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT94), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n569), .B(new_n556), .C1(new_n526), .C2(new_n566), .ZN(new_n570));
  AOI22_X1  g369(.A1(new_n568), .A2(new_n570), .B1(new_n534), .B2(new_n566), .ZN(new_n571));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT95), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n573), .ZN(new_n577));
  XOR2_X1   g376(.A(G134gat), .B(G162gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT93), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n555), .A2(KEYINPUT41), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  NAND4_X1  g380(.A1(new_n575), .A2(new_n576), .A3(new_n577), .A4(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n577), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n576), .B1(new_n571), .B2(new_n573), .ZN(new_n584));
  INV_X1    g383(.A(new_n581), .ZN(new_n585));
  OAI22_X1  g384(.A1(new_n583), .A2(new_n574), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  INV_X1    g388(.A(G78gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n590), .ZN(new_n593));
  XNOR2_X1  g392(.A(G57gat), .B(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(new_n595), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT89), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G57gat), .ZN(new_n600));
  OAI22_X1  g399(.A1(new_n597), .A2(new_n591), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n598), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n596), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT21), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n503), .B1(new_n605), .B2(new_n604), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT20), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n613), .B(KEYINPUT90), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G183gat), .B(G211gat), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n610), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n588), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G230gat), .ZN(new_n620));
  INV_X1    g419(.A(G233gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n566), .A2(new_n604), .ZN(new_n623));
  OAI221_X1 g422(.A(new_n602), .B1(new_n598), .B2(new_n600), .C1(new_n591), .C2(new_n597), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n564), .A2(new_n565), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n564), .A2(new_n565), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .A4(new_n596), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT10), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n623), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OR3_X1    g428(.A1(new_n566), .A2(new_n628), .A3(new_n604), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n622), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI211_X1 g430(.A(new_n620), .B(new_n621), .C1(new_n623), .C2(new_n627), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT96), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n633), .A2(KEYINPUT96), .A3(new_n637), .ZN(new_n640));
  AND2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n619), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n485), .A2(new_n553), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT97), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n454), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT98), .B(G1gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1324gat));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G8gat), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n644), .A2(new_n455), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n500), .B1(new_n644), .B2(new_n455), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT42), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n652), .B1(KEYINPUT42), .B2(new_n650), .ZN(G1325gat));
  INV_X1    g452(.A(G15gat), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n644), .A2(new_n654), .A3(new_n436), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n644), .A2(new_n452), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n654), .ZN(G1326gat));
  NAND2_X1  g456(.A1(new_n644), .A2(new_n453), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  AND2_X1   g459(.A1(new_n485), .A2(new_n553), .ZN(new_n661));
  INV_X1    g460(.A(new_n641), .ZN(new_n662));
  INV_X1    g461(.A(new_n618), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n587), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n664), .B(KEYINPUT100), .Z(new_n665));
  NAND4_X1  g464(.A1(new_n661), .A2(new_n504), .A3(new_n454), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n618), .B(KEYINPUT102), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n553), .A2(new_n662), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n670), .B(KEYINPUT103), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n452), .A2(new_n484), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n286), .B1(new_n404), .B2(new_n353), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n454), .A2(new_n463), .A3(new_n345), .A4(new_n461), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n479), .A2(new_n399), .A3(new_n481), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n677), .A2(new_n455), .B1(new_n285), .B2(new_n281), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n675), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n445), .B(new_n444), .C1(new_n436), .C2(KEYINPUT36), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT104), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n441), .B1(new_n674), .B2(new_n681), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n587), .A3(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n485), .B2(new_n587), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n672), .B1(new_n684), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n504), .B1(new_n688), .B2(new_n454), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n668), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n668), .B2(new_n689), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1328gat));
  NAND2_X1  g492(.A1(new_n688), .A2(new_n455), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n505), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n695), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n661), .A2(new_n665), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n698), .A2(G36gat), .A3(new_n353), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n688), .A2(G43gat), .A3(new_n452), .ZN(new_n702));
  INV_X1    g501(.A(new_n436), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n513), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n405), .A2(new_n436), .B1(new_n439), .B2(KEYINPUT35), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n673), .B1(new_n452), .B2(new_n484), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n679), .A2(KEYINPUT104), .A3(new_n680), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n683), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n588), .A3(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n453), .B(new_n671), .C1(new_n713), .C2(new_n686), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n707), .B1(new_n714), .B2(new_n520), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n286), .A2(new_n520), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n698), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(new_n714), .B2(new_n520), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n715), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI221_X4 g519(.A(new_n717), .B1(new_n707), .B2(KEYINPUT48), .C1(new_n714), .C2(new_n520), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(G1331gat));
  NOR4_X1   g521(.A1(new_n711), .A2(new_n553), .A3(new_n619), .A4(new_n662), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n454), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n455), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT49), .B(G64gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n723), .A2(new_n455), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1333gat));
  AOI21_X1  g531(.A(new_n589), .B1(new_n723), .B2(new_n452), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n703), .A2(G71gat), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n723), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n723), .A2(new_n453), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g537(.A1(new_n553), .A2(new_n618), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n641), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT110), .Z(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n713), .B2(new_n686), .ZN(new_n742));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742), .B2(new_n404), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n682), .A2(new_n587), .A3(new_n739), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n454), .A2(new_n558), .A3(new_n641), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n742), .B2(new_n353), .ZN(new_n751));
  INV_X1    g550(.A(new_n741), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n684), .B2(new_n687), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(KEYINPUT112), .A3(new_n455), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n754), .A3(G92gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n662), .A2(new_n353), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(G92gat), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(new_n746), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n744), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n744), .B2(KEYINPUT111), .ZN(new_n762));
  INV_X1    g561(.A(new_n758), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n559), .B1(new_n753), .B2(new_n455), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n766), .ZN(G1337gat));
  OAI21_X1  g566(.A(G99gat), .B1(new_n742), .B2(new_n680), .ZN(new_n768));
  OR3_X1    g567(.A1(new_n703), .A2(G99gat), .A3(new_n662), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n768), .B1(new_n747), .B2(new_n769), .ZN(G1338gat));
  NOR3_X1   g569(.A1(new_n662), .A2(new_n286), .A3(G106gat), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n761), .A2(new_n762), .A3(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT113), .B(G106gat), .Z(new_n774));
  AOI21_X1  g573(.A(new_n774), .B1(new_n753), .B2(new_n453), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT53), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n747), .B2(new_n772), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(new_n775), .ZN(G1339gat));
  INV_X1    g578(.A(new_n489), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n535), .A2(new_n536), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n539), .A2(new_n527), .A3(new_n538), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n548), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n633), .A2(new_n638), .ZN(new_n785));
  AND3_X1   g584(.A1(new_n629), .A2(new_n630), .A3(new_n622), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n786), .A2(new_n631), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  AOI211_X1 g588(.A(KEYINPUT54), .B(new_n622), .C1(new_n629), .C2(new_n630), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(new_n637), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n631), .A2(new_n787), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(KEYINPUT114), .A3(new_n638), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n788), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n785), .B1(new_n794), .B2(KEYINPUT55), .ZN(new_n795));
  INV_X1    g594(.A(new_n788), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n790), .A2(new_n789), .A3(new_n637), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT114), .B1(new_n792), .B2(new_n638), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND4_X1   g600(.A1(new_n587), .A2(new_n784), .A3(new_n795), .A4(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n549), .A2(new_n795), .A3(new_n551), .A4(new_n801), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n784), .A2(new_n641), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n802), .B1(new_n805), .B2(new_n588), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT115), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n587), .B1(new_n803), .B2(new_n804), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n802), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n807), .A2(new_n669), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n642), .A2(new_n552), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n404), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n438), .A2(new_n286), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n455), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n552), .A2(G113gat), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT118), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n453), .B1(new_n811), .B2(new_n812), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n454), .A2(new_n353), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n703), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT116), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n820), .A2(new_n825), .A3(new_n822), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n553), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n827), .A2(KEYINPUT117), .A3(G113gat), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT117), .B1(new_n827), .B2(G113gat), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n819), .B1(new_n828), .B2(new_n829), .ZN(G1340gat));
  AOI21_X1  g629(.A(G120gat), .B1(new_n816), .B2(new_n641), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n824), .A2(new_n826), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n662), .A2(new_n355), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(G1341gat));
  INV_X1    g633(.A(G127gat), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n835), .A3(new_n618), .ZN(new_n836));
  INV_X1    g635(.A(new_n669), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n838), .B2(new_n835), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n816), .A2(new_n840), .A3(new_n587), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n832), .A2(new_n587), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n840), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n452), .A2(new_n821), .ZN(new_n846));
  XNOR2_X1  g645(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n810), .A2(new_n669), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n809), .A2(new_n808), .A3(new_n802), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n812), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(new_n453), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n453), .A2(KEYINPUT57), .ZN(new_n853));
  XNOR2_X1  g652(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n799), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT121), .B1(new_n795), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n552), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n795), .A2(new_n855), .A3(KEYINPUT121), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n587), .B1(new_n859), .B2(new_n804), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n663), .B1(new_n860), .B2(new_n802), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n853), .B1(new_n861), .B2(new_n812), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n553), .B(new_n846), .C1(new_n852), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G141gat), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n452), .A2(new_n286), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n813), .A2(new_n353), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n552), .A2(G141gat), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n866), .A2(new_n867), .B1(KEYINPUT122), .B2(KEYINPUT58), .ZN(new_n868));
  OR2_X1    g667(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n864), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1344gat));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n812), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n861), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n453), .ZN(new_n876));
  AOI211_X1 g675(.A(new_n286), .B(new_n847), .C1(new_n811), .C2(new_n812), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n846), .A2(new_n641), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT59), .B(G148gat), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n852), .A2(new_n862), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n641), .A4(new_n846), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n866), .B2(new_n641), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n230), .A2(new_n232), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n880), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(G1345gat));
  NAND3_X1  g685(.A1(new_n866), .A2(new_n226), .A3(new_n618), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n881), .A2(new_n846), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n669), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n226), .ZN(G1346gat));
  NOR3_X1   g689(.A1(new_n888), .A2(new_n227), .A3(new_n588), .ZN(new_n891));
  AOI21_X1  g690(.A(G162gat), .B1(new_n866), .B2(new_n587), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n814), .A2(new_n353), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n851), .A2(new_n404), .A3(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(G169gat), .B1(new_n896), .B2(new_n553), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n404), .A2(new_n455), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n703), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n851), .A2(new_n286), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT124), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n820), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n553), .A2(G169gat), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(G1348gat));
  NAND4_X1  g705(.A1(new_n901), .A2(new_n903), .A3(G176gat), .A4(new_n641), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n907), .A2(KEYINPUT125), .ZN(new_n909));
  AOI21_X1  g708(.A(G176gat), .B1(new_n896), .B2(new_n641), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(G1349gat));
  NAND3_X1  g710(.A1(new_n901), .A2(new_n903), .A3(new_n837), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G183gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT127), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(KEYINPUT127), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n618), .A2(new_n300), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n895), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n454), .B1(new_n811), .B2(new_n812), .ZN(new_n920));
  INV_X1    g719(.A(new_n918), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n920), .A2(KEYINPUT126), .A3(new_n894), .A4(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n916), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n913), .A2(new_n915), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n915), .B1(new_n913), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1350gat));
  NAND3_X1  g725(.A1(new_n896), .A2(new_n299), .A3(new_n587), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n901), .A2(new_n903), .A3(new_n587), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n928), .A2(new_n929), .A3(G190gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n928), .B2(G190gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G1351gat));
  AND2_X1   g731(.A1(new_n920), .A2(new_n865), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(new_n455), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n553), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n878), .A2(new_n452), .A3(new_n898), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n553), .A2(G197gat), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(G1352gat));
  OR2_X1    g737(.A1(new_n876), .A2(new_n877), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n452), .A2(new_n898), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n641), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G204gat), .ZN(new_n942));
  INV_X1    g741(.A(G204gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n933), .A2(new_n943), .A3(new_n756), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n944), .A2(KEYINPUT62), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(G1353gat));
  INV_X1    g746(.A(G211gat), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n934), .A2(new_n948), .A3(new_n618), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n618), .B(new_n940), .C1(new_n876), .C2(new_n877), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  NAND3_X1  g752(.A1(new_n939), .A2(new_n587), .A3(new_n940), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G218gat), .ZN(new_n955));
  INV_X1    g754(.A(G218gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n934), .A2(new_n956), .A3(new_n587), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1355gat));
endmodule


