//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n620, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1208, new_n1209,
    new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT67), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n467), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n462), .A2(G2105), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n476), .A2(G2105), .B1(G101), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND4_X1  g055(.A1(new_n463), .A2(new_n466), .A3(G2105), .A4(new_n467), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n481), .A2(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n463), .A2(new_n466), .A3(new_n483), .A4(new_n467), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(G136), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n473), .A2(new_n467), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n492), .A2(KEYINPUT4), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G114), .C2(new_n483), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n481), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n495), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n502), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n509), .A2(new_n517), .ZN(G166));
  AOI22_X1  g093(.A1(new_n503), .A2(new_n505), .B1(new_n510), .B2(new_n511), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(G89), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n512), .A2(G51), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n526));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n506), .B2(new_n528), .ZN(new_n529));
  AOI211_X1 g104(.A(KEYINPUT70), .B(new_n527), .C1(new_n503), .C2(new_n505), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n533), .B(new_n525), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n524), .B1(new_n532), .B2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n508), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n512), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n515), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n508), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n519), .A2(G81), .B1(new_n512), .B2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  NOR2_X1   g127(.A1(KEYINPUT73), .A2(G65), .ZN(new_n553));
  AND2_X1   g128(.A1(KEYINPUT73), .A2(G65), .ZN(new_n554));
  AOI211_X1 g129(.A(new_n553), .B(new_n554), .C1(new_n503), .C2(new_n505), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n552), .B(G651), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n553), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n556), .B1(new_n506), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(KEYINPUT74), .B1(new_n559), .B2(new_n508), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n506), .A2(G91), .A3(new_n514), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n519), .A2(KEYINPUT72), .A3(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n514), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n512), .A2(new_n569), .A3(G53), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n564), .A2(new_n565), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n561), .A2(new_n571), .ZN(G299));
  XNOR2_X1  g147(.A(G171), .B(KEYINPUT75), .ZN(G301));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  NOR2_X1   g149(.A1(G168), .A2(new_n574), .ZN(new_n575));
  AOI211_X1 g150(.A(KEYINPUT76), .B(new_n524), .C1(new_n532), .C2(new_n534), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n519), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n512), .A2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(new_n506), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(KEYINPUT77), .A3(G651), .ZN(new_n590));
  INV_X1    g165(.A(G48), .ZN(new_n591));
  OAI21_X1  g166(.A(KEYINPUT78), .B1(new_n566), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n512), .A2(new_n593), .A3(G48), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n592), .A2(new_n594), .B1(G86), .B2(new_n519), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n589), .A2(new_n590), .A3(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n508), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n519), .A2(G85), .B1(new_n512), .B2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n598), .A2(KEYINPUT79), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(new_n512), .A2(G54), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(new_n503), .B2(new_n505), .ZN(new_n607));
  AND2_X1   g182(.A1(G79), .A2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(G651), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND3_X1   g184(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  AOI21_X1  g185(.A(KEYINPUT10), .B1(new_n519), .B2(G92), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n605), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n614));
  XNOR2_X1  g189(.A(G171), .B(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(G868), .ZN(G321));
  XOR2_X1   g191(.A(G321), .B(KEYINPUT80), .Z(G284));
  MUX2_X1   g192(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g193(.A(G280), .B(KEYINPUT81), .ZN(G297));
  INV_X1    g194(.A(new_n612), .ZN(new_n620));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g201(.A1(new_n493), .A2(new_n477), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n483), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n481), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n488), .B2(G135), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n630), .A2(new_n637), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n650), .B(new_n651), .Z(new_n652));
  OR2_X1    g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n649), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n658), .B2(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n659), .B2(new_n660), .ZN(new_n664));
  INV_X1    g239(.A(new_n660), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n665), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n662), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(KEYINPUT84), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n683), .B2(new_n684), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT85), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n683), .A2(new_n684), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n680), .B(KEYINPUT19), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n685), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n696), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n690), .A2(new_n691), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n689), .A2(KEYINPUT85), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n689), .A2(KEYINPUT85), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n700), .A2(KEYINPUT20), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n679), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n699), .A2(new_n702), .A3(new_n679), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n678), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n707), .A2(new_n677), .A3(new_n703), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n676), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n677), .B1(new_n707), .B2(new_n703), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(new_n678), .A3(new_n705), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(new_n711), .A3(new_n675), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n709), .A2(new_n712), .ZN(G229));
  OR2_X1    g288(.A1(G6), .A2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(G305), .B2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n715), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n715), .ZN(new_n721));
  INV_X1    g296(.A(G1971), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n715), .A2(G23), .ZN(new_n724));
  INV_X1    g299(.A(G288), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n715), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT33), .B(G1976), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n718), .A2(new_n719), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT93), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT92), .B(KEYINPUT34), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(new_n732), .ZN(new_n734));
  MUX2_X1   g309(.A(G24), .B(G290), .S(G16), .Z(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT91), .B(G1986), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT94), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT87), .B(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT88), .ZN(new_n741));
  OAI21_X1  g316(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NOR3_X1   g318(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n744));
  OAI221_X1 g319(.A(G2104), .B1(G107), .B2(new_n483), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G119), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n481), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G131), .B2(new_n488), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n741), .B1(new_n748), .B2(new_n739), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT90), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT35), .B(G1991), .Z(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n750), .B(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n738), .B(new_n753), .C1(new_n735), .C2(new_n737), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n733), .A2(new_n734), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n733), .A2(KEYINPUT36), .A3(new_n734), .A4(new_n754), .ZN(new_n758));
  NOR2_X1   g333(.A1(G171), .A2(new_n715), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G5), .B2(new_n715), .ZN(new_n760));
  INV_X1    g335(.A(G1961), .ZN(new_n761));
  NOR2_X1   g336(.A1(G16), .A2(G19), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n546), .B2(G16), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n760), .A2(new_n761), .B1(new_n763), .B2(G1341), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n761), .B2(new_n760), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n620), .A2(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G4), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2078), .ZN(new_n770));
  NOR2_X1   g345(.A1(G164), .A2(new_n739), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G27), .B2(new_n739), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G11), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(KEYINPUT31), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(KEYINPUT31), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G28), .ZN(new_n778));
  INV_X1    g353(.A(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n777), .B2(G28), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n775), .B(new_n776), .C1(new_n778), .C2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n739), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n781), .B1(new_n635), .B2(new_n782), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n783), .B1(new_n763), .B2(G1341), .C1(new_n767), .C2(new_n768), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n772), .A2(new_n770), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n765), .A2(new_n773), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n715), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n715), .ZN(new_n788));
  INV_X1    g363(.A(G2090), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n782), .A2(G35), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G162), .B2(new_n782), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT29), .Z(new_n792));
  OAI221_X1 g367(.A(new_n786), .B1(G1966), .B2(new_n788), .C1(new_n789), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n779), .A2(G32), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT26), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n797), .A2(new_n798), .B1(G105), .B2(new_n477), .ZN(new_n799));
  INV_X1    g374(.A(G141), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n487), .B2(new_n800), .ZN(new_n801));
  AND4_X1   g376(.A1(G2105), .A2(new_n463), .A3(new_n466), .A4(new_n467), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n802), .A2(KEYINPUT100), .A3(G129), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n804));
  INV_X1    g379(.A(G129), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n481), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n801), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n794), .B1(new_n807), .B2(new_n779), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT27), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(G1996), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n739), .A2(G26), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT28), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n488), .A2(G140), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n802), .A2(G128), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n483), .A2(G116), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n813), .B(new_n814), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n812), .B1(new_n821), .B2(G29), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G2067), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n810), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(G29), .A2(G33), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT96), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n483), .A2(G103), .A3(G2104), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G139), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n487), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n829), .B(KEYINPUT97), .C1(new_n830), .C2(new_n487), .ZN(new_n834));
  NAND2_X1  g409(.A1(G115), .A2(G2104), .ZN(new_n835));
  INV_X1    g410(.A(G127), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n474), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n833), .A2(new_n834), .B1(G2105), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n826), .B1(new_n838), .B2(G29), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(G2072), .Z(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT98), .B(KEYINPUT24), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(G34), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(G34), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n739), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(new_n479), .B2(new_n779), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT99), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n840), .B1(new_n846), .B2(G2084), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n792), .A2(new_n789), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n715), .A2(G20), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT23), .Z(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G299), .B2(G16), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G1956), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n788), .A2(G1966), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(G2084), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n848), .A2(new_n852), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  NOR4_X1   g430(.A1(new_n793), .A2(new_n824), .A3(new_n847), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n757), .A2(new_n758), .A3(new_n856), .ZN(G150));
  INV_X1    g432(.A(G150), .ZN(G311));
  NAND2_X1  g433(.A1(new_n620), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n861), .A2(new_n508), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n512), .A2(G55), .ZN(new_n863));
  INV_X1    g438(.A(G93), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n515), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n545), .B(new_n866), .Z(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n860), .B(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  INV_X1    g445(.A(G860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n866), .A2(new_n871), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(G145));
  NAND2_X1  g451(.A1(new_n488), .A2(G142), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n802), .A2(G130), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n483), .A2(G118), .ZN(new_n879));
  OAI21_X1  g454(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n878), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n628), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n748), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n833), .A2(new_n834), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n837), .A2(G2105), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n807), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n807), .B1(new_n838), .B2(KEYINPUT101), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n495), .A2(new_n499), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n894), .A2(new_n895), .A3(new_n821), .ZN(new_n896));
  INV_X1    g471(.A(new_n821), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n838), .A2(KEYINPUT101), .A3(new_n807), .ZN(new_n899));
  OAI21_X1  g474(.A(G164), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n885), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n821), .B1(new_n894), .B2(new_n895), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n897), .A3(new_n901), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n904), .A2(new_n905), .A3(new_n884), .A4(new_n883), .ZN(new_n906));
  XOR2_X1   g481(.A(G162), .B(new_n635), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(G160), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n903), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n883), .B1(new_n896), .B2(new_n902), .ZN(new_n911));
  INV_X1    g486(.A(new_n883), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n912), .A2(new_n904), .A3(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n910), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(G395));
  XNOR2_X1  g493(.A(new_n867), .B(new_n623), .ZN(new_n919));
  AOI21_X1  g494(.A(KEYINPUT104), .B1(G299), .B2(new_n620), .ZN(new_n920));
  NAND2_X1  g495(.A1(G299), .A2(new_n620), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n612), .A2(new_n561), .A3(new_n571), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(new_n923), .B2(KEYINPUT104), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(KEYINPUT105), .ZN(new_n927));
  INV_X1    g502(.A(new_n919), .ZN(new_n928));
  INV_X1    g503(.A(new_n922), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n612), .B1(new_n561), .B2(new_n571), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT104), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n920), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n923), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n926), .A2(KEYINPUT105), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n927), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT42), .ZN(new_n941));
  XNOR2_X1  g516(.A(G288), .B(KEYINPUT107), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n942), .A2(G305), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(G305), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(G290), .A2(G166), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n602), .A2(G303), .A3(new_n603), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n943), .A2(new_n946), .A3(new_n947), .A4(new_n944), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n927), .A2(new_n952), .A3(new_n938), .A4(new_n939), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n941), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n941), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G868), .B2(new_n866), .ZN(G295));
  OAI21_X1  g532(.A(new_n956), .B1(G868), .B2(new_n866), .ZN(G331));
  AND3_X1   g533(.A1(new_n504), .A2(KEYINPUT5), .A3(G543), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT5), .B1(new_n504), .B2(G543), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n528), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT70), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n506), .A2(new_n526), .A3(new_n528), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n533), .B1(new_n964), .B2(new_n525), .ZN(new_n965));
  INV_X1    g540(.A(new_n534), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n523), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT76), .ZN(new_n968));
  NAND2_X1  g543(.A1(G168), .A2(new_n574), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(G171), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G301), .A2(G168), .ZN(new_n971));
  AND3_X1   g546(.A1(new_n970), .A2(new_n867), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n867), .B1(new_n970), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n937), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G171), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n575), .A2(new_n576), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n615), .A2(new_n967), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n868), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n970), .A2(new_n867), .A3(new_n971), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n925), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n980), .A3(new_n951), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(new_n915), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n921), .A2(KEYINPUT41), .A3(new_n922), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(new_n924), .B2(new_n933), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n972), .B2(new_n973), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n980), .ZN(new_n988));
  INV_X1    g563(.A(new_n951), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI211_X1 g565(.A(KEYINPUT108), .B(new_n951), .C1(new_n987), .C2(new_n980), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n982), .B(new_n983), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n981), .A2(new_n915), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n951), .B1(new_n974), .B2(new_n980), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT43), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT44), .ZN(new_n997));
  INV_X1    g572(.A(new_n994), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n982), .A2(new_n983), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT109), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n982), .A2(new_n1001), .A3(new_n983), .A4(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n988), .A2(new_n989), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT108), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n988), .A2(new_n984), .A3(new_n989), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n993), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1000), .B(new_n1002), .C1(new_n983), .C2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n997), .B1(KEYINPUT44), .B2(new_n1007), .ZN(G397));
  INV_X1    g583(.A(G2067), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n821), .B(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1996), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n807), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n495), .B2(new_n499), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n471), .A2(G40), .A3(new_n478), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1012), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1011), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n807), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n748), .B(new_n752), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1024), .B1(new_n1018), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G290), .A2(G1986), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1018), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G305), .A2(G1981), .ZN(new_n1032));
  INV_X1    g607(.A(G1981), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n589), .A2(new_n1033), .A3(new_n590), .A4(new_n595), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1032), .A2(new_n1037), .A3(new_n1034), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT114), .B(G8), .C1(new_n1017), .C2(new_n1014), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1017), .B2(new_n1014), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1036), .A2(new_n1038), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  OAI211_X1 g620(.A(G303), .B(G8), .C1(new_n1045), .C2(KEYINPUT55), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(G166), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1017), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1014), .A2(KEYINPUT50), .ZN(new_n1052));
  NOR2_X1   g627(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n495), .B2(new_n499), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n893), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(new_n1051), .A3(new_n1016), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1055), .A2(new_n789), .B1(new_n1057), .B2(new_n722), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1050), .B1(new_n1058), .B2(new_n1048), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1042), .A2(new_n1039), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G288), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1060), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1060), .B1(new_n725), .B2(G1976), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1063), .B(new_n1067), .C1(new_n1042), .C2(new_n1039), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1044), .A2(new_n1059), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1054), .B(KEYINPUT111), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1017), .B1(KEYINPUT50), .B2(new_n1014), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n789), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1057), .A2(new_n722), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1077), .A2(new_n1050), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1057), .B2(G2078), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n761), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1057), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT122), .B(new_n1080), .C1(new_n1057), .C2(G2078), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1083), .A2(new_n1085), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n615), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1070), .A2(new_n1079), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1966), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1057), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1084), .B2(G2084), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(G8), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G168), .A2(new_n1048), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1095), .B(new_n1097), .C1(KEYINPUT120), .C2(KEYINPUT51), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT51), .B1(new_n1097), .B2(KEYINPUT120), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(G8), .C1(new_n1094), .C2(new_n967), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT62), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1098), .A2(new_n1100), .A3(new_n1104), .A4(new_n1101), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1091), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1043), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n725), .A2(new_n1062), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1034), .B1(new_n1043), .B2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1079), .A2(new_n1107), .B1(new_n1109), .B2(new_n1061), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1050), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1107), .A2(new_n1111), .A3(KEYINPUT115), .ZN(new_n1112));
  OR3_X1    g687(.A1(new_n1077), .A2(new_n1050), .A3(new_n1078), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1095), .A2(G286), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(KEYINPUT63), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT115), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1112), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1070), .A2(new_n1079), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT63), .B1(new_n1118), .B2(new_n1114), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1106), .B(new_n1110), .C1(new_n1117), .C2(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1083), .A2(new_n1088), .A3(new_n1085), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1121), .A2(new_n1122), .A3(G301), .A4(new_n1087), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT124), .B1(new_n1089), .B2(new_n615), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1081), .A2(new_n1082), .B1(new_n761), .B2(new_n1084), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1056), .A2(new_n1016), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1086), .B1(new_n1051), .B2(KEYINPUT123), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1126), .B(new_n1127), .C1(KEYINPUT123), .C2(new_n1051), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1088), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1123), .A2(KEYINPUT54), .A3(new_n1124), .A4(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1125), .A2(G301), .A3(new_n1088), .A4(new_n1128), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1090), .A2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(new_n1118), .A3(new_n1135), .A4(new_n1102), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1055), .A2(G1956), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1056), .A2(new_n1051), .A3(new_n1016), .A4(new_n1138), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n1139), .A2(KEYINPUT116), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(KEYINPUT116), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1137), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(G299), .B(KEYINPUT57), .Z(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1137), .A2(new_n1140), .A3(new_n1143), .A4(new_n1141), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1148), .B(new_n1149), .C1(new_n1146), .C2(new_n1145), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n546), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1126), .A2(new_n1011), .A3(new_n1051), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1017), .A2(new_n1014), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT58), .B(G1341), .Z(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1149), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1147), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1155), .A2(G2067), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1163), .B1(new_n1084), .B2(new_n768), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(KEYINPUT119), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(KEYINPUT119), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n620), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(KEYINPUT119), .A3(new_n612), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1150), .B(new_n1162), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1164), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1147), .A2(new_n620), .A3(new_n1173), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1174), .A2(new_n1145), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1136), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1031), .B1(new_n1120), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1029), .A2(new_n1018), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT48), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n897), .A2(new_n1009), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n748), .A2(new_n751), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1024), .B2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1027), .A2(new_n1179), .B1(new_n1182), .B2(new_n1018), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1010), .A2(new_n807), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  XNOR2_X1  g760(.A(new_n1020), .B(KEYINPUT110), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1184), .A2(new_n1018), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1022), .A2(KEYINPUT125), .A3(KEYINPUT46), .ZN(new_n1188));
  AOI21_X1  g763(.A(KEYINPUT125), .B1(new_n1022), .B2(KEYINPUT46), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1187), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT47), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1183), .B1(new_n1192), .B2(KEYINPUT126), .ZN(new_n1193));
  XNOR2_X1  g768(.A(new_n1190), .B(KEYINPUT47), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1177), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g773(.A1(new_n672), .A2(new_n655), .A3(G319), .A4(new_n673), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n709), .B2(new_n712), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n916), .A2(new_n1201), .ZN(new_n1202));
  AOI211_X1 g776(.A(KEYINPUT127), .B(new_n1202), .C1(new_n992), .C2(new_n995), .ZN(new_n1203));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n1204));
  INV_X1    g778(.A(new_n1202), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1204), .B1(new_n996), .B2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g780(.A1(new_n1203), .A2(new_n1206), .ZN(G308));
  NAND2_X1  g781(.A1(new_n996), .A2(new_n1205), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1208), .A2(KEYINPUT127), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n996), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1210), .ZN(G225));
endmodule


