//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G250), .B1(G257), .B2(G264), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(new_n212), .B2(new_n213), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G77), .ZN(new_n227));
  INV_X1    g0027(.A(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G107), .ZN(new_n229));
  INV_X1    g0029(.A(G264), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n226), .B1(new_n227), .B2(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n208), .B1(new_n225), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n219), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n244), .B(new_n245), .Z(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  NAND2_X1  g0050(.A1(KEYINPUT66), .A2(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT8), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(new_n206), .A3(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n253), .B(new_n254), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n214), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n260), .B1(new_n205), .B2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G20), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n261), .B(new_n263), .C1(G50), .C2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G41), .ZN(new_n270));
  OAI211_X1 g0070(.A(G1), .B(G13), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n271), .A2(G274), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n275), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  XOR2_X1   g0077(.A(KEYINPUT65), .B(G1698), .Z(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(G222), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G1698), .ZN(new_n282));
  OAI221_X1 g0082(.A(new_n280), .B1(new_n227), .B2(new_n279), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  AOI211_X1 g0083(.A(new_n274), .B(new_n277), .C1(new_n283), .C2(new_n275), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G190), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n268), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G200), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n288), .B1(KEYINPUT69), .B2(KEYINPUT10), .ZN(new_n289));
  NAND2_X1  g0089(.A1(KEYINPUT69), .A2(KEYINPUT10), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n284), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n267), .B1(new_n284), .B2(G169), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n266), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n252), .ZN(new_n297));
  INV_X1    g0097(.A(new_n262), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n252), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G58), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(new_n221), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(new_n201), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(G20), .B1(G159), .B2(new_n256), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT3), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n307));
  AOI21_X1  g0107(.A(G20), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n308), .A2(KEYINPUT7), .B1(new_n309), .B2(new_n279), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n310), .A2(new_n311), .A3(G68), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n310), .B2(G68), .ZN(new_n313));
  OAI211_X1 g0113(.A(KEYINPUT16), .B(new_n304), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n260), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT73), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n305), .A2(KEYINPUT73), .A3(G33), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(new_n307), .ZN(new_n319));
  INV_X1    g0119(.A(new_n309), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(KEYINPUT74), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n279), .B2(G20), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT74), .B1(new_n319), .B2(new_n320), .ZN(new_n325));
  OAI21_X1  g0125(.A(G68), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT16), .B1(new_n326), .B2(new_n304), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n300), .B1(new_n315), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n274), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n275), .A2(new_n273), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G232), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n306), .A2(new_n307), .A3(G226), .A4(G1698), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G87), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT65), .A2(G1698), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n335), .A2(new_n306), .A3(new_n307), .A4(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n333), .B(new_n334), .C1(new_n337), .C2(new_n281), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT75), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n271), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n278), .A2(G223), .A3(new_n279), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n333), .A4(new_n334), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n332), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G179), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n343), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n328), .A2(KEYINPUT18), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT76), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT76), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n328), .A2(new_n349), .A3(KEYINPUT18), .A4(new_n346), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT18), .ZN(new_n351));
  INV_X1    g0151(.A(new_n260), .ZN(new_n352));
  INV_X1    g0152(.A(new_n304), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n309), .B1(new_n306), .B2(new_n307), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n305), .A2(G33), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n206), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n354), .B1(new_n357), .B2(new_n322), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT72), .B1(new_n358), .B2(new_n221), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n310), .A2(new_n311), .A3(G68), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n353), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n352), .B1(new_n361), .B2(KEYINPUT16), .ZN(new_n362));
  INV_X1    g0162(.A(new_n327), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n299), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n343), .A2(new_n345), .ZN(new_n365));
  AOI211_X1 g0165(.A(new_n292), .B(new_n332), .C1(new_n340), .C2(new_n342), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n351), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n348), .A2(new_n350), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  AOI211_X1 g0170(.A(new_n370), .B(new_n332), .C1(new_n340), .C2(new_n342), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n338), .A2(new_n339), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(new_n342), .A3(new_n275), .ZN(new_n373));
  INV_X1    g0173(.A(new_n332), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n287), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n325), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n377), .A2(new_n323), .A3(new_n321), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n353), .B1(new_n378), .B2(G68), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n314), .B(new_n260), .C1(new_n379), .C2(KEYINPUT16), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n376), .A2(new_n380), .A3(KEYINPUT77), .A4(new_n300), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n364), .A2(KEYINPUT77), .A3(KEYINPUT17), .A4(new_n376), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n369), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT12), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n266), .B2(G68), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n296), .A2(KEYINPUT12), .A3(new_n221), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n388), .B(new_n389), .C1(new_n298), .C2(new_n221), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT71), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n391), .ZN(new_n393));
  INV_X1    g0193(.A(G50), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n257), .A2(new_n394), .B1(new_n206), .B2(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n206), .A2(G33), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n396), .A2(new_n227), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n260), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT11), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(new_n393), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT14), .ZN(new_n401));
  NAND2_X1  g0201(.A1(G33), .A2(G97), .ZN(new_n402));
  OAI221_X1 g0202(.A(new_n402), .B1(new_n337), .B2(new_n276), .C1(new_n236), .C2(new_n282), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n275), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n274), .B1(G238), .B2(new_n330), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n406), .A2(new_n408), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n401), .B(G169), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n404), .A2(new_n405), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n407), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(G179), .C1(new_n415), .C2(new_n413), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n409), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n401), .B1(new_n418), .B2(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n400), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(G200), .ZN(new_n421));
  INV_X1    g0221(.A(new_n400), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n414), .B(G190), .C1(new_n415), .C2(new_n413), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(KEYINPUT15), .B(G87), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n426), .A2(new_n396), .B1(new_n206), .B2(new_n227), .ZN(new_n427));
  XNOR2_X1  g0227(.A(KEYINPUT8), .B(G58), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT67), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n427), .B1(new_n429), .B2(new_n256), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n352), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n296), .A2(new_n227), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n298), .B2(new_n227), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT68), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n274), .B1(G244), .B2(new_n330), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n337), .A2(new_n236), .B1(new_n229), .B2(new_n279), .ZN(new_n437));
  INV_X1    g0237(.A(new_n282), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n437), .B1(G238), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n436), .B1(new_n439), .B2(new_n271), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(G200), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n370), .B2(new_n440), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n435), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n440), .A2(G179), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n345), .B2(new_n440), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n435), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NOR4_X1   g0247(.A1(new_n295), .A2(new_n386), .A3(new_n425), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n306), .A2(new_n307), .A3(G244), .A4(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G116), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(new_n450), .C1(new_n337), .C2(new_n222), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n278), .A2(G238), .A3(new_n279), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n449), .A4(new_n450), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n271), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n272), .A2(G1), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n271), .A2(new_n458), .A3(G250), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n271), .A2(G274), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n458), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n292), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n345), .B1(new_n456), .B2(new_n461), .ZN(new_n464));
  INV_X1    g0264(.A(G97), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n223), .A2(new_n465), .A3(new_n229), .ZN(new_n466));
  XNOR2_X1  g0266(.A(new_n466), .B(KEYINPUT80), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n402), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G20), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n279), .A2(new_n206), .A3(G68), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n468), .B1(new_n396), .B2(new_n465), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n260), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n296), .A2(new_n426), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n205), .A2(G33), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n352), .A2(new_n266), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n475), .B(new_n476), .C1(new_n426), .C2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n463), .A2(new_n464), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(G200), .B1(new_n456), .B2(new_n461), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n352), .A2(new_n266), .A3(new_n477), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G87), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n475), .A2(new_n476), .A3(new_n483), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n456), .A2(new_n461), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n481), .B(new_n484), .C1(new_n485), .C2(new_n370), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n206), .A2(G107), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT23), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n206), .B2(G107), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n279), .A2(new_n206), .A3(G87), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT22), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT22), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n279), .A2(new_n496), .A3(new_n206), .A4(G87), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(KEYINPUT24), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n260), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n265), .A2(new_n487), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n503));
  OR2_X1    g0303(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT84), .A2(KEYINPUT25), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n265), .A2(new_n487), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n503), .B(new_n506), .C1(new_n478), .C2(new_n229), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n507), .B(KEYINPUT85), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n279), .A2(G257), .A3(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(G294), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n512));
  OAI21_X1  g0312(.A(G33), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n509), .B(new_n513), .C1(new_n224), .C2(new_n337), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n275), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT5), .B(G41), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n457), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n517), .A2(new_n460), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n275), .B1(new_n457), .B2(new_n516), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G264), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n515), .A2(G190), .A3(new_n521), .A4(new_n519), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n501), .A2(new_n508), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n480), .A2(new_n486), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n520), .A2(G257), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n519), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G283), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(KEYINPUT4), .B1(new_n337), .B2(new_n228), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n278), .A2(new_n534), .A3(G244), .A4(new_n279), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT78), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n275), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI211_X1 g0338(.A(KEYINPUT78), .B(new_n532), .C1(new_n533), .C2(new_n535), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n529), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n345), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n266), .A2(G97), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(new_n482), .B2(G97), .ZN(new_n543));
  XNOR2_X1  g0343(.A(G97), .B(G107), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n545), .A2(new_n465), .A3(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n548), .A2(new_n206), .B1(new_n227), .B2(new_n257), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(new_n378), .B2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n543), .B1(new_n550), .B2(new_n352), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n292), .B(new_n529), .C1(new_n538), .C2(new_n539), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n541), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n540), .A2(new_n287), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n370), .B(new_n529), .C1(new_n538), .C2(new_n539), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g0356(.A1(new_n526), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT83), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n531), .B(new_n206), .C1(G33), .C2(new_n465), .ZN(new_n559));
  INV_X1    g0359(.A(G116), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n260), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n266), .A2(G116), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n482), .B2(G116), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n517), .A2(G270), .A3(new_n271), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT81), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n520), .A2(KEYINPUT81), .A3(G270), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n279), .A2(G257), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n335), .A2(new_n336), .ZN(new_n575));
  INV_X1    g0375(.A(G303), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n279), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n282), .A2(new_n230), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n275), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n573), .A2(new_n579), .A3(new_n519), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n558), .B(new_n568), .C1(new_n580), .C2(new_n287), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n518), .B1(new_n571), .B2(new_n572), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n287), .B1(new_n582), .B2(new_n579), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT83), .B1(new_n583), .B2(new_n567), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n580), .A2(G190), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n573), .A2(new_n579), .A3(new_n519), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n345), .B1(new_n564), .B2(new_n566), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT82), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n567), .A2(new_n582), .A3(G179), .A4(new_n579), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n590), .B1(new_n587), .B2(new_n588), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n500), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n260), .B1(new_n498), .B2(KEYINPUT24), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n508), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n522), .A2(new_n345), .ZN(new_n599));
  OR2_X1    g0399(.A1(new_n522), .A2(G179), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n586), .A2(new_n595), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n448), .A2(new_n557), .A3(new_n602), .ZN(G372));
  NOR2_X1   g0403(.A1(new_n293), .A2(new_n294), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n368), .A2(new_n347), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n420), .ZN(new_n607));
  INV_X1    g0407(.A(new_n446), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n424), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n383), .A2(new_n384), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n604), .B1(new_n611), .B2(new_n291), .ZN(new_n612));
  INV_X1    g0412(.A(new_n448), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n486), .A2(new_n480), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT26), .B1(new_n614), .B2(new_n553), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n486), .A2(new_n480), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n541), .A2(new_n551), .A3(new_n552), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n480), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n553), .A2(new_n556), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n480), .A2(new_n486), .A3(new_n525), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(KEYINPUT87), .A3(new_n622), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n593), .A2(new_n594), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT88), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n598), .A2(new_n626), .A3(new_n599), .A4(new_n600), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n554), .A2(new_n555), .ZN(new_n629));
  INV_X1    g0429(.A(new_n551), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n622), .A2(new_n617), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT87), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n628), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n620), .B1(new_n623), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n612), .B1(new_n613), .B2(new_n635), .ZN(G369));
  NAND2_X1  g0436(.A1(new_n265), .A2(new_n206), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT89), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n567), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n586), .A2(new_n595), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n595), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n598), .A2(new_n643), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n601), .A2(new_n525), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n643), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n601), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n595), .A2(new_n643), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n625), .A2(new_n627), .ZN(new_n656));
  OAI22_X1  g0456(.A1(new_n655), .A2(new_n650), .B1(new_n656), .B2(new_n643), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(G399));
  NOR2_X1   g0459(.A1(new_n210), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n467), .A2(new_n560), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(G1), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n216), .B2(new_n661), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n665), .B(KEYINPUT28), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT31), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n587), .A2(new_n292), .A3(new_n522), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n540), .A3(new_n485), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n540), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n587), .A2(new_n292), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT90), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n515), .A2(new_n521), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n462), .B2(new_n675), .ZN(new_n676));
  NOR4_X1   g0476(.A1(new_n456), .A2(new_n674), .A3(KEYINPUT90), .A4(new_n461), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n671), .B(new_n672), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT30), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n670), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n540), .A2(new_n292), .A3(new_n587), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n681), .B(KEYINPUT30), .C1(new_n677), .C2(new_n676), .ZN(new_n682));
  AOI211_X1 g0482(.A(new_n667), .B(new_n651), .C1(new_n680), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n679), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n684), .A2(new_n682), .A3(new_n669), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT31), .B1(new_n685), .B2(new_n643), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n621), .A2(new_n602), .A3(new_n622), .A4(new_n651), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n557), .A2(KEYINPUT91), .A3(new_n602), .A4(new_n651), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G330), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT92), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n635), .B2(new_n643), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT93), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n631), .A2(new_n617), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n633), .B1(new_n700), .B2(new_n526), .ZN(new_n701));
  INV_X1    g0501(.A(new_n628), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n623), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n480), .ZN(new_n704));
  INV_X1    g0504(.A(new_n619), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n618), .B1(new_n616), .B2(new_n617), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(KEYINPUT92), .A3(new_n651), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n698), .A2(new_n699), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n601), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n557), .B1(new_n624), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n643), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n698), .A2(new_n710), .A3(new_n709), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT93), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n696), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n666), .B1(new_n719), .B2(G1), .ZN(G364));
  NOR2_X1   g0520(.A1(new_n264), .A2(G20), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n205), .B1(new_n721), .B2(G45), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n660), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n648), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G330), .B2(new_n646), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n209), .A2(new_n279), .ZN(new_n727));
  INV_X1    g0527(.A(G355), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n727), .A2(new_n728), .B1(G116), .B2(new_n209), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n210), .A2(new_n279), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n731), .B1(new_n272), .B2(new_n217), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n246), .A2(new_n272), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G13), .A2(G33), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G20), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n214), .B1(G20), .B2(new_n345), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n724), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  AND3_X1   g0541(.A1(KEYINPUT94), .A2(G20), .A3(G179), .ZN(new_n742));
  AOI21_X1  g0542(.A(KEYINPUT94), .B1(G20), .B2(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n370), .A2(new_n287), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n287), .A2(G190), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(KEYINPUT33), .B(G317), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G326), .A2(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n206), .A2(G179), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n749), .ZN(new_n755));
  INV_X1    g0555(.A(G283), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n306), .A2(new_n307), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n746), .A2(new_n754), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n759), .B2(new_n576), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G190), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g0563(.A(new_n757), .B(new_n760), .C1(G329), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n511), .A2(new_n512), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n292), .A2(new_n287), .A3(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n745), .A2(new_n761), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR3_X1   g0571(.A1(new_n744), .A2(new_n370), .A3(G200), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n771), .A2(G311), .B1(G322), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n753), .A2(new_n764), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n227), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n763), .A2(KEYINPUT32), .A3(G159), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT32), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n781), .B1(new_n762), .B2(new_n782), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n751), .A2(G68), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n748), .A2(G50), .B1(G58), .B2(new_n772), .ZN(new_n785));
  INV_X1    g0585(.A(new_n768), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n465), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n759), .A2(new_n223), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n755), .A2(new_n229), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n758), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n784), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n774), .B1(new_n779), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n741), .B1(new_n792), .B2(new_n738), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n737), .B(KEYINPUT96), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n646), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n726), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NAND2_X1  g0597(.A1(new_n435), .A2(new_n643), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n443), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n446), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n608), .A2(new_n651), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n698), .A2(new_n709), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n802), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n708), .A2(new_n804), .A3(new_n651), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n696), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n724), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n696), .A2(new_n803), .A3(new_n805), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n738), .A2(new_n735), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n724), .B1(G77), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n772), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n813), .A2(new_n510), .B1(new_n576), .B2(new_n747), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G283), .B2(new_n751), .ZN(new_n815));
  INV_X1    g0615(.A(G311), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n759), .A2(new_n229), .B1(new_n762), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n758), .B1(new_n755), .B2(new_n223), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n787), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n815), .B(new_n819), .C1(new_n560), .C2(new_n778), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n751), .A2(G150), .B1(G143), .B2(new_n772), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n747), .C1(new_n778), .C2(new_n782), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT97), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n279), .B1(new_n755), .B2(new_n221), .ZN(new_n826));
  INV_X1    g0626(.A(G132), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n759), .A2(new_n394), .B1(new_n762), .B2(new_n827), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(G58), .C2(new_n768), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n824), .A2(KEYINPUT34), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n820), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n812), .B1(new_n832), .B2(new_n738), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT98), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n835), .B(new_n836), .C1(new_n735), .C2(new_n802), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n809), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G384));
  INV_X1    g0639(.A(new_n548), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n840), .A2(KEYINPUT35), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(KEYINPUT35), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n841), .A2(G116), .A3(new_n215), .A4(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT36), .Z(new_n844));
  OR3_X1    g0644(.A1(new_n216), .A2(new_n227), .A3(new_n302), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n394), .A2(G68), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n205), .B(G13), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT101), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n364), .A2(new_n376), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n361), .A2(KEYINPUT16), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n300), .B1(new_n315), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n641), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n852), .A2(new_n346), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n850), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n856), .A2(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n328), .A2(new_n346), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n328), .A2(new_n853), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n850), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT99), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n368), .A2(new_n350), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n610), .B1(new_n864), .B2(new_n348), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n863), .B1(new_n865), .B2(new_n854), .ZN(new_n866));
  INV_X1    g0666(.A(new_n854), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n386), .A2(KEYINPUT99), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n862), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n849), .B1(new_n869), .B2(KEYINPUT38), .ZN(new_n870));
  INV_X1    g0670(.A(new_n862), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n865), .A2(new_n863), .A3(new_n854), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT99), .B1(new_n386), .B2(new_n867), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(KEYINPUT101), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT100), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n866), .A2(new_n868), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT38), .B1(new_n857), .B2(new_n861), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g0681(.A(KEYINPUT100), .B(new_n879), .C1(new_n866), .C2(new_n868), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n870), .B(new_n876), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n805), .A2(new_n801), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n651), .A2(new_n422), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n425), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n425), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n883), .A2(new_n891), .B1(new_n605), .B2(new_n641), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n878), .A2(new_n880), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT103), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n605), .B1(new_n894), .B2(new_n610), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n385), .A2(KEYINPUT103), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n859), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n860), .A2(KEYINPUT102), .A3(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n875), .B1(new_n897), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n893), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n883), .B2(KEYINPUT39), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n607), .A2(new_n651), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n892), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n718), .A2(new_n448), .A3(new_n715), .A4(new_n711), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(new_n612), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n909), .B(new_n911), .ZN(new_n912));
  NOR4_X1   g0712(.A1(new_n694), .A2(new_n890), .A3(KEYINPUT40), .A4(new_n802), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n883), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n893), .A2(new_n904), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n693), .A2(new_n804), .A3(new_n889), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT40), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n448), .A3(new_n693), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n883), .A2(new_n913), .B1(new_n917), .B2(KEYINPUT40), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n613), .B2(new_n694), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n920), .A2(G330), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n912), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n205), .B2(new_n721), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n912), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n848), .B1(new_n925), .B2(new_n926), .ZN(G367));
  OAI221_X1 g0727(.A(new_n739), .B1(new_n209), .B2(new_n426), .C1(new_n731), .C2(new_n242), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n724), .ZN(new_n929));
  INV_X1    g0729(.A(G143), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n813), .A2(new_n255), .B1(new_n930), .B2(new_n747), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G159), .B2(new_n751), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n786), .A2(new_n221), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n759), .A2(new_n301), .B1(new_n762), .B2(new_n822), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n279), .B1(new_n755), .B2(new_n227), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n932), .B(new_n936), .C1(new_n394), .C2(new_n778), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n778), .A2(new_n756), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n759), .A2(new_n560), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n939), .A2(KEYINPUT46), .B1(new_n786), .B2(new_n229), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(KEYINPUT46), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(G317), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n758), .B1(new_n762), .B2(new_n942), .C1(new_n465), .C2(new_n755), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G311), .B2(new_n748), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n751), .A2(new_n766), .B1(G303), .B2(new_n772), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n941), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n937), .B1(new_n938), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT47), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n929), .B1(new_n948), .B2(new_n738), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n651), .A2(new_n484), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n614), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n480), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n949), .B1(new_n794), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT105), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n630), .A2(new_n651), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(new_n552), .A3(new_n541), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n954), .B(new_n956), .C1(new_n700), .C2(new_n955), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n956), .A2(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n655), .A2(new_n650), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n617), .B1(new_n959), .B2(new_n601), .ZN(new_n963));
  AOI22_X1  g0763(.A1(KEYINPUT42), .A2(new_n962), .B1(new_n963), .B2(new_n651), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT106), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n962), .A2(KEYINPUT42), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n964), .A2(new_n965), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT107), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n970), .A2(KEYINPUT107), .A3(new_n971), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n952), .B(KEYINPUT43), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n972), .A2(new_n973), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n653), .A2(new_n959), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n975), .B(new_n976), .Z(new_n977));
  INV_X1    g0777(.A(new_n961), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n652), .B2(new_n654), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(new_n648), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n719), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n960), .A2(new_n658), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT44), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n959), .A2(new_n657), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT45), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n653), .A2(KEYINPUT108), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n982), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n719), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n660), .B(KEYINPUT41), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n723), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n953), .B1(new_n977), .B2(new_n994), .ZN(G387));
  NOR2_X1   g0795(.A1(new_n982), .A2(new_n661), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n719), .B2(new_n980), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n652), .A2(new_n794), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n429), .A2(new_n394), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT109), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n999), .A2(KEYINPUT50), .B1(new_n662), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(KEYINPUT50), .B2(new_n999), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n272), .B1(new_n221), .B2(new_n227), .C1(new_n662), .C2(new_n1000), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n730), .B1(new_n272), .B2(new_n239), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(G107), .B2(new_n209), .C1(new_n663), .C2(new_n727), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n739), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n724), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n759), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(G77), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n255), .B2(new_n762), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n755), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n758), .B(new_n1010), .C1(G97), .C2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n786), .A2(new_n426), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n748), .A2(G159), .B1(G50), .B2(new_n772), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G68), .A2(new_n771), .B1(new_n751), .B2(new_n252), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n763), .A2(G326), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n279), .B1(new_n1011), .B2(G116), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n813), .A2(new_n942), .B1(new_n816), .B2(new_n750), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G322), .B2(new_n748), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n576), .B2(new_n778), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT48), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n766), .A2(new_n1008), .B1(new_n768), .B2(G283), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1018), .B(new_n1019), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1017), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n998), .B(new_n1007), .C1(new_n1031), .C2(new_n738), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n980), .B2(new_n723), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n997), .A2(new_n1033), .ZN(G393));
  XOR2_X1   g0834(.A(new_n987), .B(new_n653), .Z(new_n1035));
  OAI211_X1 g0835(.A(new_n990), .B(new_n660), .C1(new_n982), .C2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n730), .A2(new_n249), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n739), .C1(new_n465), .C2(new_n209), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n724), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT110), .Z(new_n1040));
  AOI22_X1  g0840(.A1(new_n751), .A2(G303), .B1(G116), .B2(new_n768), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n510), .B2(new_n770), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT111), .Z(new_n1043));
  OAI22_X1  g0843(.A1(new_n813), .A2(new_n816), .B1(new_n942), .B2(new_n747), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n789), .A2(new_n279), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G283), .A2(new_n1008), .B1(new_n763), .B2(G322), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT112), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n748), .A2(G150), .B1(G159), .B2(new_n772), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT51), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n786), .A2(new_n227), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G68), .A2(new_n1008), .B1(new_n763), .B2(G143), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n279), .C1(new_n223), .C2(new_n755), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(G50), .C2(new_n751), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1051), .B(new_n1056), .C1(new_n429), .C2(new_n777), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1049), .A2(new_n1057), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1058), .A2(KEYINPUT113), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n738), .B1(new_n1058), .B2(KEYINPUT113), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1040), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n737), .B2(new_n959), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n1035), .B2(new_n723), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1036), .A2(new_n1063), .ZN(G390));
  AOI22_X1  g0864(.A1(new_n714), .A2(new_n800), .B1(new_n608), .B2(new_n651), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n908), .B1(new_n1065), .B2(new_n890), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n893), .B2(new_n904), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n908), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n884), .B2(new_n889), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n907), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT114), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n695), .B(new_n802), .C1(new_n687), .C2(new_n692), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n889), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n693), .A2(G330), .A3(new_n889), .A4(new_n804), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT115), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT115), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n906), .B(new_n1069), .C1(new_n883), .C2(KEYINPUT39), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1081), .B(new_n1077), .C1(new_n1082), .C2(new_n1067), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n693), .A2(G330), .A3(new_n804), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n890), .ZN(new_n1086));
  AND3_X1   g0886(.A1(new_n1086), .A2(new_n1065), .A3(new_n1075), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1086), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n884), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n696), .A2(new_n448), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n910), .A2(new_n612), .A3(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1084), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .A4(new_n1092), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n660), .A3(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1079), .A2(new_n723), .A3(new_n1083), .A4(new_n1080), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n724), .B1(new_n252), .B2(new_n811), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n777), .A2(G97), .B1(G107), .B2(new_n751), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT117), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1052), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1101), .B1(new_n221), .B2(new_n755), .C1(new_n510), .C2(new_n762), .ZN(new_n1102));
  OR3_X1    g0902(.A1(new_n788), .A2(KEYINPUT118), .A3(new_n279), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT118), .B1(new_n788), .B2(new_n279), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n756), .C2(new_n747), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1102), .B(new_n1105), .C1(G116), .C2(new_n772), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(G128), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n813), .A2(new_n827), .B1(new_n1108), .B2(new_n747), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G137), .B2(new_n751), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1008), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT53), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n759), .B2(new_n255), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n1111), .A2(new_n1113), .B1(G159), .B2(new_n768), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n777), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(G125), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n279), .B1(new_n762), .B2(new_n1118), .C1(new_n394), .C2(new_n755), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT116), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1110), .A2(new_n1114), .A3(new_n1117), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1107), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1098), .B1(new_n1122), .B2(new_n738), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n907), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n736), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1097), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1096), .A2(new_n1127), .ZN(G378));
  OAI21_X1  g0928(.A(new_n724), .B1(G50), .B2(new_n811), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT121), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n853), .A2(new_n267), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n295), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n295), .A2(new_n1132), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1135), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1139), .A2(new_n736), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n933), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1011), .A2(G58), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n758), .A2(new_n270), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G283), .B2(new_n763), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1141), .A2(new_n1009), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n813), .A2(new_n229), .B1(new_n426), .B2(new_n770), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n465), .A2(new_n750), .B1(new_n747), .B2(new_n560), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1145), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(G50), .B1(new_n269), .B2(new_n270), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1148), .A2(KEYINPUT58), .B1(new_n1143), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n772), .A2(G128), .B1(new_n1008), .B2(new_n1116), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT119), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n750), .A2(new_n827), .B1(new_n255), .B2(new_n786), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n1118), .A2(new_n747), .B1(new_n770), .B2(new_n822), .ZN(new_n1154));
  NOR3_X1   g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT59), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT120), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n269), .B(new_n270), .C1(new_n755), .C2(new_n782), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G124), .B2(new_n763), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1156), .A2(KEYINPUT120), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1150), .B1(KEYINPUT58), .B2(new_n1148), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1130), .B(new_n1140), .C1(new_n738), .C2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n919), .A2(new_n1139), .A3(G330), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1138), .B1(new_n921), .B2(new_n695), .ZN(new_n1165));
  AND4_X1   g0965(.A1(KEYINPUT122), .A2(new_n1164), .A3(new_n1165), .A4(new_n909), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1164), .A2(new_n1165), .B1(new_n909), .B2(KEYINPUT122), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1163), .B1(new_n1168), .B2(new_n723), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1091), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1095), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1139), .B1(new_n919), .B2(G330), .ZN(new_n1173));
  NOR3_X1   g0973(.A1(new_n921), .A2(new_n1138), .A3(new_n695), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n909), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1124), .A2(new_n1068), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1164), .A2(new_n1176), .A3(new_n1165), .A4(new_n892), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1172), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1171), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n660), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT57), .B1(new_n1171), .B2(new_n1168), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1169), .B1(new_n1180), .B2(new_n1181), .ZN(G375));
  NAND2_X1  g0982(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1093), .A2(new_n993), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n890), .A2(new_n735), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n724), .B1(G68), .B2(new_n811), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G132), .A2(new_n748), .B1(new_n751), .B2(new_n1116), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n822), .B2(new_n813), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT125), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n786), .A2(new_n394), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G159), .A2(new_n1008), .B1(new_n763), .B2(G128), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n279), .A3(new_n1142), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G150), .C2(new_n771), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1189), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1188), .A2(KEYINPUT125), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT124), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n747), .A2(new_n510), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT123), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n759), .A2(new_n465), .B1(new_n762), .B2(new_n576), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n813), .A2(new_n756), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1198), .B(new_n1201), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n758), .B1(new_n755), .B2(new_n227), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1203), .B(new_n1013), .C1(new_n751), .C2(G116), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1204), .C1(new_n229), .C2(new_n778), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1196), .B1(new_n1197), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1197), .B2(new_n1205), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1186), .B1(new_n1207), .B2(new_n738), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1185), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1089), .B2(new_n722), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1184), .A2(new_n1211), .ZN(G381));
  OR4_X1    g1012(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1213), .A2(G387), .A3(G381), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n661), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1126), .B1(new_n1215), .B2(new_n1095), .ZN(new_n1216));
  INV_X1    g1016(.A(G375), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1214), .A2(new_n1216), .A3(new_n1217), .ZN(G407));
  NAND2_X1  g1018(.A1(new_n642), .A2(G213), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1216), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(G407), .A2(new_n1221), .A3(G213), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT126), .ZN(G409));
  NAND2_X1  g1023(.A1(new_n1088), .A2(new_n884), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1087), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1091), .A2(new_n1224), .A3(KEYINPUT60), .A4(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1226), .A2(new_n660), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT60), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1183), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G384), .B1(new_n1230), .B2(new_n1211), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n838), .B(new_n1210), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT127), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1220), .A2(G2897), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1234), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1236), .B1(new_n1237), .B2(KEYINPUT127), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1233), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1235), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1169), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1171), .A2(new_n1168), .A3(new_n993), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n722), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(new_n1163), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1216), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1219), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1241), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT63), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1237), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G387), .A2(new_n1036), .A3(new_n1063), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(G393), .B(new_n796), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n953), .B(G390), .C1(new_n977), .C2(new_n994), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1220), .B1(new_n1242), .B2(new_n1246), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(KEYINPUT63), .A3(new_n1237), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1249), .A2(new_n1252), .A3(new_n1258), .A4(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT62), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1259), .A2(new_n1262), .A3(new_n1237), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1259), .B2(new_n1240), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1262), .B1(new_n1259), .B2(new_n1237), .ZN(new_n1266));
  NOR3_X1   g1066(.A1(new_n1263), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1267), .B2(new_n1258), .ZN(G405));
  AND2_X1   g1068(.A1(G375), .A2(new_n1216), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1242), .ZN(new_n1270));
  OR3_X1    g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1237), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1237), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1258), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1271), .A2(new_n1258), .A3(new_n1272), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(G402));
endmodule


