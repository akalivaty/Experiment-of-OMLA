//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  XNOR2_X1  g000(.A(G116), .B(G119), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT64), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G137), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n193), .A2(new_n195), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n197), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n192), .A2(G137), .ZN(new_n200));
  OAI21_X1  g014(.A(G131), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  AND4_X1   g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .A4(G128), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n205), .B(G146), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n203), .A3(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n198), .B(new_n201), .C1(new_n207), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n193), .A2(new_n197), .A3(new_n195), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n206), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G143), .B(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n217), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n215), .A2(new_n198), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n190), .B1(new_n213), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n189), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n188), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n215), .A2(new_n198), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n222), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n229), .A3(new_n212), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT28), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n233), .B(G101), .ZN(new_n234));
  INV_X1    g048(.A(G237), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G237), .ZN(new_n238));
  AOI21_X1  g052(.A(G953), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G210), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n234), .B(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n230), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n232), .A2(KEYINPUT29), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G902), .ZN(new_n245));
  AND2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XOR2_X1   g060(.A(new_n246), .B(KEYINPUT69), .Z(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n242), .B1(new_n224), .B2(new_n230), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n230), .A2(new_n242), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n241), .ZN(new_n254));
  INV_X1    g068(.A(new_n230), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT30), .B1(new_n213), .B2(new_n223), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n229), .A2(new_n257), .A3(new_n212), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n255), .B1(new_n259), .B2(new_n190), .ZN(new_n260));
  INV_X1    g074(.A(new_n241), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT29), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(G472), .B1(new_n247), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(G472), .A2(G902), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n213), .A2(new_n223), .A3(KEYINPUT30), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n257), .B1(new_n229), .B2(new_n212), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n190), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(new_n230), .A3(new_n241), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT31), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n260), .A2(new_n271), .A3(new_n241), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n241), .B1(new_n251), .B2(new_n252), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT32), .B(new_n265), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT70), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n265), .B1(new_n273), .B2(new_n274), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT67), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT67), .B(new_n265), .C1(new_n273), .C2(new_n274), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT68), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT68), .ZN(new_n284));
  AOI211_X1 g098(.A(new_n284), .B(KEYINPUT32), .C1(new_n279), .C2(new_n280), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n264), .B(new_n276), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n287));
  INV_X1    g101(.A(G953), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(G221), .A3(G234), .ZN(new_n289));
  OR2_X1    g103(.A1(new_n289), .A2(KEYINPUT22), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(KEYINPUT22), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(G137), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(G137), .B1(new_n290), .B2(new_n291), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n287), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n294), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT71), .A3(new_n292), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n300), .A2(KEYINPUT16), .A3(G140), .ZN(new_n301));
  XNOR2_X1  g115(.A(G125), .B(G140), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(KEYINPUT16), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(G146), .ZN(new_n304));
  INV_X1    g118(.A(G119), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G128), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n305), .A2(KEYINPUT23), .A3(G128), .ZN(new_n309));
  OAI22_X1  g123(.A1(new_n308), .A2(new_n309), .B1(G119), .B2(new_n208), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n208), .A2(G119), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(new_n306), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT24), .B(G110), .Z(new_n313));
  AOI22_X1  g127(.A1(new_n310), .A2(G110), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n303), .A2(G146), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n302), .A2(new_n203), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI22_X1  g131(.A1(new_n310), .A2(G110), .B1(new_n312), .B2(new_n313), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n304), .A2(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT72), .B1(new_n299), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n304), .A2(new_n314), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n317), .A2(new_n318), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n298), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n319), .A2(new_n292), .A3(new_n296), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G217), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(G234), .B2(new_n245), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n327), .A2(G902), .A3(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n320), .A2(new_n324), .A3(new_n245), .A4(new_n326), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n331), .A2(KEYINPUT73), .A3(KEYINPUT25), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT25), .B1(new_n331), .B2(KEYINPUT73), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n330), .B1(new_n334), .B2(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n286), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G478), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(KEYINPUT15), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n208), .A2(G143), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n205), .A2(G128), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n192), .ZN(new_n342));
  INV_X1    g156(.A(G122), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G116), .ZN(new_n344));
  INV_X1    g158(.A(G116), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G122), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G107), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n351));
  INV_X1    g165(.A(new_n339), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n340), .B1(new_n351), .B2(new_n352), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT93), .A3(new_n339), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n342), .B(new_n349), .C1(new_n357), .C2(new_n192), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n343), .A2(G116), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT14), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n344), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT95), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g177(.A(KEYINPUT95), .B(new_n344), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n363), .B(new_n364), .C1(KEYINPUT14), .C2(new_n346), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G107), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n347), .A2(new_n348), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT94), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n341), .B(new_n192), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n358), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT9), .B(G234), .Z(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n373), .A2(new_n328), .A3(G953), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n358), .A2(new_n370), .A3(new_n374), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(KEYINPUT96), .A3(new_n377), .ZN(new_n378));
  OR3_X1    g192(.A1(new_n371), .A2(KEYINPUT96), .A3(new_n375), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(new_n245), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n338), .B1(new_n380), .B2(KEYINPUT97), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(KEYINPUT97), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n378), .A2(new_n379), .A3(new_n383), .A4(new_n245), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n381), .B1(new_n385), .B2(new_n338), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n237), .A2(G237), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n388));
  OAI211_X1 g202(.A(G214), .B(new_n288), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n205), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n239), .A2(G143), .A3(G214), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n196), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT87), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  INV_X1    g209(.A(new_n391), .ZN(new_n396));
  AOI21_X1  g210(.A(G143), .B1(new_n239), .B2(G214), .ZN(new_n397));
  OAI21_X1  g211(.A(G131), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n390), .A2(KEYINPUT87), .A3(new_n391), .A4(new_n196), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n394), .A2(new_n395), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n304), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT89), .B1(new_n398), .B2(new_n395), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n390), .A2(new_n391), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT17), .A4(G131), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n400), .A2(new_n401), .A3(new_n402), .A4(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(KEYINPUT18), .A3(G131), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n302), .A2(new_n203), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT86), .A3(new_n316), .ZN(new_n409));
  NAND2_X1  g223(.A1(KEYINPUT18), .A2(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n390), .A2(new_n391), .A3(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n408), .A2(KEYINPUT86), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n407), .A2(new_n409), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n415));
  XOR2_X1   g229(.A(G113), .B(G122), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT88), .ZN(new_n417));
  INV_X1    g231(.A(G104), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n406), .A2(new_n413), .A3(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT91), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n419), .B1(new_n406), .B2(new_n413), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n245), .B(new_n421), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G475), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n394), .A2(new_n398), .A3(new_n399), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n302), .B(KEYINPUT19), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n203), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(new_n315), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n420), .ZN(new_n432));
  AOI21_X1  g246(.A(G475), .B1(new_n432), .B2(new_n422), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(KEYINPUT90), .A3(new_n434), .A4(new_n245), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G952), .A3(new_n288), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT21), .B(G898), .Z(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G475), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n406), .A2(new_n413), .A3(new_n419), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n419), .B1(new_n430), .B2(new_n413), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n443), .B(new_n245), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT20), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n433), .A2(new_n434), .A3(new_n245), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND4_X1   g264(.A1(new_n386), .A2(new_n437), .A3(new_n442), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n221), .A2(new_n202), .A3(G128), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n210), .A3(new_n209), .ZN(new_n453));
  INV_X1    g267(.A(G101), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n418), .A2(G107), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n348), .A2(G104), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT3), .B1(new_n418), .B2(G107), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n348), .A3(G104), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n459), .A2(new_n461), .A3(new_n454), .A4(new_n455), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT75), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n462), .A2(new_n463), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n453), .B(new_n458), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT10), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n459), .A2(new_n461), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n468), .A2(KEYINPUT75), .A3(new_n454), .A4(new_n455), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n463), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n457), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT10), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n453), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n227), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n459), .A2(new_n461), .A3(new_n455), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G101), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT4), .B(new_n477), .C1(new_n464), .C2(new_n465), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n477), .A2(KEYINPUT4), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n228), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n474), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G140), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n288), .A2(G227), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n482), .B(new_n483), .Z(new_n484));
  AND2_X1   g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n466), .A2(KEYINPUT10), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n472), .B1(new_n471), .B2(new_n453), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n227), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n474), .A2(new_n475), .A3(new_n480), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n458), .B1(new_n464), .B2(new_n465), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n210), .A3(new_n209), .A4(new_n452), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n466), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n227), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(KEYINPUT12), .A3(new_n227), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n491), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n484), .B(KEYINPUT74), .Z(new_n500));
  OAI211_X1 g314(.A(new_n490), .B(G469), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(G469), .A2(G902), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n484), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n475), .B1(new_n474), .B2(new_n480), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n504), .B1(new_n491), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n489), .A2(new_n481), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT77), .A3(new_n504), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT76), .B1(new_n491), .B2(new_n504), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n497), .A2(new_n498), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT76), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n481), .A2(new_n514), .A3(new_n484), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G469), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n503), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G221), .B1(new_n373), .B2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT78), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT77), .B1(new_n509), .B2(new_n504), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n507), .B(new_n484), .C1(new_n489), .C2(new_n481), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(new_n518), .A3(new_n245), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT12), .B1(new_n494), .B2(new_n227), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n496), .B(new_n475), .C1(new_n493), .C2(new_n466), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n481), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n500), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n529), .A2(new_n530), .B1(new_n485), .B2(new_n489), .ZN(new_n531));
  OAI21_X1  g345(.A(G469), .B1(new_n531), .B2(G902), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n520), .ZN(new_n535));
  OAI21_X1  g349(.A(G214), .B1(G237), .B2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT6), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n187), .A2(KEYINPUT5), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n345), .A2(KEYINPUT5), .A3(G119), .ZN(new_n540));
  INV_X1    g354(.A(G113), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n539), .A2(new_n542), .B1(new_n225), .B2(new_n187), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n543), .B(new_n458), .C1(new_n464), .C2(new_n465), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT80), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT80), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n471), .A2(new_n546), .A3(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n478), .A2(new_n190), .A3(new_n479), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT79), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n478), .A2(KEYINPUT79), .A3(new_n190), .A4(new_n479), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(G110), .B(G122), .Z(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n538), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n551), .A2(new_n552), .ZN(new_n557));
  INV_X1    g371(.A(new_n548), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n554), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n220), .A2(G125), .A3(new_n222), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(KEYINPUT83), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT83), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n453), .B2(G125), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n288), .A2(G224), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT84), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n566), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT82), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n570), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NOR4_X1   g388(.A1(new_n553), .A2(KEYINPUT82), .A3(new_n555), .A4(new_n572), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n561), .B(new_n569), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n553), .A2(new_n555), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n567), .A2(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n565), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n566), .A2(KEYINPUT7), .A3(new_n567), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT85), .B1(new_n471), .B2(new_n543), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n471), .B2(new_n543), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n554), .B(KEYINPUT8), .Z(new_n583));
  INV_X1    g397(.A(KEYINPUT85), .ZN(new_n584));
  OR3_X1    g398(.A1(new_n471), .A2(new_n584), .A3(new_n543), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n577), .A2(new_n579), .A3(new_n580), .A4(new_n586), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n587), .A2(new_n245), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(G210), .B1(G237), .B2(G902), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n576), .A2(new_n588), .A3(new_n590), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n537), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n451), .A2(new_n522), .A3(new_n535), .A4(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n336), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(new_n454), .ZN(G3));
  OAI21_X1  g411(.A(new_n245), .B1(new_n273), .B2(new_n274), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT98), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT98), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(new_n245), .C1(new_n273), .C2(new_n274), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(G472), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n602), .A2(new_n335), .A3(new_n281), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n522), .A2(new_n535), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n437), .A2(new_n450), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n376), .A2(new_n607), .A3(new_n377), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n376), .B1(new_n607), .B2(new_n377), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT33), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n378), .A2(new_n379), .A3(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n610), .A2(G478), .A3(new_n245), .A4(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT100), .B(G478), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n380), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n606), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n576), .A2(new_n588), .A3(new_n590), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n590), .B1(new_n576), .B2(new_n588), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n536), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n442), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n617), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n605), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT34), .B(G104), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  XOR2_X1   g439(.A(new_n442), .B(KEYINPUT101), .Z(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n536), .B(new_n627), .C1(new_n618), .C2(new_n619), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n385), .A2(new_n338), .ZN(new_n629));
  INV_X1    g443(.A(new_n381), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n447), .A2(new_n449), .B1(new_n425), .B2(G475), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n604), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(KEYINPUT35), .B(G107), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND2_X1  g450(.A1(new_n334), .A2(new_n329), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n298), .A2(KEYINPUT36), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(new_n319), .Z(new_n639));
  OAI211_X1 g453(.A(new_n639), .B(new_n245), .C1(new_n328), .C2(G234), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT102), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n602), .A2(new_n281), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n595), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT37), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G110), .ZN(G12));
  AOI21_X1  g461(.A(new_n534), .B1(new_n533), .B2(new_n520), .ZN(new_n648));
  AOI211_X1 g462(.A(KEYINPUT78), .B(new_n521), .C1(new_n526), .C2(new_n532), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n439), .B1(new_n441), .B2(G900), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n631), .A2(new_n632), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n620), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n650), .A2(new_n286), .A3(new_n653), .A4(new_n642), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  XOR2_X1   g469(.A(new_n651), .B(KEYINPUT39), .Z(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT40), .Z(new_n659));
  NOR2_X1   g473(.A1(new_n260), .A2(new_n261), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n245), .B1(new_n231), .B2(new_n241), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G472), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n276), .B(new_n663), .C1(new_n283), .C2(new_n285), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n643), .A2(new_n536), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n386), .B1(new_n437), .B2(new_n450), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n592), .A2(new_n593), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT103), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n659), .A2(new_n665), .A3(new_n666), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  AND3_X1   g485(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n616), .B(new_n651), .C1(new_n672), .C2(new_n436), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT104), .B1(new_n620), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n650), .A2(new_n674), .A3(new_n286), .A4(new_n642), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n620), .A2(new_n673), .A3(KEYINPUT104), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n203), .ZN(G48));
  NAND2_X1  g492(.A1(new_n525), .A2(new_n245), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G469), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n520), .A3(new_n526), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n622), .A2(new_n286), .A3(new_n335), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  INV_X1    g498(.A(new_n628), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n286), .A2(new_n335), .A3(new_n685), .A4(new_n681), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(new_n633), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  NAND3_X1  g502(.A1(new_n680), .A2(new_n520), .A3(new_n526), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n620), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n286), .A2(new_n690), .A3(new_n642), .A4(new_n451), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT105), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NAND2_X1  g507(.A1(new_n598), .A2(G472), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n241), .B1(new_n232), .B2(new_n243), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n265), .B1(new_n273), .B2(new_n695), .ZN(new_n696));
  AND4_X1   g510(.A1(new_n335), .A2(new_n627), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n681), .A2(new_n697), .A3(new_n594), .A4(new_n666), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n690), .A2(KEYINPUT106), .A3(new_n666), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT107), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n343), .ZN(G24));
  NAND2_X1  g518(.A1(new_n694), .A2(new_n696), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n673), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n690), .A2(new_n642), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  XOR2_X1   g522(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n709));
  NOR2_X1   g523(.A1(new_n519), .A2(new_n521), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n592), .A2(new_n536), .A3(new_n593), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n286), .A2(new_n335), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n709), .B1(new_n713), .B2(new_n673), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n277), .A2(new_n282), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n264), .A2(new_n275), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n716), .A2(new_n335), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n711), .A2(new_n673), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n710), .A4(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT109), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n714), .A2(KEYINPUT109), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  NOR2_X1   g539(.A1(new_n713), .A2(new_n652), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n192), .ZN(G36));
  NOR2_X1   g541(.A1(new_n672), .A2(new_n436), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n616), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n729), .B(new_n730), .C1(KEYINPUT110), .C2(new_n606), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n728), .B(new_n616), .C1(new_n732), .C2(KEYINPUT43), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n644), .A3(new_n642), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n531), .A2(KEYINPUT45), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n531), .A2(KEYINPUT45), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(G469), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT46), .B1(new_n740), .B2(new_n502), .ZN(new_n741));
  INV_X1    g555(.A(new_n526), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(KEYINPUT46), .A3(new_n502), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n520), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n656), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n735), .A2(new_n736), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n737), .A2(new_n712), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G137), .ZN(G39));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n745), .A2(new_n752), .A3(new_n520), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n752), .B1(new_n745), .B2(new_n520), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n755), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(KEYINPUT47), .A3(new_n753), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n286), .ZN(new_n760));
  INV_X1    g574(.A(new_n335), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n718), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT112), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(KEYINPUT112), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  INV_X1    g580(.A(new_n669), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n680), .A2(new_n526), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT114), .Z(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT49), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n761), .A2(new_n521), .A3(new_n537), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n729), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n771), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n664), .B1(KEYINPUT113), .B2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n767), .A2(new_n770), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n761), .A2(new_n705), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n439), .B1(new_n731), .B2(new_n733), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT117), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n778), .A2(KEYINPUT117), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n681), .B(new_n777), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(G952), .B(new_n288), .C1(new_n782), .C2(new_n620), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n711), .A2(new_n689), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n785), .A2(new_n664), .A3(new_n761), .A4(new_n439), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT120), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT120), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n606), .A2(new_n616), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n784), .B1(new_n780), .B2(new_n781), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n643), .A3(new_n705), .ZN(new_n792));
  INV_X1    g606(.A(new_n777), .ZN(new_n793));
  INV_X1    g607(.A(new_n781), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(new_n779), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n669), .A2(new_n536), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT50), .A4(new_n681), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n767), .A2(new_n537), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n799), .B2(new_n782), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n790), .B(new_n792), .C1(new_n797), .C2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n795), .A2(new_n712), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n769), .A2(new_n521), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n756), .A2(new_n758), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n783), .B1(new_n801), .B2(new_n806), .ZN(new_n807));
  XOR2_X1   g621(.A(new_n804), .B(KEYINPUT119), .Z(new_n808));
  AND3_X1   g622(.A1(new_n756), .A2(new_n758), .A3(KEYINPUT118), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT118), .B1(new_n756), .B2(new_n758), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n803), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n792), .B1(new_n800), .B2(new_n797), .ZN(new_n813));
  INV_X1    g627(.A(new_n790), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n802), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n698), .A2(new_n699), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n698), .A2(new_n699), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n817), .A2(new_n818), .B1(new_n633), .B2(new_n686), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n682), .A2(new_n691), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n714), .A2(KEYINPUT109), .A3(new_n719), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT109), .B1(new_n714), .B2(new_n719), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n604), .A2(new_n617), .A3(new_n628), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT115), .B1(new_n596), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n617), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n650), .A2(new_n827), .A3(new_n603), .A4(new_n685), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n828), .B(new_n829), .C1(new_n336), .C2(new_n595), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n726), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n706), .A2(new_n710), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n632), .A2(new_n651), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n650), .A2(new_n286), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n835), .B2(new_n631), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n642), .A3(new_n712), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n606), .A2(new_n386), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n650), .A2(new_n838), .A3(new_n603), .A4(new_n685), .ZN(new_n839));
  INV_X1    g653(.A(new_n644), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n650), .A2(new_n451), .A3(new_n594), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(new_n643), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n831), .A2(new_n832), .A3(new_n837), .A4(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n824), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n654), .B(new_n707), .C1(new_n675), .C2(new_n676), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n664), .A2(new_n637), .A3(new_n640), .A4(new_n651), .ZN(new_n849));
  INV_X1    g663(.A(new_n710), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n594), .A2(new_n666), .ZN(new_n851));
  OR3_X1    g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n847), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n846), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n858));
  INV_X1    g672(.A(new_n707), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n286), .A2(new_n650), .A3(new_n674), .A4(new_n642), .ZN(new_n860));
  INV_X1    g674(.A(new_n676), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(KEYINPUT52), .A3(new_n852), .A4(new_n654), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n855), .B1(new_n847), .B2(new_n854), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(KEYINPUT116), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n845), .A2(new_n857), .A3(new_n858), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n864), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n687), .A2(new_n682), .A3(new_n691), .A4(new_n702), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n722), .B2(new_n723), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n726), .B(new_n842), .C1(new_n826), .C2(new_n830), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n867), .A2(new_n869), .A3(new_n837), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n866), .A2(new_n872), .A3(KEYINPUT54), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n858), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n720), .A2(KEYINPUT53), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n844), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n857), .A3(new_n821), .A4(new_n865), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n874), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n807), .A2(new_n816), .A3(new_n873), .A4(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n787), .A2(new_n788), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n881), .A2(new_n827), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n717), .B(new_n784), .C1(new_n780), .C2(new_n781), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT48), .Z(new_n884));
  NOR3_X1   g698(.A1(new_n880), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(G952), .A2(G953), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n776), .B1(new_n885), .B2(new_n886), .ZN(G75));
  OAI21_X1  g701(.A(new_n561), .B1(new_n574), .B2(new_n575), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n569), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n875), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n870), .A2(new_n821), .A3(new_n837), .A4(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n863), .A2(KEYINPUT116), .A3(new_n864), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT116), .B1(new_n863), .B2(new_n864), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n845), .B2(new_n867), .ZN(new_n896));
  OAI211_X1 g710(.A(G210), .B(G902), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT55), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n897), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n898), .B1(new_n897), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n890), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(G210), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n905), .B(new_n245), .C1(new_n874), .C2(new_n877), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT55), .B1(new_n906), .B2(new_n900), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n897), .A2(new_n898), .A3(new_n901), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n889), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n288), .A2(G952), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT122), .Z(new_n911));
  AND3_X1   g725(.A1(new_n904), .A2(new_n909), .A3(new_n911), .ZN(G51));
  NAND2_X1  g726(.A1(new_n874), .A2(new_n877), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(KEYINPUT123), .A3(new_n879), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n916), .A3(KEYINPUT54), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n502), .B(KEYINPUT57), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n525), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n895), .A2(new_n896), .ZN(new_n921));
  OR3_X1    g735(.A1(new_n921), .A2(new_n245), .A3(new_n740), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n910), .B1(new_n920), .B2(new_n922), .ZN(G54));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n245), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n422), .A3(new_n432), .ZN(new_n926));
  INV_X1    g740(.A(new_n910), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n432), .A2(new_n422), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .A4(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n873), .B2(new_n879), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n610), .A2(new_n612), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n911), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n915), .A2(new_n917), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n932), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n935), .B1(new_n937), .B2(new_n934), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT124), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n913), .A2(new_n639), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n911), .ZN(new_n943));
  AOI22_X1  g757(.A1(new_n913), .A2(new_n941), .B1(new_n326), .B2(new_n325), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g760(.A(new_n288), .B1(new_n440), .B2(G224), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n821), .A2(new_n843), .A3(new_n831), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n288), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n888), .B1(G898), .B2(new_n288), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n949), .B(new_n951), .ZN(G69));
  XNOR2_X1  g766(.A(new_n259), .B(new_n428), .ZN(new_n953));
  NAND2_X1  g767(.A1(G900), .A2(G953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n737), .A2(new_n712), .A3(new_n748), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n717), .A2(new_n594), .A3(new_n666), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n747), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n847), .A2(new_n726), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n724), .A3(new_n765), .A4(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n953), .B(new_n954), .C1(new_n960), .C2(G953), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n670), .A2(new_n848), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n827), .A2(new_n838), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n658), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n336), .A2(new_n711), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n967), .B(new_n968), .C1(new_n965), .C2(new_n966), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n749), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n964), .A2(new_n765), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n971), .A2(new_n288), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n961), .B1(new_n972), .B2(new_n953), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n288), .B1(G227), .B2(G900), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n974), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n961), .B(new_n976), .C1(new_n972), .C2(new_n953), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n971), .B2(new_n948), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n660), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n960), .B2(new_n948), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n983), .A2(new_n260), .A3(new_n261), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n982), .A2(new_n927), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n980), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n660), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n866), .A2(new_n262), .A3(new_n872), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(G57));
endmodule


