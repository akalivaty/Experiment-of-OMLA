//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n820, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G169gat), .ZN(new_n212));
  INV_X1    g011(.A(G176gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n211), .A2(new_n217), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  AND2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT24), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(new_n225), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(KEYINPUT23), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n218), .A2(KEYINPUT25), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT64), .B(KEYINPUT23), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(new_n214), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n228), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n223), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n207), .A2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(new_n208), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT28), .A3(new_n208), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n247), .A3(new_n231), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n214), .A2(KEYINPUT26), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n218), .A3(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n246), .A2(new_n250), .A3(KEYINPUT67), .A4(new_n204), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n225), .B1(new_n243), .B2(new_n245), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT67), .B1(new_n253), .B2(new_n250), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n203), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT72), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G197gat), .B(G204gat), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G211gat), .B(G218gat), .Z(new_n263));
  OR2_X1    g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n263), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n246), .A2(new_n250), .A3(new_n204), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(new_n251), .A3(new_n237), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT72), .A3(new_n203), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n237), .A2(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n202), .B1(new_n272), .B2(KEYINPUT29), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n257), .A2(new_n266), .A3(new_n271), .A4(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n203), .A2(KEYINPUT29), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n270), .A2(new_n275), .B1(new_n272), .B2(new_n203), .ZN(new_n276));
  INV_X1    g075(.A(new_n266), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT73), .ZN(new_n280));
  XOR2_X1   g079(.A(G64gat), .B(G92gat), .Z(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n274), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT75), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n274), .A2(KEYINPUT75), .A3(new_n278), .A4(new_n282), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n274), .A2(new_n278), .A3(new_n282), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n278), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n282), .B(KEYINPUT74), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n289), .A2(KEYINPUT30), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n294));
  OR2_X1    g093(.A1(G127gat), .A2(G134gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n296), .A2(new_n297), .B1(G127gat), .B2(G134gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n295), .B(new_n298), .C1(new_n299), .C2(KEYINPUT1), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n295), .ZN(new_n301));
  INV_X1    g100(.A(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G113gat), .ZN(new_n303));
  INV_X1    g102(.A(G113gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G120gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT1), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n300), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G148gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT76), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G148gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n312), .A3(G141gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G141gat), .B2(new_n309), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT77), .ZN(new_n315));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(KEYINPUT2), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n315), .A3(KEYINPUT2), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G155gat), .B(G162gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G155gat), .ZN(new_n323));
  INV_X1    g122(.A(G162gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(G141gat), .B(G148gat), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n316), .B(new_n325), .C1(new_n326), .C2(KEYINPUT2), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n308), .A2(new_n322), .A3(KEYINPUT4), .A4(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT4), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n316), .A2(new_n315), .A3(KEYINPUT2), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n321), .B1(new_n330), .B2(new_n317), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n309), .A2(G141gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT76), .B(G148gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(G141gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n327), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n300), .A2(new_n307), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n329), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n328), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n335), .A2(KEYINPUT3), .B1(new_n307), .B2(new_n300), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n342), .B(new_n327), .C1(new_n331), .C2(new_n334), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n341), .B1(new_n340), .B2(new_n343), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n339), .B(KEYINPUT5), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G57gat), .B(G85gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT80), .ZN(new_n348));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n328), .A2(new_n337), .A3(new_n338), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(new_n343), .A3(new_n336), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(KEYINPUT78), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n335), .B(new_n336), .ZN(new_n360));
  INV_X1    g159(.A(new_n338), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n346), .B(new_n352), .C1(new_n358), .C2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n366));
  INV_X1    g165(.A(new_n362), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n352), .B1(new_n368), .B2(new_n346), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n294), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n352), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n358), .A2(new_n362), .ZN(new_n372));
  INV_X1    g171(.A(new_n346), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n374), .A2(KEYINPUT81), .A3(new_n364), .A4(new_n363), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n376));
  OR3_X1    g175(.A1(new_n363), .A2(new_n376), .A3(new_n364), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n376), .B1(new_n363), .B2(new_n364), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n370), .A2(new_n375), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n293), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n343), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n277), .A2(new_n382), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n383), .A2(KEYINPUT83), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n342), .B1(new_n277), .B2(KEYINPUT29), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n335), .ZN(new_n386));
  NAND2_X1  g185(.A1(G228gat), .A2(G233gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n383), .A2(KEYINPUT83), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n384), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n266), .A2(KEYINPUT84), .A3(new_n381), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT84), .B1(new_n266), .B2(new_n381), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n342), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n382), .B(KEYINPUT85), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n392), .A2(new_n335), .B1(new_n277), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n389), .B1(new_n394), .B2(new_n387), .ZN(new_n395));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT31), .B(G50gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G22gat), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n389), .B(new_n399), .C1(new_n394), .C2(new_n387), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n380), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n336), .B1(new_n252), .B2(new_n254), .ZN(new_n406));
  INV_X1    g205(.A(G227gat), .ZN(new_n407));
  INV_X1    g206(.A(G233gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n269), .A2(new_n308), .A3(new_n251), .A4(new_n237), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT69), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n410), .B1(new_n406), .B2(new_n411), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(KEYINPUT33), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT32), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n411), .ZN(new_n424));
  AOI221_X4 g223(.A(new_n421), .B1(KEYINPUT33), .B2(new_n418), .C1(new_n424), .C2(new_n409), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n414), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n409), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n427), .A2(KEYINPUT32), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n418), .ZN(new_n431));
  INV_X1    g230(.A(new_n413), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n412), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n422), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n426), .A2(new_n435), .A3(KEYINPUT36), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT36), .B1(new_n426), .B2(new_n435), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n404), .A2(new_n405), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n403), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n293), .B2(new_n379), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n436), .A2(new_n437), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT86), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n282), .B1(new_n290), .B2(KEYINPUT37), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT87), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n274), .B2(new_n278), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n448), .B2(new_n282), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n274), .A2(new_n447), .A3(new_n278), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT38), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  INV_X1    g254(.A(new_n450), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n444), .B2(KEYINPUT87), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n457), .B2(new_n449), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT88), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n374), .A2(new_n364), .A3(new_n363), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n377), .A2(new_n460), .A3(new_n378), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n447), .B1(new_n276), .B2(new_n266), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n257), .A2(new_n271), .A3(new_n273), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(new_n266), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(new_n450), .A3(new_n455), .A4(new_n291), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n285), .A3(new_n287), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n454), .A2(new_n459), .A3(new_n467), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n337), .B(new_n328), .C1(new_n344), .C2(new_n345), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n361), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT39), .ZN(new_n471));
  INV_X1    g270(.A(new_n360), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(new_n338), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n352), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n469), .A2(new_n471), .A3(new_n361), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(KEYINPUT40), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n363), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT40), .B1(new_n474), .B2(new_n475), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n288), .A2(new_n292), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n403), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n439), .A2(new_n443), .B1(new_n468), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n426), .A2(new_n435), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(new_n403), .ZN(new_n484));
  XOR2_X1   g283(.A(KEYINPUT89), .B(KEYINPUT35), .Z(new_n485));
  AND3_X1   g284(.A1(new_n484), .A2(new_n461), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n379), .A3(new_n293), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n486), .A2(new_n293), .B1(new_n487), .B2(KEYINPUT35), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT90), .B1(new_n482), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n467), .B1(new_n458), .B2(KEYINPUT88), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n452), .A2(new_n453), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n481), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n405), .B1(new_n404), .B2(new_n438), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT86), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n486), .A2(new_n293), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n487), .A2(KEYINPUT35), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(G183gat), .B(G211gat), .Z(new_n502));
  INV_X1    g301(.A(KEYINPUT98), .ZN(new_n503));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G71gat), .B(G78gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT21), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT99), .ZN(new_n511));
  INV_X1    g310(.A(G231gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n408), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT99), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n510), .B(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(G231gat), .A3(G233gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G127gat), .B(G155gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(new_n516), .A3(new_n518), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n523), .B1(new_n520), .B2(new_n521), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n527));
  XOR2_X1   g326(.A(G15gat), .B(G22gat), .Z(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(G1gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n527), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n508), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(KEYINPUT21), .B2(new_n538), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n525), .A2(new_n526), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n539), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n520), .A2(new_n521), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n522), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n543), .B2(new_n524), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n502), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n539), .B1(new_n525), .B2(new_n526), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(new_n541), .A3(new_n524), .ZN(new_n547));
  INV_X1    g346(.A(new_n502), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G43gat), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT15), .B1(new_n551), .B2(G50gat), .ZN(new_n552));
  INV_X1    g351(.A(G50gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(G43gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OR3_X1    g354(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  INV_X1    g359(.A(G29gat), .ZN(new_n561));
  INV_X1    g360(.A(G36gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n555), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n555), .A2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n556), .A2(new_n558), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT92), .B(G43gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n554), .B1(new_n568), .B2(new_n553), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n565), .B(new_n566), .C1(new_n569), .C2(KEYINPUT15), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT7), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT8), .ZN(new_n574));
  AND2_X1   g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  OAI221_X1 g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .C1(G85gat), .C2(G92gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G99gat), .B(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n576), .B(new_n577), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT100), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n571), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT101), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n564), .A2(new_n570), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n581), .A2(KEYINPUT100), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n584), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n588), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT101), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n597), .B(KEYINPUT102), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n590), .A2(KEYINPUT17), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT93), .B(KEYINPUT17), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n571), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n591), .A2(new_n592), .A3(new_n599), .A4(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n596), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(new_n596), .B2(new_n602), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT103), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n606), .B(new_n607), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n593), .A2(KEYINPUT101), .A3(new_n594), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n602), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n598), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n598), .A3(new_n602), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n605), .A2(new_n609), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n614), .A2(new_n615), .A3(new_n608), .A4(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n536), .A2(KEYINPUT95), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n621), .A2(new_n599), .A3(new_n601), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n590), .A2(new_n536), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT18), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n624), .B(KEYINPUT13), .Z(new_n630));
  NOR2_X1   g429(.A1(new_n626), .A2(KEYINPUT97), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT97), .B1(new_n590), .B2(new_n536), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n625), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n630), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n628), .B1(new_n627), .B2(KEYINPUT96), .ZN(new_n636));
  XNOR2_X1  g435(.A(G113gat), .B(G141gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT11), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(new_n212), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G197gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT12), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n635), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n635), .B2(new_n636), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI211_X1 g446(.A(KEYINPUT10), .B(new_n538), .C1(new_n582), .C2(new_n585), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n581), .A2(new_n508), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n583), .A2(new_n538), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n648), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n650), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n653), .B1(new_n654), .B2(new_n647), .ZN(new_n655));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n550), .A2(new_n620), .A3(new_n645), .A4(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n501), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n379), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n529), .ZN(G1324gat));
  NAND3_X1  g467(.A1(new_n501), .A2(new_n480), .A3(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(G8gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT42), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT16), .B(G8gat), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g472(.A(new_n671), .B(KEYINPUT42), .S(new_n673), .Z(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n666), .B2(new_n438), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n483), .A2(G15gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n666), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n666), .A2(new_n440), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n620), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n489), .A2(new_n500), .A3(KEYINPUT44), .A4(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n645), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n550), .A2(new_n683), .A3(new_n662), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n441), .A2(new_n442), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n492), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n499), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n681), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n682), .A2(new_n684), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n379), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n682), .A2(new_n690), .A3(KEYINPUT106), .A4(new_n684), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT107), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n693), .A2(new_n698), .A3(new_n694), .A4(new_n695), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n697), .A2(G29gat), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n501), .A2(new_n681), .A3(new_n684), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n694), .A2(new_n561), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT105), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n700), .A2(new_n706), .ZN(G1328gat));
  NAND2_X1  g506(.A1(new_n480), .A2(new_n562), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT46), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n693), .A2(new_n480), .A3(new_n695), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n562), .B2(new_n711), .ZN(G1329gat));
  OAI21_X1  g511(.A(new_n568), .B1(new_n691), .B2(new_n438), .ZN(new_n713));
  INV_X1    g512(.A(new_n483), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n567), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n713), .B(KEYINPUT47), .C1(new_n701), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n715), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n693), .A2(new_n442), .A3(new_n695), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n568), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n719), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g519(.A(G50gat), .B1(new_n691), .B2(new_n440), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n403), .A2(new_n553), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n721), .B(KEYINPUT48), .C1(new_n701), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n701), .A2(new_n722), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n693), .A2(new_n403), .A3(new_n695), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(G50gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n723), .B1(new_n726), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g526(.A1(new_n545), .A2(new_n549), .ZN(new_n728));
  NOR4_X1   g527(.A1(new_n728), .A2(new_n681), .A3(new_n645), .A4(new_n663), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n687), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n694), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g533(.A(new_n293), .B(KEYINPUT109), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT110), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n738), .B(new_n740), .ZN(G1333gat));
  NAND3_X1  g540(.A1(new_n732), .A2(G71gat), .A3(new_n442), .ZN(new_n742));
  INV_X1    g541(.A(G71gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n731), .B2(new_n483), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n742), .A2(KEYINPUT50), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT50), .B1(new_n742), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1334gat));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n403), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g548(.A1(new_n550), .A2(new_n645), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n687), .A2(KEYINPUT51), .A3(new_n681), .A4(new_n750), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n751), .A2(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(KEYINPUT111), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n687), .A2(new_n681), .A3(new_n750), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n752), .A2(new_n753), .A3(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n663), .A2(G85gat), .A3(new_n379), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n682), .A2(new_n662), .A3(new_n690), .A4(new_n750), .ZN(new_n760));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760), .B2(new_n379), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n759), .A2(new_n761), .ZN(G1336gat));
  NOR3_X1   g561(.A1(new_n736), .A2(G92gat), .A3(new_n663), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G92gat), .B1(new_n760), .B2(new_n736), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n760), .A2(new_n293), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n756), .A2(new_n751), .ZN(new_n769));
  AOI22_X1  g568(.A1(new_n768), .A2(G92gat), .B1(new_n769), .B2(new_n763), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n770), .B2(new_n766), .ZN(G1337gat));
  XOR2_X1   g570(.A(KEYINPUT112), .B(G99gat), .Z(new_n772));
  NAND4_X1  g571(.A1(new_n757), .A2(new_n714), .A3(new_n662), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n760), .A2(new_n438), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n772), .ZN(G1338gat));
  OR2_X1    g574(.A1(new_n760), .A2(new_n440), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n663), .A2(G106gat), .A3(new_n440), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT53), .B1(new_n757), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n776), .A2(G106gat), .B1(new_n769), .B2(new_n778), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n648), .A2(new_n652), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n646), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n648), .A2(new_n652), .A3(new_n647), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n786), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n659), .B1(new_n653), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n661), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT55), .B1(new_n788), .B2(new_n790), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n645), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n631), .A2(new_n633), .A3(new_n630), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n624), .B1(new_n623), .B2(new_n626), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n640), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n662), .A2(new_n643), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(new_n620), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n793), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n661), .A3(new_n791), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n643), .A2(new_n799), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n619), .B(new_n618), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(new_n728), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n550), .A2(new_n683), .A3(new_n620), .A4(new_n663), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n379), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(new_n736), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n484), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n645), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n784), .B1(new_n812), .B2(G113gat), .ZN(new_n813));
  AOI211_X1 g612(.A(KEYINPUT113), .B(new_n304), .C1(new_n811), .C2(new_n645), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n645), .A2(new_n304), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  OAI22_X1  g615(.A1(new_n813), .A2(new_n814), .B1(new_n810), .B2(new_n816), .ZN(G1340gat));
  NOR2_X1   g616(.A1(new_n810), .A2(new_n663), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(new_n302), .ZN(G1341gat));
  NAND2_X1  g618(.A1(new_n811), .A2(new_n550), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g620(.A1(new_n620), .A2(new_n480), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n808), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(G134gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n484), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n810), .B2(new_n620), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1343gat));
  AOI211_X1 g632(.A(KEYINPUT57), .B(new_n440), .C1(new_n806), .C2(new_n807), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n438), .A2(new_n694), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(new_n735), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(G141gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n683), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n728), .A2(new_n681), .A3(new_n645), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n841), .A2(new_n663), .B1(new_n806), .B2(KEYINPUT117), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n801), .A2(new_n728), .A3(new_n843), .A4(new_n805), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n440), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n838), .B(new_n840), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n442), .A2(new_n440), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n808), .A2(new_n736), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n839), .B1(new_n849), .B2(new_n683), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n847), .A2(KEYINPUT58), .A3(new_n850), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n853), .B1(new_n855), .B2(new_n856), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n806), .A2(new_n807), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n403), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT57), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n858), .A2(new_n846), .A3(new_n403), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n836), .B(KEYINPUT119), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n860), .A2(new_n662), .A3(new_n861), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G148gat), .B1(new_n863), .B2(KEYINPUT120), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n846), .B1(new_n858), .B2(new_n403), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n834), .A3(new_n663), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(new_n862), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT59), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n333), .A2(KEYINPUT59), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n838), .B1(new_n845), .B2(new_n846), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n663), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n849), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n333), .A3(new_n662), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1345gat));
  OAI21_X1  g675(.A(G155gat), .B1(new_n871), .B2(new_n728), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n874), .A2(new_n323), .A3(new_n550), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1346gat));
  NAND3_X1  g678(.A1(new_n823), .A2(new_n324), .A3(new_n848), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n806), .A2(KEYINPUT117), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n807), .A3(new_n844), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n846), .B1(new_n882), .B2(new_n403), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n861), .A2(new_n836), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n883), .A2(new_n884), .A3(new_n620), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n885), .B2(new_n324), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n694), .A2(new_n293), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n858), .A2(new_n484), .A3(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(new_n212), .A3(new_n683), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n858), .B2(new_n379), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT122), .B(new_n694), .C1(new_n806), .C2(new_n807), .ZN(new_n894));
  OR2_X1    g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n484), .A3(new_n735), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n645), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n891), .B1(new_n898), .B2(new_n212), .ZN(G1348gat));
  OAI21_X1  g698(.A(G176gat), .B1(new_n890), .B2(new_n663), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n662), .A2(new_n213), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n896), .B2(new_n901), .ZN(G1349gat));
  OAI21_X1  g701(.A(G183gat), .B1(new_n890), .B2(new_n728), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n550), .A2(new_n244), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n896), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g705(.A1(new_n897), .A2(new_n208), .A3(new_n681), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n620), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT61), .B1(new_n908), .B2(new_n208), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G190gat), .B1(new_n890), .B2(new_n620), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(KEYINPUT61), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n909), .A2(new_n910), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(G1351gat));
  OAI211_X1 g714(.A(new_n735), .B(new_n848), .C1(new_n893), .C2(new_n894), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n683), .A2(G197gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n919), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n889), .A2(new_n438), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n860), .A2(new_n645), .A3(new_n861), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(G197gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n920), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT125), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n920), .A2(new_n929), .A3(new_n926), .A4(new_n922), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1352gat));
  NOR3_X1   g730(.A1(new_n916), .A2(G204gat), .A3(new_n663), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT62), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n867), .A2(new_n924), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G204gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1353gat));
  INV_X1    g735(.A(G211gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n937), .A3(new_n550), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n860), .A2(new_n550), .A3(new_n861), .A4(new_n924), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n866), .A2(new_n834), .A3(new_n923), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n937), .B1(new_n942), .B2(new_n550), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(KEYINPUT63), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n938), .B1(new_n944), .B2(new_n945), .ZN(G1354gat));
  NAND2_X1  g745(.A1(new_n942), .A2(new_n681), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G218gat), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n620), .A2(G218gat), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n917), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n948), .A2(KEYINPUT127), .A3(new_n950), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1355gat));
endmodule


