//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(G15gat), .ZN(new_n208));
  INV_X1    g007(.A(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G15gat), .A2(G22gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT16), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(G1gat), .ZN(new_n214));
  INV_X1    g013(.A(G1gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n210), .A2(new_n215), .A3(new_n211), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(G8gat), .B1(new_n216), .B2(KEYINPUT86), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n214), .B(new_n216), .C1(KEYINPUT86), .C2(G8gat), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT87), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n220), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT87), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT83), .B(G43gat), .Z(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT84), .B(G50gat), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n226), .A2(G50gat), .B1(new_n227), .B2(G43gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229));
  OR2_X1    g028(.A1(G43gat), .A2(G50gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(G43gat), .A2(G50gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT14), .ZN(new_n233));
  INV_X1    g032(.A(G29gat), .ZN(new_n234));
  INV_X1    g033(.A(G36gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n236), .A2(new_n237), .B1(G29gat), .B2(G36gat), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n228), .A2(new_n229), .B1(new_n232), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT85), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(G29gat), .A2(G36gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT85), .B1(new_n242), .B2(new_n233), .ZN(new_n243));
  OAI22_X1  g042(.A1(new_n241), .A2(new_n243), .B1(new_n234), .B2(new_n235), .ZN(new_n244));
  INV_X1    g043(.A(new_n232), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n239), .A2(KEYINPUT17), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT17), .B1(new_n239), .B2(new_n246), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n223), .B(new_n225), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G229gat), .A2(G233gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n221), .A2(new_n246), .A3(new_n239), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n207), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n246), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT88), .B1(new_n257), .B2(new_n224), .ZN(new_n258));
  OR2_X1    g057(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n250), .B(KEYINPUT13), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n251), .A2(new_n258), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n249), .A2(KEYINPUT18), .A3(new_n250), .A4(new_n251), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n254), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n256), .A2(new_n265), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269));
  INV_X1    g068(.A(G85gat), .ZN(new_n270));
  INV_X1    g069(.A(G92gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(KEYINPUT8), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT7), .ZN(new_n273));
  OAI22_X1  g072(.A1(new_n270), .A2(new_n271), .B1(new_n273), .B2(KEYINPUT97), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT97), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n275), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n272), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G99gat), .B(G106gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n272), .A2(new_n278), .A3(new_n274), .A4(new_n276), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT98), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n280), .A2(KEYINPUT98), .A3(new_n281), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n284), .A2(new_n285), .A3(new_n246), .A4(new_n239), .ZN(new_n286));
  AND3_X1   g085(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  AND3_X1   g087(.A1(new_n286), .A2(KEYINPUT99), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT99), .B1(new_n286), .B2(new_n288), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n247), .A2(new_n248), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n284), .A2(new_n285), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  OAI22_X1  g092(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT101), .ZN(new_n295));
  XOR2_X1   g094(.A(G190gat), .B(G218gat), .Z(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n295), .B1(new_n294), .B2(new_n297), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n286), .A2(new_n288), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT99), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n286), .A2(KEYINPUT99), .A3(new_n288), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n247), .A2(new_n248), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n303), .A2(new_n304), .B1(new_n292), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n296), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT96), .B(G134gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(G162gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n310));
  XOR2_X1   g109(.A(new_n309), .B(new_n310), .Z(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n300), .B(new_n307), .C1(KEYINPUT100), .C2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G57gat), .B(G64gat), .Z(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT90), .ZN(new_n315));
  XNOR2_X1  g114(.A(G57gat), .B(G64gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT90), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(KEYINPUT9), .A3(new_n318), .ZN(new_n319));
  OR2_X1    g118(.A1(G71gat), .A2(G78gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(G71gat), .A2(G78gat), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n314), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT91), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n314), .A3(KEYINPUT91), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(KEYINPUT95), .B(G183gat), .Z(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  NAND2_X1  g136(.A1(G231gat), .A2(G233gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n224), .B1(new_n331), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(G211gat), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n319), .A2(new_n322), .B1(new_n328), .B2(new_n329), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT21), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n342), .B1(new_n344), .B2(new_n224), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n338), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(G211gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(new_n342), .A3(new_n224), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(G231gat), .A3(new_n348), .A4(G233gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G127gat), .B(G155gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n346), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n353), .B1(new_n346), .B2(new_n349), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n337), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n335), .B(new_n336), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n354), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT101), .B1(new_n306), .B2(new_n296), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(new_n363), .A3(new_n307), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n362), .A2(KEYINPUT100), .A3(new_n363), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n311), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n313), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT102), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT102), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n313), .A2(new_n361), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n378), .A2(new_n379), .B1(KEYINPUT23), .B2(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(KEYINPUT23), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT25), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT67), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT65), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(KEYINPUT65), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n378), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT66), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT66), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n393), .A3(new_n378), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  OAI211_X1 g195(.A(KEYINPUT25), .B(new_n396), .C1(new_n380), .C2(KEYINPUT23), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n380), .A2(KEYINPUT64), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT64), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(G169gat), .B2(G176gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n397), .B1(new_n401), .B2(KEYINPUT23), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n386), .B1(new_n395), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n390), .A2(new_n393), .A3(new_n378), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n393), .B1(new_n390), .B2(new_n378), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n386), .B(new_n402), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n385), .B1(new_n403), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT27), .B(G183gat), .ZN(new_n409));
  INV_X1    g208(.A(G190gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT28), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT68), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT26), .B1(new_n398), .B2(new_n400), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT26), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n396), .B1(new_n380), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n413), .B(new_n377), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n377), .B1(new_n414), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT68), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n412), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n422), .B(KEYINPUT75), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT67), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n384), .B1(new_n429), .B2(new_n406), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n427), .B1(new_n430), .B2(new_n420), .ZN(new_n431));
  AND2_X1   g230(.A1(G211gat), .A2(G218gat), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(KEYINPUT22), .ZN(new_n433));
  NOR2_X1   g232(.A1(KEYINPUT71), .A2(G204gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(KEYINPUT71), .A2(G204gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n203), .A3(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(KEYINPUT71), .A2(G204gat), .ZN(new_n438));
  OAI21_X1  g237(.A(G197gat), .B1(new_n438), .B2(new_n434), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n433), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(G211gat), .A2(G218gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G211gat), .A2(G218gat), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT72), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT72), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n432), .B2(new_n441), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n441), .ZN(new_n449));
  AOI211_X1 g248(.A(new_n433), .B(new_n449), .C1(new_n437), .C2(new_n439), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT73), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT73), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n440), .B2(new_n447), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n425), .A2(new_n431), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT74), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n451), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n451), .B2(new_n453), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n431), .B2(new_n425), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n374), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n457), .A2(new_n458), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n408), .A2(new_n421), .B1(new_n426), .B2(new_n424), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n430), .A2(new_n420), .A3(new_n423), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n374), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n425), .A2(new_n431), .A3(new_n454), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(KEYINPUT30), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n465), .A2(new_n470), .A3(new_n466), .A4(new_n467), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(G127gat), .B(G134gat), .Z(new_n475));
  XNOR2_X1  g274(.A(G113gat), .B(G120gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(KEYINPUT1), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G113gat), .B(G120gat), .Z(new_n478));
  INV_X1    g277(.A(KEYINPUT1), .ZN(new_n479));
  XNOR2_X1  g278(.A(G127gat), .B(G134gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G141gat), .B(G148gat), .Z(new_n483));
  NAND2_X1  g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT2), .ZN(new_n485));
  INV_X1    g284(.A(G155gat), .ZN(new_n486));
  INV_X1    g285(.A(G162gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n484), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G141gat), .B(G148gat), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n484), .B(new_n488), .C1(new_n491), .C2(KEYINPUT2), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n490), .A2(new_n477), .A3(new_n481), .A4(new_n492), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n474), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT76), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT4), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n482), .B2(new_n493), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n473), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n490), .A2(new_n492), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT3), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n477), .A2(new_n481), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n492), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n495), .A2(KEYINPUT76), .A3(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT5), .B(new_n497), .C1(new_n502), .C2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(G1gat), .B(G29gat), .Z(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n515));
  OR2_X1    g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G57gat), .B(G85gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n519), .A3(new_n517), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n474), .A2(KEYINPUT5), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n508), .B(new_n524), .C1(new_n501), .C2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT80), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n523), .B1(new_n511), .B2(new_n526), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n528), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n472), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n429), .A2(new_n406), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n420), .B1(new_n540), .B2(new_n385), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT69), .B1(new_n541), .B2(new_n482), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n543));
  NOR4_X1   g342(.A1(new_n430), .A2(new_n543), .A3(new_n505), .A4(new_n420), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G227gat), .A2(G233gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n505), .B1(new_n430), .B2(new_n420), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n545), .A2(KEYINPUT34), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n408), .A2(new_n482), .A3(new_n421), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(new_n543), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n408), .A2(KEYINPUT69), .A3(new_n482), .A4(new_n421), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n550), .A2(new_n546), .A3(new_n547), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT34), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n539), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT32), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n550), .A2(new_n547), .A3(new_n551), .ZN(new_n558));
  INV_X1    g357(.A(new_n546), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT33), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G43gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(G71gat), .B(G99gat), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  AOI221_X4 g365(.A(new_n557), .B1(KEYINPUT33), .B2(new_n564), .C1(new_n558), .C2(new_n559), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n556), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n482), .B1(new_n408), .B2(new_n421), .ZN(new_n569));
  NOR3_X1   g368(.A1(new_n542), .A2(new_n544), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT32), .B1(new_n570), .B2(new_n546), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n570), .B2(new_n546), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n573), .A3(new_n564), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n560), .B1(new_n561), .B2(new_n565), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n548), .A2(new_n539), .A3(new_n554), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n555), .ZN(new_n577));
  XOR2_X1   g376(.A(G78gat), .B(G106gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT81), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT31), .B(G50gat), .Z(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G228gat), .A2(G233gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n454), .A2(new_n426), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n493), .B1(new_n584), .B2(new_n506), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n507), .A2(new_n426), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n587), .B1(new_n457), .B2(new_n458), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n583), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n440), .A2(new_n432), .A3(new_n441), .ZN(new_n590));
  INV_X1    g389(.A(new_n450), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT29), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n503), .B1(new_n592), .B2(KEYINPUT3), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n451), .A2(new_n453), .A3(new_n587), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n583), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n589), .A2(G22gat), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n588), .ZN(new_n598));
  OAI211_X1 g397(.A(G228gat), .B(G233gat), .C1(new_n598), .C2(new_n585), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n209), .B1(new_n599), .B2(new_n595), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n582), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(G22gat), .B1(new_n589), .B2(new_n596), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n209), .A3(new_n595), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n581), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  AND4_X1   g404(.A1(new_n538), .A2(new_n568), .A3(new_n577), .A4(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT35), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n469), .A2(new_n471), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n529), .A2(new_n534), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n609), .A2(new_n536), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT82), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n612), .A2(new_n577), .A3(new_n568), .A4(new_n605), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n607), .B1(new_n611), .B2(KEYINPUT82), .ZN(new_n614));
  OAI22_X1  g413(.A1(new_n606), .A2(new_n607), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n568), .A2(new_n577), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT36), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT39), .B(new_n473), .C1(new_n494), .C2(new_n496), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n508), .B1(new_n501), .B2(new_n525), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT39), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n523), .B(new_n618), .C1(new_n620), .C2(new_n473), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n469), .A2(new_n534), .A3(new_n471), .A4(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n621), .A2(new_n622), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n454), .B1(new_n425), .B2(new_n431), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT37), .B1(new_n465), .B2(new_n467), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n626), .B(new_n374), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n468), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n536), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n629), .B1(new_n455), .B2(new_n460), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n465), .A2(KEYINPUT37), .A3(new_n467), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n466), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n634), .B1(new_n637), .B2(new_n626), .ZN(new_n638));
  OAI221_X1 g437(.A(new_n605), .B1(new_n624), .B2(new_n625), .C1(new_n633), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n605), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n537), .B2(new_n472), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT36), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n568), .A2(new_n577), .A3(new_n642), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n617), .A2(new_n639), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n268), .B(new_n371), .C1(new_n615), .C2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(G230gat), .ZN(new_n646));
  INV_X1    g445(.A(G233gat), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n282), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n280), .A2(KEYINPUT103), .A3(new_n281), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n331), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n343), .A2(new_n650), .A3(new_n282), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n292), .A2(new_n656), .A3(new_n331), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n649), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n654), .A3(new_n648), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n658), .B2(new_n659), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n645), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n537), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n268), .B1(new_n615), .B2(new_n644), .ZN(new_n673));
  INV_X1    g472(.A(new_n371), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n673), .A2(new_n668), .A3(new_n472), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT16), .B(G8gat), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(KEYINPUT42), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n675), .A2(G8gat), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n645), .A2(new_n668), .A3(new_n472), .A4(new_n678), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT42), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n672), .B1(new_n680), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n681), .B2(new_n682), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(new_n679), .A3(KEYINPUT104), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(new_n616), .ZN(new_n690));
  AOI21_X1  g489(.A(G15gat), .B1(new_n669), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n617), .A2(new_n643), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n208), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n669), .B2(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n669), .A2(new_n640), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  NAND2_X1  g497(.A1(new_n615), .A2(new_n644), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n256), .B(new_n265), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n361), .A2(new_n667), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n313), .A2(new_n366), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT105), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n703), .A2(KEYINPUT105), .ZN(new_n705));
  AND4_X1   g504(.A1(new_n699), .A2(new_n700), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n234), .A3(new_n537), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n699), .B2(new_n702), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n364), .A2(new_n365), .A3(new_n311), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n364), .B1(new_n365), .B2(new_n311), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n714));
  AOI211_X1 g513(.A(new_n713), .B(new_n714), .C1(new_n615), .C2(new_n644), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n700), .B(new_n701), .C1(new_n710), .C2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n537), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n708), .A2(new_n718), .ZN(G1328gat));
  NAND3_X1  g518(.A1(new_n673), .A2(new_n704), .A3(new_n705), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G36gat), .A3(new_n608), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT46), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n716), .B2(new_n608), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1329gat));
  INV_X1    g523(.A(new_n226), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(new_n716), .B2(new_n693), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n706), .A2(KEYINPUT107), .A3(new_n690), .A4(new_n226), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n673), .A2(new_n690), .A3(new_n704), .A4(new_n705), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n725), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n726), .A2(KEYINPUT47), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1330gat));
  INV_X1    g535(.A(new_n227), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n605), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n714), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n699), .A2(new_n702), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n713), .B1(new_n615), .B2(new_n644), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(new_n709), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n742), .A2(new_n640), .A3(new_n700), .A4(new_n701), .ZN(new_n743));
  AOI211_X1 g542(.A(KEYINPUT48), .B(new_n738), .C1(new_n743), .C2(new_n737), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n737), .B1(new_n716), .B2(new_n605), .ZN(new_n746));
  INV_X1    g545(.A(new_n738), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n744), .A2(new_n748), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n371), .A2(new_n700), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n699), .A2(new_n667), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n717), .ZN(new_n752));
  XOR2_X1   g551(.A(new_n752), .B(G57gat), .Z(G1332gat));
  AOI21_X1  g552(.A(new_n668), .B1(new_n615), .B2(new_n644), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n754), .A2(KEYINPUT108), .A3(new_n750), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT108), .B1(new_n754), .B2(new_n750), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(new_n608), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  NOR3_X1   g561(.A1(new_n751), .A2(G71gat), .A3(new_n616), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n692), .B1(new_n755), .B2(new_n756), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n763), .B1(new_n764), .B2(G71gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI211_X1 g566(.A(KEYINPUT50), .B(new_n763), .C1(new_n764), .C2(G71gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(G1334gat));
  OAI21_X1  g568(.A(new_n640), .B1(new_n755), .B2(new_n756), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n700), .A2(new_n361), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g572(.A(new_n713), .B(new_n773), .C1(new_n615), .C2(new_n644), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n702), .A4(new_n772), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n741), .A2(new_n772), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n775), .A2(new_n778), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n781), .A2(new_n668), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n782), .A2(new_n270), .A3(new_n537), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n667), .B(new_n772), .C1(new_n710), .C2(new_n715), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n717), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1336gat));
  OAI21_X1  g585(.A(G92gat), .B1(new_n784), .B2(new_n608), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n788));
  NAND3_X1  g587(.A1(new_n472), .A2(new_n271), .A3(new_n667), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT110), .Z(new_n790));
  OAI211_X1 g589(.A(new_n787), .B(new_n788), .C1(new_n781), .C2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  OR2_X1    g591(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n793));
  NAND2_X1  g592(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n780), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT109), .B1(new_n774), .B2(KEYINPUT51), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n776), .A2(new_n777), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n790), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n742), .A2(new_n667), .A3(new_n472), .A4(new_n772), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(G92gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n791), .B1(new_n792), .B2(new_n801), .ZN(G1337gat));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(G99gat), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n782), .A2(new_n690), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n784), .B2(new_n693), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1338gat));
  OAI21_X1  g606(.A(G106gat), .B1(new_n784), .B2(new_n605), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n809));
  NOR3_X1   g608(.A1(new_n605), .A2(G106gat), .A3(new_n668), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT114), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n808), .B(new_n809), .C1(new_n781), .C2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n811), .B(KEYINPUT115), .Z(new_n814));
  NAND4_X1  g613(.A1(new_n742), .A2(new_n667), .A3(new_n640), .A4(new_n772), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n798), .A2(new_n814), .B1(new_n815), .B2(G106gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n812), .B1(new_n813), .B2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(G113gat), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n254), .A2(new_n207), .A3(new_n263), .A4(new_n264), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n261), .B1(new_n259), .B2(new_n262), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n250), .B1(new_n249), .B2(new_n251), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n206), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n819), .B(new_n822), .C1(new_n665), .C2(new_n666), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n653), .A2(new_n654), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n656), .ZN(new_n826));
  INV_X1    g625(.A(new_n657), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n648), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n828), .A2(KEYINPUT54), .A3(new_n658), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n649), .C1(new_n655), .C2(new_n657), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n662), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n824), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n658), .A3(KEYINPUT54), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n662), .A4(new_n831), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n664), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n823), .B1(new_n268), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n713), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n819), .A2(new_n822), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n833), .A2(new_n664), .A3(new_n835), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n702), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n361), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n368), .A2(new_n668), .A3(new_n268), .A4(new_n370), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n717), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n616), .A2(new_n640), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n608), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n846), .A2(KEYINPUT117), .A3(new_n608), .A4(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n818), .B1(new_n852), .B2(new_n700), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  INV_X1    g654(.A(new_n848), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n268), .A2(G113gat), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT118), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n854), .A2(new_n855), .A3(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n859), .ZN(new_n861));
  OAI21_X1  g660(.A(KEYINPUT119), .B1(new_n853), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(G1340gat));
  INV_X1    g662(.A(new_n852), .ZN(new_n864));
  OAI21_X1  g663(.A(G120gat), .B1(new_n864), .B2(new_n668), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n668), .A2(G120gat), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT120), .Z(new_n867));
  OAI21_X1  g666(.A(new_n865), .B1(new_n848), .B2(new_n867), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n856), .A2(new_n869), .A3(new_n361), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n843), .B1(new_n850), .B2(new_n851), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n869), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n872), .B(new_n873), .ZN(G1342gat));
  NOR3_X1   g673(.A1(new_n848), .A2(G134gat), .A3(new_n713), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT56), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n864), .B2(new_n713), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1343gat));
  NOR3_X1   g677(.A1(new_n692), .A2(new_n717), .A3(new_n472), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  INV_X1    g679(.A(new_n845), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n361), .B1(new_n838), .B2(new_n841), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n640), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n823), .B(KEYINPUT122), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n835), .A2(new_n664), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n833), .A2(KEYINPUT123), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(new_n824), .C1(new_n829), .C2(new_n832), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n700), .A2(new_n885), .A3(new_n886), .A4(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n702), .B1(new_n884), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n841), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n843), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n605), .B1(new_n892), .B2(new_n845), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n879), .B(new_n883), .C1(new_n893), .C2(new_n880), .ZN(new_n894));
  OAI21_X1  g693(.A(G141gat), .B1(new_n894), .B2(new_n268), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n846), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n605), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n692), .B1(new_n846), .B2(new_n896), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n608), .A3(new_n899), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n268), .A2(G141gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n895), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT58), .B1(new_n895), .B2(KEYINPUT125), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI221_X1 g703(.A(new_n895), .B1(KEYINPUT125), .B2(KEYINPUT58), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(G1344gat));
  NOR2_X1   g705(.A1(new_n668), .A2(G148gat), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n898), .A2(new_n608), .A3(new_n899), .A4(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n909), .B(G148gat), .C1(new_n894), .C2(new_n668), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n840), .B1(new_n711), .B2(new_n712), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n702), .A2(new_n914), .A3(new_n840), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n839), .A3(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n890), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n361), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n880), .B(new_n640), .C1(new_n918), .C2(new_n881), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n640), .B1(new_n881), .B2(new_n882), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT57), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n919), .A2(new_n921), .A3(new_n667), .A4(new_n879), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n909), .B1(new_n922), .B2(G148gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n908), .B1(new_n911), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT127), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n926), .B(new_n908), .C1(new_n911), .C2(new_n923), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1345gat));
  NOR3_X1   g727(.A1(new_n894), .A2(new_n486), .A3(new_n843), .ZN(new_n929));
  INV_X1    g728(.A(new_n900), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n361), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n931), .B2(new_n486), .ZN(G1346gat));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n487), .A3(new_n702), .ZN(new_n933));
  OAI21_X1  g732(.A(G162gat), .B1(new_n894), .B2(new_n713), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1347gat));
  AOI211_X1 g734(.A(new_n616), .B(new_n640), .C1(new_n844), .C2(new_n845), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n537), .A2(new_n608), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n700), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n667), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(G176gat), .ZN(G1349gat));
  AND3_X1   g741(.A1(new_n936), .A2(new_n361), .A3(new_n937), .ZN(new_n943));
  INV_X1    g742(.A(G183gat), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n409), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1350gat));
  NAND2_X1  g750(.A1(new_n938), .A2(new_n702), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(new_n410), .ZN(new_n954));
  XOR2_X1   g753(.A(KEYINPUT61), .B(G190gat), .Z(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n952), .B2(new_n955), .ZN(G1351gat));
  NAND2_X1  g755(.A1(new_n693), .A2(new_n937), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n957), .A2(new_n920), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n203), .A3(new_n700), .ZN(new_n959));
  AND4_X1   g758(.A1(new_n693), .A2(new_n919), .A3(new_n921), .A4(new_n937), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(new_n700), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n959), .B1(new_n961), .B2(new_n203), .ZN(G1352gat));
  NOR4_X1   g761(.A1(new_n957), .A2(new_n920), .A3(G204gat), .A4(new_n668), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n919), .A2(new_n667), .A3(new_n921), .ZN(new_n965));
  OAI21_X1  g764(.A(G204gat), .B1(new_n965), .B2(new_n957), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n342), .A3(new_n361), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n960), .A2(new_n361), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  AOI21_X1  g771(.A(G218gat), .B1(new_n958), .B2(new_n702), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n702), .A2(G218gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n973), .B1(new_n960), .B2(new_n974), .ZN(G1355gat));
endmodule


