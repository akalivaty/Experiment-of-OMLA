

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757;

  XNOR2_X1 U367 ( .A(n513), .B(n512), .ZN(n729) );
  BUF_X1 U368 ( .A(G116), .Z(n401) );
  XNOR2_X1 U369 ( .A(G119), .B(G116), .ZN(n373) );
  AND2_X2 U370 ( .A1(n736), .A2(n437), .ZN(n376) );
  NAND2_X2 U371 ( .A1(n380), .A2(n379), .ZN(n368) );
  XNOR2_X1 U372 ( .A(G113), .B(KEYINPUT74), .ZN(n374) );
  NAND2_X2 U373 ( .A1(n393), .A2(n347), .ZN(n421) );
  AND2_X2 U374 ( .A1(n424), .A2(n423), .ZN(n422) );
  XNOR2_X1 U375 ( .A(n616), .B(KEYINPUT86), .ZN(n748) );
  INV_X1 U376 ( .A(n608), .ZN(n686) );
  NAND2_X1 U377 ( .A1(n539), .A2(n685), .ZN(n370) );
  NAND2_X1 U378 ( .A1(n408), .A2(n573), .ZN(n616) );
  OR2_X2 U379 ( .A1(n411), .A2(n413), .ZN(n539) );
  XNOR2_X1 U380 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U381 ( .A(n515), .B(n365), .ZN(n364) );
  INV_X2 U382 ( .A(G953), .ZN(n751) );
  INV_X2 U383 ( .A(KEYINPUT4), .ZN(n366) );
  XNOR2_X1 U384 ( .A(G113), .B(KEYINPUT74), .ZN(n477) );
  XNOR2_X1 U385 ( .A(KEYINPUT75), .B(KEYINPUT3), .ZN(n479) );
  NAND2_X1 U386 ( .A1(n442), .A2(n440), .ZN(n345) );
  NAND2_X1 U387 ( .A1(n442), .A2(n440), .ZN(n620) );
  XNOR2_X1 U388 ( .A(n390), .B(KEYINPUT32), .ZN(n346) );
  XNOR2_X1 U389 ( .A(n390), .B(KEYINPUT32), .ZN(n755) );
  XNOR2_X1 U390 ( .A(n364), .B(G137), .ZN(n361) );
  INV_X1 U391 ( .A(G472), .ZN(n436) );
  NOR2_X1 U392 ( .A1(n636), .A2(G902), .ZN(n482) );
  NAND2_X1 U393 ( .A1(n416), .A2(G902), .ZN(n414) );
  XNOR2_X1 U394 ( .A(n487), .B(n367), .ZN(n731) );
  INV_X1 U395 ( .A(G107), .ZN(n367) );
  XNOR2_X1 U396 ( .A(G104), .B(G110), .ZN(n487) );
  XNOR2_X1 U397 ( .A(n731), .B(KEYINPUT76), .ZN(n514) );
  INV_X1 U398 ( .A(KEYINPUT78), .ZN(n382) );
  XNOR2_X1 U399 ( .A(n460), .B(G128), .ZN(n419) );
  INV_X1 U400 ( .A(G143), .ZN(n460) );
  INV_X1 U401 ( .A(KEYINPUT48), .ZN(n430) );
  NAND2_X1 U402 ( .A1(G234), .A2(G237), .ZN(n508) );
  XNOR2_X1 U403 ( .A(n385), .B(n474), .ZN(n476) );
  XNOR2_X1 U404 ( .A(n473), .B(n386), .ZN(n385) );
  INV_X1 U405 ( .A(KEYINPUT80), .ZN(n386) );
  XNOR2_X1 U406 ( .A(n493), .B(n495), .ZN(n433) );
  XOR2_X1 U407 ( .A(G131), .B(G140), .Z(n488) );
  XNOR2_X1 U408 ( .A(n516), .B(G146), .ZN(n471) );
  XNOR2_X1 U409 ( .A(n525), .B(n524), .ZN(n643) );
  XNOR2_X1 U410 ( .A(n729), .B(n514), .ZN(n525) );
  AND2_X1 U411 ( .A1(n349), .A2(n675), .ZN(n427) );
  XNOR2_X1 U412 ( .A(n384), .B(n383), .ZN(n554) );
  INV_X1 U413 ( .A(KEYINPUT109), .ZN(n383) );
  XNOR2_X1 U414 ( .A(n435), .B(n535), .ZN(n434) );
  XNOR2_X1 U415 ( .A(n501), .B(n500), .ZN(n502) );
  INV_X1 U416 ( .A(KEYINPUT25), .ZN(n500) );
  XNOR2_X1 U417 ( .A(n690), .B(n356), .ZN(n357) );
  INV_X1 U418 ( .A(KEYINPUT6), .ZN(n356) );
  INV_X1 U419 ( .A(KEYINPUT1), .ZN(n420) );
  XNOR2_X1 U420 ( .A(n466), .B(n406), .ZN(n721) );
  XNOR2_X1 U421 ( .A(n468), .B(n362), .ZN(n406) );
  XNOR2_X1 U422 ( .A(n401), .B(G107), .ZN(n464) );
  INV_X1 U423 ( .A(KEYINPUT72), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n359) );
  INV_X1 U425 ( .A(G137), .ZN(n363) );
  NOR2_X1 U426 ( .A1(n399), .A2(n566), .ZN(n410) );
  NAND2_X1 U427 ( .A1(n491), .A2(n484), .ZN(n412) );
  XNOR2_X2 U428 ( .A(G119), .B(G116), .ZN(n478) );
  INV_X1 U429 ( .A(G134), .ZN(n461) );
  XNOR2_X1 U430 ( .A(G113), .B(G122), .ZN(n449) );
  XOR2_X1 U431 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n450) );
  XNOR2_X1 U432 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U433 ( .A(G143), .B(G104), .ZN(n452) );
  NOR2_X1 U434 ( .A1(G953), .A2(G237), .ZN(n472) );
  NAND2_X1 U435 ( .A1(n443), .A2(n441), .ZN(n440) );
  XOR2_X1 U436 ( .A(KEYINPUT70), .B(G101), .Z(n516) );
  XNOR2_X1 U437 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n519) );
  INV_X1 U438 ( .A(G237), .ZN(n483) );
  INV_X1 U439 ( .A(KEYINPUT38), .ZN(n387) );
  NAND2_X1 U440 ( .A1(n543), .A2(KEYINPUT89), .ZN(n423) );
  NOR2_X1 U441 ( .A1(n533), .A2(n534), .ZN(n540) );
  XNOR2_X1 U442 ( .A(KEYINPUT15), .B(G902), .ZN(n618) );
  XNOR2_X1 U443 ( .A(KEYINPUT16), .B(G122), .ZN(n512) );
  XNOR2_X1 U444 ( .A(n402), .B(n463), .ZN(n465) );
  XNOR2_X1 U445 ( .A(n462), .B(n403), .ZN(n402) );
  INV_X1 U446 ( .A(KEYINPUT101), .ZN(n403) );
  XNOR2_X1 U447 ( .A(n370), .B(n369), .ZN(n511) );
  INV_X1 U448 ( .A(KEYINPUT106), .ZN(n369) );
  XNOR2_X1 U449 ( .A(n405), .B(n404), .ZN(n653) );
  INV_X1 U450 ( .A(KEYINPUT103), .ZN(n404) );
  BUF_X1 U451 ( .A(n690), .Z(n400) );
  XNOR2_X1 U452 ( .A(n481), .B(n394), .ZN(n636) );
  XNOR2_X1 U453 ( .A(n432), .B(n431), .ZN(n725) );
  XNOR2_X1 U454 ( .A(n498), .B(n351), .ZN(n431) );
  XNOR2_X1 U455 ( .A(n497), .B(n433), .ZN(n432) );
  XNOR2_X1 U456 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U457 ( .A(n488), .B(n446), .ZN(n489) );
  AND2_X1 U458 ( .A1(G227), .A2(n751), .ZN(n446) );
  XNOR2_X1 U459 ( .A(n645), .B(n644), .ZN(n646) );
  AND2_X1 U460 ( .A1(n439), .A2(n438), .ZN(n710) );
  XNOR2_X1 U461 ( .A(n568), .B(n542), .ZN(n544) );
  NOR2_X1 U462 ( .A1(n554), .A2(n553), .ZN(n662) );
  XNOR2_X1 U463 ( .A(n723), .B(n722), .ZN(n398) );
  NOR2_X1 U464 ( .A1(n543), .A2(KEYINPUT89), .ZN(n347) );
  NOR2_X1 U465 ( .A1(n572), .A2(n653), .ZN(n348) );
  XOR2_X1 U466 ( .A(n486), .B(n485), .Z(n349) );
  XNOR2_X1 U467 ( .A(n529), .B(n528), .ZN(n350) );
  XNOR2_X1 U468 ( .A(n419), .B(n461), .ZN(n470) );
  INV_X1 U469 ( .A(n470), .ZN(n362) );
  XOR2_X1 U470 ( .A(n492), .B(n494), .Z(n351) );
  AND2_X1 U471 ( .A1(n736), .A2(n445), .ZN(n352) );
  XOR2_X1 U472 ( .A(KEYINPUT69), .B(KEYINPUT0), .Z(n353) );
  XNOR2_X1 U473 ( .A(n503), .B(n502), .ZN(n607) );
  INV_X1 U474 ( .A(n607), .ZN(n395) );
  INV_X1 U475 ( .A(G902), .ZN(n484) );
  XNOR2_X1 U476 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n354) );
  OR2_X1 U477 ( .A1(KEYINPUT44), .A2(KEYINPUT77), .ZN(n355) );
  INV_X1 U478 ( .A(n357), .ZN(n396) );
  NAND2_X1 U479 ( .A1(n541), .A2(n357), .ZN(n568) );
  NAND2_X1 U480 ( .A1(n396), .A2(n607), .ZN(n587) );
  NOR2_X1 U481 ( .A1(n609), .A2(n357), .ZN(n610) );
  NAND2_X2 U482 ( .A1(n360), .A2(n358), .ZN(n744) );
  NAND2_X1 U483 ( .A1(n359), .A2(n362), .ZN(n358) );
  NAND2_X1 U484 ( .A1(n361), .A2(n470), .ZN(n360) );
  XNOR2_X2 U485 ( .A(n744), .B(n471), .ZN(n394) );
  XNOR2_X2 U486 ( .A(n366), .B(KEYINPUT71), .ZN(n515) );
  XNOR2_X2 U487 ( .A(n368), .B(n479), .ZN(n513) );
  INV_X1 U488 ( .A(n370), .ZN(n594) );
  BUF_X1 U489 ( .A(n513), .Z(n371) );
  XNOR2_X1 U490 ( .A(n620), .B(n619), .ZN(n372) );
  XNOR2_X1 U491 ( .A(n345), .B(n619), .ZN(n720) );
  BUF_X2 U492 ( .A(n372), .Z(n724) );
  XNOR2_X1 U493 ( .A(n417), .B(KEYINPUT81), .ZN(n375) );
  XNOR2_X1 U494 ( .A(n417), .B(KEYINPUT81), .ZN(n428) );
  OR2_X2 U495 ( .A1(n599), .A2(n396), .ZN(n575) );
  BUF_X1 U496 ( .A(n643), .Z(n645) );
  XNOR2_X1 U497 ( .A(n391), .B(KEYINPUT35), .ZN(n641) );
  NAND2_X1 U498 ( .A1(n373), .A2(n374), .ZN(n379) );
  NAND2_X1 U499 ( .A1(n377), .A2(n378), .ZN(n380) );
  INV_X1 U500 ( .A(n478), .ZN(n377) );
  INV_X1 U501 ( .A(n477), .ZN(n378) );
  NAND2_X1 U502 ( .A1(n690), .A2(n540), .ZN(n435) );
  XNOR2_X2 U503 ( .A(n482), .B(n436), .ZN(n690) );
  NAND2_X1 U504 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U505 ( .A1(n567), .A2(n381), .ZN(n399) );
  XNOR2_X1 U506 ( .A(n565), .B(n382), .ZN(n381) );
  NAND2_X1 U507 ( .A1(n434), .A2(n539), .ZN(n384) );
  INV_X1 U508 ( .A(n388), .ZN(n393) );
  NAND2_X1 U509 ( .A1(n388), .A2(KEYINPUT89), .ZN(n424) );
  XNOR2_X2 U510 ( .A(n530), .B(n350), .ZN(n388) );
  XNOR2_X1 U511 ( .A(n393), .B(n387), .ZN(n675) );
  NOR2_X1 U512 ( .A1(n549), .A2(n388), .ZN(n550) );
  AND2_X1 U513 ( .A1(n388), .A2(n571), .ZN(n633) );
  NOR2_X2 U514 ( .A1(n641), .A2(n389), .ZN(n593) );
  NAND2_X1 U515 ( .A1(n592), .A2(n755), .ZN(n389) );
  NAND2_X2 U516 ( .A1(n611), .A2(n589), .ZN(n390) );
  NAND2_X1 U517 ( .A1(n392), .A2(n582), .ZN(n391) );
  XNOR2_X1 U518 ( .A(n581), .B(KEYINPUT34), .ZN(n392) );
  XNOR2_X1 U519 ( .A(n394), .B(n490), .ZN(n715) );
  XNOR2_X2 U520 ( .A(n397), .B(n353), .ZN(n601) );
  NOR2_X2 U521 ( .A1(n580), .A2(n579), .ZN(n397) );
  XNOR2_X2 U522 ( .A(n552), .B(n551), .ZN(n580) );
  NAND2_X2 U523 ( .A1(n422), .A2(n421), .ZN(n552) );
  NOR2_X2 U524 ( .A1(n596), .A2(n705), .ZN(n581) );
  XNOR2_X2 U525 ( .A(n601), .B(KEYINPUT93), .ZN(n596) );
  NAND2_X1 U526 ( .A1(n561), .A2(n562), .ZN(n563) );
  NOR2_X1 U527 ( .A1(n398), .A2(n728), .ZN(G63) );
  NOR2_X1 U528 ( .A1(n564), .A2(KEYINPUT47), .ZN(n565) );
  NAND2_X1 U529 ( .A1(n560), .A2(n662), .ZN(n564) );
  NAND2_X1 U530 ( .A1(n556), .A2(n555), .ZN(n405) );
  NAND2_X1 U531 ( .A1(n407), .A2(n410), .ZN(n409) );
  XNOR2_X1 U532 ( .A(n538), .B(KEYINPUT46), .ZN(n407) );
  NOR2_X1 U533 ( .A1(n572), .A2(n557), .ZN(n532) );
  XNOR2_X1 U534 ( .A(n429), .B(n531), .ZN(n572) );
  NAND2_X1 U535 ( .A1(n511), .A2(n510), .ZN(n417) );
  NAND2_X1 U536 ( .A1(n617), .A2(n736), .ZN(n443) );
  XNOR2_X2 U537 ( .A(n425), .B(n354), .ZN(n736) );
  XNOR2_X1 U538 ( .A(n409), .B(n430), .ZN(n408) );
  NOR2_X1 U539 ( .A1(n715), .A2(n412), .ZN(n411) );
  NAND2_X1 U540 ( .A1(n715), .A2(n416), .ZN(n415) );
  INV_X1 U541 ( .A(n491), .ZN(n416) );
  NAND2_X1 U542 ( .A1(n418), .A2(n375), .ZN(n634) );
  AND2_X1 U543 ( .A1(n550), .A2(n349), .ZN(n418) );
  XNOR2_X1 U544 ( .A(n419), .B(n517), .ZN(n521) );
  XNOR2_X2 U545 ( .A(n539), .B(n420), .ZN(n608) );
  NAND2_X1 U546 ( .A1(n426), .A2(n615), .ZN(n425) );
  XNOR2_X1 U547 ( .A(n593), .B(n355), .ZN(n426) );
  NAND2_X1 U548 ( .A1(n428), .A2(n427), .ZN(n429) );
  NAND2_X1 U549 ( .A1(n376), .A2(n444), .ZN(n442) );
  NOR2_X1 U550 ( .A1(n618), .A2(KEYINPUT2), .ZN(n437) );
  NAND2_X1 U551 ( .A1(n443), .A2(KEYINPUT2), .ZN(n438) );
  NAND2_X1 U552 ( .A1(n352), .A2(n444), .ZN(n439) );
  NOR2_X1 U553 ( .A1(n618), .A2(n445), .ZN(n441) );
  INV_X1 U554 ( .A(n748), .ZN(n444) );
  INV_X1 U555 ( .A(KEYINPUT2), .ZN(n445) );
  XNOR2_X2 U556 ( .A(n575), .B(n574), .ZN(n705) );
  OR2_X1 U557 ( .A1(n547), .A2(n556), .ZN(n447) );
  INV_X1 U558 ( .A(KEYINPUT100), .ZN(n451) );
  XNOR2_X1 U559 ( .A(n454), .B(n453), .ZN(n456) );
  INV_X1 U560 ( .A(KEYINPUT110), .ZN(n542) );
  INV_X1 U561 ( .A(KEYINPUT65), .ZN(n619) );
  BUF_X1 U562 ( .A(n580), .Z(n553) );
  XNOR2_X1 U563 ( .A(n715), .B(n716), .ZN(n717) );
  XNOR2_X1 U564 ( .A(n545), .B(KEYINPUT36), .ZN(n546) );
  XNOR2_X1 U565 ( .A(n718), .B(n717), .ZN(n719) );
  BUF_X1 U566 ( .A(n641), .Z(n642) );
  XNOR2_X1 U567 ( .A(KEYINPUT13), .B(G475), .ZN(n459) );
  INV_X1 U568 ( .A(G146), .ZN(n448) );
  XNOR2_X1 U569 ( .A(n448), .B(G125), .ZN(n517) );
  XNOR2_X1 U570 ( .A(n517), .B(KEYINPUT10), .ZN(n498) );
  XNOR2_X1 U571 ( .A(n488), .B(n498), .ZN(n745) );
  XNOR2_X1 U572 ( .A(n450), .B(n449), .ZN(n454) );
  NAND2_X1 U573 ( .A1(G214), .A2(n472), .ZN(n455) );
  XNOR2_X1 U574 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U575 ( .A(n745), .B(n457), .Z(n624) );
  NOR2_X1 U576 ( .A1(G902), .A2(n624), .ZN(n458) );
  XNOR2_X1 U577 ( .A(n459), .B(n458), .ZN(n547) );
  INV_X1 U578 ( .A(n547), .ZN(n555) );
  XOR2_X1 U579 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n463) );
  XNOR2_X1 U580 ( .A(G122), .B(KEYINPUT102), .ZN(n462) );
  XNOR2_X1 U581 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U582 ( .A1(G234), .A2(n751), .ZN(n467) );
  XOR2_X1 U583 ( .A(KEYINPUT8), .B(n467), .Z(n496) );
  NAND2_X1 U584 ( .A1(G217), .A2(n496), .ZN(n468) );
  NOR2_X1 U585 ( .A1(n721), .A2(G902), .ZN(n469) );
  XOR2_X1 U586 ( .A(n469), .B(G478), .Z(n556) );
  NOR2_X2 U587 ( .A1(n555), .A2(n556), .ZN(n664) );
  INV_X1 U588 ( .A(n664), .ZN(n557) );
  XOR2_X1 U589 ( .A(KEYINPUT107), .B(KEYINPUT30), .Z(n486) );
  XOR2_X1 U590 ( .A(KEYINPUT79), .B(KEYINPUT96), .Z(n474) );
  NAND2_X1 U591 ( .A1(n472), .A2(G210), .ZN(n473) );
  XNOR2_X1 U592 ( .A(G131), .B(KEYINPUT5), .ZN(n475) );
  XNOR2_X1 U593 ( .A(n476), .B(n475), .ZN(n480) );
  XNOR2_X1 U594 ( .A(n371), .B(n480), .ZN(n481) );
  NAND2_X1 U595 ( .A1(n484), .A2(n483), .ZN(n526) );
  NAND2_X1 U596 ( .A1(n526), .A2(G214), .ZN(n674) );
  NAND2_X1 U597 ( .A1(n690), .A2(n674), .ZN(n485) );
  XNOR2_X1 U598 ( .A(n514), .B(n489), .ZN(n490) );
  XNOR2_X1 U599 ( .A(KEYINPUT73), .B(G469), .ZN(n491) );
  XOR2_X1 U600 ( .A(G140), .B(G110), .Z(n493) );
  XNOR2_X1 U601 ( .A(G137), .B(G128), .ZN(n492) );
  XOR2_X1 U602 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n495) );
  XNOR2_X1 U603 ( .A(G119), .B(KEYINPUT94), .ZN(n494) );
  NAND2_X1 U604 ( .A1(n496), .A2(G221), .ZN(n497) );
  NOR2_X1 U605 ( .A1(G902), .A2(n725), .ZN(n503) );
  NAND2_X1 U606 ( .A1(G234), .A2(n618), .ZN(n499) );
  XNOR2_X1 U607 ( .A(KEYINPUT20), .B(n499), .ZN(n504) );
  NAND2_X1 U608 ( .A1(G217), .A2(n504), .ZN(n501) );
  NAND2_X1 U609 ( .A1(n504), .A2(G221), .ZN(n505) );
  XOR2_X1 U610 ( .A(KEYINPUT21), .B(n505), .Z(n683) );
  XNOR2_X1 U611 ( .A(KEYINPUT95), .B(n683), .ZN(n583) );
  NOR2_X1 U612 ( .A1(n607), .A2(n583), .ZN(n685) );
  NOR2_X1 U613 ( .A1(G900), .A2(n751), .ZN(n506) );
  NAND2_X1 U614 ( .A1(n506), .A2(G902), .ZN(n507) );
  NAND2_X1 U615 ( .A1(G952), .A2(n751), .ZN(n576) );
  NAND2_X1 U616 ( .A1(n507), .A2(n576), .ZN(n509) );
  XNOR2_X1 U617 ( .A(n508), .B(KEYINPUT14), .ZN(n701) );
  NAND2_X1 U618 ( .A1(n509), .A2(n701), .ZN(n534) );
  INV_X1 U619 ( .A(n534), .ZN(n510) );
  XNOR2_X1 U620 ( .A(n516), .B(n515), .ZN(n523) );
  NAND2_X1 U621 ( .A1(n751), .A2(G224), .ZN(n518) );
  XNOR2_X1 U622 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U624 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U625 ( .A1(n643), .A2(n618), .ZN(n530) );
  NAND2_X1 U626 ( .A1(n526), .A2(G210), .ZN(n529) );
  INV_X1 U627 ( .A(KEYINPUT83), .ZN(n527) );
  XNOR2_X1 U628 ( .A(n527), .B(KEYINPUT92), .ZN(n528) );
  XOR2_X1 U629 ( .A(KEYINPUT88), .B(KEYINPUT39), .Z(n531) );
  XNOR2_X1 U630 ( .A(n532), .B(KEYINPUT40), .ZN(n756) );
  XOR2_X1 U631 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n535) );
  NAND2_X1 U632 ( .A1(n607), .A2(n683), .ZN(n533) );
  NAND2_X1 U633 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U634 ( .A1(n447), .A2(n679), .ZN(n536) );
  XNOR2_X1 U635 ( .A(KEYINPUT41), .B(n536), .ZN(n704) );
  NOR2_X1 U636 ( .A1(n554), .A2(n704), .ZN(n537) );
  XNOR2_X1 U637 ( .A(KEYINPUT42), .B(n537), .ZN(n757) );
  NOR2_X1 U638 ( .A1(n756), .A2(n757), .ZN(n538) );
  AND2_X1 U639 ( .A1(n664), .A2(n540), .ZN(n541) );
  INV_X1 U640 ( .A(n674), .ZN(n543) );
  NAND2_X1 U641 ( .A1(n544), .A2(n552), .ZN(n545) );
  NOR2_X1 U642 ( .A1(n608), .A2(n546), .ZN(n673) );
  XNOR2_X1 U643 ( .A(n673), .B(KEYINPUT87), .ZN(n567) );
  NAND2_X1 U644 ( .A1(n556), .A2(n547), .ZN(n548) );
  XNOR2_X1 U645 ( .A(n548), .B(KEYINPUT105), .ZN(n582) );
  INV_X1 U646 ( .A(n582), .ZN(n549) );
  XOR2_X1 U647 ( .A(KEYINPUT85), .B(n634), .Z(n562) );
  XNOR2_X1 U648 ( .A(KEYINPUT68), .B(KEYINPUT19), .ZN(n551) );
  NAND2_X1 U649 ( .A1(n557), .A2(n653), .ZN(n559) );
  INV_X1 U650 ( .A(KEYINPUT104), .ZN(n558) );
  XNOR2_X1 U651 ( .A(n559), .B(n558), .ZN(n678) );
  INV_X1 U652 ( .A(n678), .ZN(n560) );
  NAND2_X1 U653 ( .A1(KEYINPUT47), .A2(n564), .ZN(n561) );
  XNOR2_X1 U654 ( .A(KEYINPUT84), .B(n563), .ZN(n566) );
  NOR2_X1 U655 ( .A1(n686), .A2(n568), .ZN(n569) );
  NAND2_X1 U656 ( .A1(n569), .A2(n674), .ZN(n570) );
  XNOR2_X1 U657 ( .A(KEYINPUT43), .B(n570), .ZN(n571) );
  NOR2_X1 U658 ( .A1(n633), .A2(n348), .ZN(n573) );
  NAND2_X1 U659 ( .A1(n686), .A2(n685), .ZN(n599) );
  INV_X1 U660 ( .A(KEYINPUT33), .ZN(n574) );
  NOR2_X1 U661 ( .A1(G898), .A2(n751), .ZN(n735) );
  NAND2_X1 U662 ( .A1(n735), .A2(G902), .ZN(n577) );
  NAND2_X1 U663 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U664 ( .A1(n701), .A2(n578), .ZN(n579) );
  NOR2_X1 U665 ( .A1(n583), .A2(n447), .ZN(n584) );
  NAND2_X1 U666 ( .A1(n601), .A2(n584), .ZN(n586) );
  XOR2_X1 U667 ( .A(KEYINPUT22), .B(KEYINPUT66), .Z(n585) );
  XNOR2_X2 U668 ( .A(n586), .B(n585), .ZN(n611) );
  NOR2_X1 U669 ( .A1(n608), .A2(n587), .ZN(n588) );
  XNOR2_X1 U670 ( .A(KEYINPUT82), .B(n588), .ZN(n589) );
  NAND2_X1 U671 ( .A1(n608), .A2(n607), .ZN(n590) );
  NOR2_X1 U672 ( .A1(n590), .A2(n400), .ZN(n591) );
  AND2_X1 U673 ( .A1(n611), .A2(n591), .ZN(n659) );
  INV_X1 U674 ( .A(n659), .ZN(n592) );
  INV_X1 U675 ( .A(n400), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n598), .A2(n594), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U678 ( .A(KEYINPUT97), .B(n597), .Z(n654) );
  OR2_X1 U679 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U680 ( .A(n600), .B(KEYINPUT98), .ZN(n694) );
  BUF_X1 U681 ( .A(n601), .Z(n602) );
  INV_X1 U682 ( .A(n602), .ZN(n603) );
  NOR2_X1 U683 ( .A1(n694), .A2(n603), .ZN(n605) );
  XNOR2_X1 U684 ( .A(KEYINPUT31), .B(KEYINPUT99), .ZN(n604) );
  XNOR2_X1 U685 ( .A(n605), .B(n604), .ZN(n667) );
  NOR2_X1 U686 ( .A1(n654), .A2(n667), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n606), .A2(n678), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n608), .A2(n395), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n651) );
  NAND2_X1 U690 ( .A1(KEYINPUT44), .A2(KEYINPUT77), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n651), .A2(n612), .ZN(n613) );
  NOR2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  INV_X1 U693 ( .A(n616), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n720), .A2(G475), .ZN(n626) );
  XOR2_X1 U695 ( .A(KEYINPUT90), .B(KEYINPUT122), .Z(n622) );
  XNOR2_X1 U696 ( .A(KEYINPUT59), .B(KEYINPUT67), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n626), .B(n625), .ZN(n630) );
  INV_X1 U699 ( .A(G952), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n627), .A2(G953), .ZN(n629) );
  INV_X1 U701 ( .A(KEYINPUT91), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(n714) );
  NAND2_X1 U703 ( .A1(n630), .A2(n714), .ZN(n632) );
  INV_X1 U704 ( .A(KEYINPUT60), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n632), .B(n631), .ZN(G60) );
  XOR2_X1 U706 ( .A(n633), .B(G140), .Z(G42) );
  XNOR2_X1 U707 ( .A(n634), .B(G143), .ZN(G45) );
  NAND2_X1 U708 ( .A1(n372), .A2(G472), .ZN(n638) );
  XNOR2_X1 U709 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n639), .A2(n714), .ZN(n640) );
  XNOR2_X1 U712 ( .A(n640), .B(KEYINPUT63), .ZN(G57) );
  XOR2_X1 U713 ( .A(n642), .B(G122), .Z(G24) );
  NAND2_X1 U714 ( .A1(n720), .A2(G210), .ZN(n647) );
  XOR2_X1 U715 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n644) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n648), .A2(n714), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT121), .B(KEYINPUT56), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(G51) );
  XNOR2_X1 U720 ( .A(G101), .B(n651), .ZN(G3) );
  NAND2_X1 U721 ( .A1(n664), .A2(n654), .ZN(n652) );
  XNOR2_X1 U722 ( .A(G104), .B(n652), .ZN(G6) );
  XNOR2_X1 U723 ( .A(KEYINPUT27), .B(KEYINPUT112), .ZN(n658) );
  XOR2_X1 U724 ( .A(G107), .B(KEYINPUT26), .Z(n656) );
  INV_X1 U725 ( .A(n653), .ZN(n666) );
  NAND2_X1 U726 ( .A1(n654), .A2(n666), .ZN(n655) );
  XNOR2_X1 U727 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(G9) );
  XOR2_X1 U729 ( .A(G110), .B(n659), .Z(G12) );
  XOR2_X1 U730 ( .A(G128), .B(KEYINPUT29), .Z(n661) );
  NAND2_X1 U731 ( .A1(n662), .A2(n666), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(G30) );
  NAND2_X1 U733 ( .A1(n662), .A2(n664), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(G146), .ZN(G48) );
  NAND2_X1 U735 ( .A1(n667), .A2(n664), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n665), .B(G113), .ZN(G15) );
  XOR2_X1 U737 ( .A(n401), .B(KEYINPUT113), .Z(n669) );
  NAND2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U739 ( .A(n669), .B(n668), .ZN(G18) );
  XOR2_X1 U740 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n671) );
  XNOR2_X1 U741 ( .A(G125), .B(KEYINPUT37), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n673), .B(n672), .ZN(G27) );
  XOR2_X1 U744 ( .A(G134), .B(n348), .Z(G36) );
  NOR2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n447), .A2(n676), .ZN(n677) );
  XOR2_X1 U747 ( .A(KEYINPUT117), .B(n677), .Z(n681) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U750 ( .A1(n705), .A2(n682), .ZN(n698) );
  NOR2_X1 U751 ( .A1(n395), .A2(n683), .ZN(n684) );
  XNOR2_X1 U752 ( .A(KEYINPUT49), .B(n684), .ZN(n692) );
  XOR2_X1 U753 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n688) );
  OR2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n400), .A2(n689), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U759 ( .A(KEYINPUT51), .B(n695), .ZN(n696) );
  NOR2_X1 U760 ( .A1(n696), .A2(n704), .ZN(n697) );
  NOR2_X1 U761 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U762 ( .A(KEYINPUT118), .B(KEYINPUT52), .ZN(n699) );
  XNOR2_X1 U763 ( .A(n700), .B(n699), .ZN(n703) );
  NAND2_X1 U764 ( .A1(n701), .A2(G952), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U766 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U767 ( .A(n706), .B(KEYINPUT119), .Z(n707) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U770 ( .A1(G953), .A2(n711), .ZN(n713) );
  XNOR2_X1 U771 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n713), .B(n712), .ZN(G75) );
  INV_X1 U773 ( .A(n714), .ZN(n728) );
  NAND2_X1 U774 ( .A1(n724), .A2(G469), .ZN(n718) );
  XOR2_X1 U775 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n716) );
  NOR2_X1 U776 ( .A1(n728), .A2(n719), .ZN(G54) );
  NAND2_X1 U777 ( .A1(n724), .A2(G478), .ZN(n723) );
  XOR2_X1 U778 ( .A(n721), .B(KEYINPUT123), .Z(n722) );
  NAND2_X1 U779 ( .A1(n724), .A2(G217), .ZN(n726) );
  XNOR2_X1 U780 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U781 ( .A1(n728), .A2(n727), .ZN(G66) );
  BUF_X1 U782 ( .A(n729), .Z(n730) );
  XNOR2_X1 U783 ( .A(n731), .B(KEYINPUT125), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n730), .B(n732), .ZN(n733) );
  XOR2_X1 U785 ( .A(G101), .B(n733), .Z(n734) );
  NOR2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n743) );
  NAND2_X1 U787 ( .A1(n736), .A2(n751), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n737), .B(KEYINPUT124), .ZN(n741) );
  NAND2_X1 U789 ( .A1(G953), .A2(G224), .ZN(n738) );
  XNOR2_X1 U790 ( .A(KEYINPUT61), .B(n738), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n739), .A2(G898), .ZN(n740) );
  NAND2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n744), .B(n745), .ZN(n749) );
  XNOR2_X1 U795 ( .A(G227), .B(n749), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U797 ( .A1(n747), .A2(G953), .ZN(n754) );
  XNOR2_X1 U798 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U799 ( .A(n750), .B(KEYINPUT126), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n754), .A2(n753), .ZN(G72) );
  XNOR2_X1 U802 ( .A(n346), .B(G119), .ZN(G21) );
  XOR2_X1 U803 ( .A(n756), .B(G131), .Z(G33) );
  XOR2_X1 U804 ( .A(G137), .B(n757), .Z(G39) );
endmodule

