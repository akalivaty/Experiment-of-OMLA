//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n206), .B2(G1gat), .ZN(new_n207));
  INV_X1    g006(.A(G8gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT89), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT88), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n212), .B(G8gat), .C1(KEYINPUT88), .C2(new_n204), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(G43gat), .B(G50gat), .Z(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n215), .A2(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT86), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT14), .ZN(new_n223));
  OR2_X1    g022(.A1(new_n222), .A2(KEYINPUT14), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n217), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n215), .A2(new_n216), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n226), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n228), .A2(new_n217), .A3(new_n223), .A4(new_n224), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(KEYINPUT17), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n229), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n213), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n231), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n237), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n236), .B(new_n231), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n235), .B(KEYINPUT13), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n241), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G197gat), .ZN(new_n247));
  XOR2_X1   g046(.A(KEYINPUT11), .B(G169gat), .Z(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT12), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n240), .A2(new_n250), .A3(new_n241), .A4(new_n244), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n252), .A2(KEYINPUT90), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT90), .B1(new_n252), .B2(new_n253), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT75), .ZN(new_n259));
  XOR2_X1   g058(.A(G57gat), .B(G85gat), .Z(new_n260));
  OR2_X1    g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n260), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n261), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267));
  INV_X1    g066(.A(G134gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G127gat), .ZN(new_n269));
  INV_X1    g068(.A(G127gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G134gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G113gat), .B(G120gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(KEYINPUT1), .ZN(new_n274));
  INV_X1    g073(.A(G120gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G113gat), .ZN(new_n276));
  INV_X1    g075(.A(G113gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G120gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(KEYINPUT72), .A2(G155gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(KEYINPUT72), .A2(G155gat), .ZN(new_n285));
  OAI21_X1  g084(.A(G162gat), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT2), .ZN(new_n287));
  OR2_X1    g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288));
  INV_X1    g087(.A(G162gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G155gat), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(G162gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293));
  AND4_X1   g092(.A1(new_n288), .A2(new_n290), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT2), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n288), .A2(new_n295), .A3(new_n293), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n290), .A2(new_n292), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n287), .A2(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT4), .B1(new_n283), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n297), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(G155gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n295), .B1(new_n301), .B2(G162gat), .ZN(new_n302));
  NAND4_X1  g101(.A1(new_n288), .A2(new_n290), .A3(new_n292), .A4(new_n293), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n274), .A2(new_n282), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n267), .B1(new_n299), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XOR2_X1   g109(.A(KEYINPUT73), .B(KEYINPUT3), .Z(new_n311));
  OAI211_X1 g110(.A(new_n300), .B(new_n311), .C1(new_n302), .C2(new_n303), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n312), .A2(new_n305), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n310), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT5), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n306), .B1(new_n304), .B2(new_n305), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n283), .A2(new_n298), .A3(KEYINPUT4), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT76), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n308), .A2(new_n315), .A3(new_n316), .A4(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n305), .A3(new_n312), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n321), .A2(new_n317), .A3(new_n318), .A4(new_n309), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n283), .A2(new_n298), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n305), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n316), .B1(new_n325), .B2(new_n310), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  AOI211_X1 g126(.A(KEYINPUT78), .B(new_n266), .C1(new_n320), .C2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n327), .ZN(new_n330));
  INV_X1    g129(.A(new_n266), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n320), .A2(new_n327), .A3(new_n266), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT6), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n334), .A2(KEYINPUT77), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT77), .B1(new_n334), .B2(new_n335), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n329), .B(new_n333), .C1(new_n336), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT79), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n266), .B1(new_n320), .B2(new_n327), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(new_n328), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n343), .B(new_n344), .C1(new_n337), .C2(new_n336), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(KEYINPUT6), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n339), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT23), .ZN(new_n351));
  XNOR2_X1  g150(.A(G183gat), .B(G190gat), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n349), .B(new_n351), .C1(new_n352), .C2(new_n348), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n354), .A2(new_n355), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n350), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT25), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(KEYINPUT27), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G183gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n365), .A3(new_n361), .ZN(new_n366));
  OR2_X1    g165(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n367));
  NAND2_X1  g166(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n362), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT26), .ZN(new_n371));
  INV_X1    g170(.A(G169gat), .ZN(new_n372));
  INV_X1    g171(.A(G176gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT67), .ZN(new_n375));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n371), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n373), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n350), .A2(new_n380), .A3(new_n371), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n375), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT27), .B(G183gat), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n383), .A2(new_n361), .A3(new_n367), .A4(new_n368), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n370), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n355), .A2(G176gat), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT25), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n376), .B1(KEYINPUT65), .B2(KEYINPUT23), .ZN(new_n391));
  INV_X1    g190(.A(new_n357), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n378), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n361), .A2(G183gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n360), .A2(G190gat), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT24), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n390), .A2(new_n393), .A3(new_n396), .A4(new_n349), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n359), .A2(new_n385), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n305), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n359), .A2(new_n385), .A3(new_n283), .A4(new_n397), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G227gat), .ZN(new_n402));
  INV_X1    g201(.A(G233gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT32), .ZN(new_n406));
  XNOR2_X1  g205(.A(G15gat), .B(G43gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G71gat), .B(G99gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT69), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n409), .B1(new_n405), .B2(KEYINPUT32), .ZN(new_n415));
  INV_X1    g214(.A(new_n410), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n401), .B2(new_n404), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n414), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n409), .ZN(new_n420));
  INV_X1    g219(.A(new_n404), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n421), .B1(new_n399), .B2(new_n400), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT32), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n424), .A2(KEYINPUT69), .A3(new_n417), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n413), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n399), .A2(new_n421), .A3(new_n400), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT34), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT31), .B(G50gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  XNOR2_X1  g231(.A(G197gat), .B(G204gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G211gat), .B(G218gat), .ZN(new_n434));
  INV_X1    g233(.A(G218gat), .ZN(new_n435));
  INV_X1    g234(.A(G211gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT70), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G211gat), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n433), .B(new_n434), .C1(new_n440), .C2(KEYINPUT22), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT22), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT70), .B(G211gat), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n435), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n434), .B1(new_n445), .B2(new_n433), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n312), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n434), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n437), .A2(new_n439), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT22), .B1(new_n452), .B2(G218gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n433), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n451), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n441), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n287), .A2(new_n294), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT29), .B1(new_n457), .B2(new_n300), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G228gat), .A2(G233gat), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n304), .B2(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n450), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n460), .ZN(new_n464));
  INV_X1    g263(.A(new_n311), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n456), .A2(new_n458), .B1(new_n304), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n466), .B2(new_n450), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n463), .A2(new_n467), .A3(G22gat), .ZN(new_n468));
  INV_X1    g267(.A(G22gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n304), .A2(new_n465), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n304), .A2(new_n448), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n447), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT29), .B1(new_n298), .B2(new_n311), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n456), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n460), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n469), .B1(new_n475), .B2(new_n462), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n432), .B1(new_n468), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT80), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT80), .B(new_n432), .C1(new_n468), .C2(new_n476), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n463), .A2(new_n467), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n432), .B1(new_n481), .B2(new_n469), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n476), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(G22gat), .B1(new_n463), .B2(new_n467), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n479), .A2(new_n480), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n415), .A2(new_n414), .A3(new_n418), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT69), .B1(new_n424), .B2(new_n417), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n428), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n413), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n429), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n398), .A2(G226gat), .A3(G233gat), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n398), .A2(new_n448), .B1(G226gat), .B2(G233gat), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n495), .A2(new_n496), .A3(new_n447), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G8gat), .B(G36gat), .Z(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT71), .ZN(new_n500));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n500), .B(new_n501), .Z(new_n502));
  OAI21_X1  g301(.A(new_n447), .B1(new_n495), .B2(new_n496), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n498), .A2(KEYINPUT30), .A3(new_n502), .A4(new_n503), .ZN(new_n507));
  INV_X1    g306(.A(new_n502), .ZN(new_n508));
  INV_X1    g307(.A(new_n503), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(new_n497), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n347), .A2(new_n494), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT35), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT82), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n334), .A2(new_n335), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(new_n340), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT83), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n346), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n332), .A2(KEYINPUT82), .A3(new_n335), .A4(new_n334), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n340), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT35), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n512), .A2(new_n522), .A3(new_n523), .A4(new_n488), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n429), .A2(KEYINPUT84), .A3(new_n493), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n492), .B1(new_n491), .B2(new_n413), .ZN(new_n529));
  AOI211_X1 g328(.A(new_n428), .B(new_n412), .C1(new_n489), .C2(new_n490), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n525), .A2(new_n526), .A3(new_n527), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n527), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT85), .B1(new_n533), .B2(new_n524), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n514), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n529), .A2(new_n530), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT36), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n308), .A2(new_n319), .A3(new_n321), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n310), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT39), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n539), .B(KEYINPUT39), .C1(new_n310), .C2(new_n325), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n266), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT40), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n340), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n544), .B(new_n511), .C1(new_n543), .C2(new_n542), .ZN(new_n545));
  OR3_X1    g344(.A1(new_n509), .A2(KEYINPUT37), .A3(new_n497), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT37), .B1(new_n509), .B2(new_n497), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n508), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT38), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT38), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n546), .A2(new_n550), .A3(new_n508), .A4(new_n547), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n504), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n545), .B(new_n488), .C1(new_n552), .C2(new_n522), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n347), .A2(new_n512), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n537), .B(new_n553), .C1(new_n554), .C2(new_n488), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n257), .B1(new_n535), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  INV_X1    g356(.A(G85gat), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(KEYINPUT8), .A2(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT94), .B(KEYINPUT7), .ZN(new_n561));
  NAND2_X1  g360(.A1(G85gat), .A2(G92gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g362(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n564));
  NAND2_X1  g363(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n564), .A2(new_n565), .B1(G85gat), .B2(G92gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n560), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G99gat), .B(G106gat), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n562), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(G85gat), .A3(G92gat), .A4(new_n565), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n568), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(new_n560), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n233), .A2(new_n230), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT41), .ZN(new_n579));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n572), .A2(new_n573), .A3(new_n560), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n573), .B1(new_n572), .B2(new_n560), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n581), .B1(new_n231), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n577), .A2(KEYINPUT95), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  XOR2_X1   g387(.A(G134gat), .B(G162gat), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n580), .A2(new_n579), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n588), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  XOR2_X1   g392(.A(G71gat), .B(G78gat), .Z(new_n594));
  OR2_X1    g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G57gat), .A2(G64gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT92), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT91), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(KEYINPUT9), .A3(new_n596), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n594), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n594), .A2(new_n603), .A3(new_n602), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n214), .B1(new_n593), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n593), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n607), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT93), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n611), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(KEYINPUT97), .B(KEYINPUT10), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n604), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n594), .A2(new_n603), .A3(new_n602), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n625), .A2(new_n626), .B1(new_n600), .B2(new_n598), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n574), .A2(KEYINPUT96), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n575), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n574), .B(new_n569), .C1(new_n606), .C2(KEYINPUT96), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n601), .B(KEYINPUT10), .C1(new_n604), .C2(new_n605), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT98), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n584), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT98), .B1(new_n575), .B2(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n622), .B1(new_n631), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n629), .A2(new_n630), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n622), .B2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G120gat), .B(G148gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT99), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n640), .A2(new_n644), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n592), .A2(new_n621), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n556), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n347), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n203), .ZN(G1324gat));
  OAI21_X1  g452(.A(G8gat), .B1(new_n651), .B2(new_n512), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT16), .B(G8gat), .Z(new_n656));
  NAND4_X1  g455(.A1(new_n556), .A2(new_n511), .A3(new_n650), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n655), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(KEYINPUT100), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(KEYINPUT100), .ZN(new_n660));
  OAI221_X1 g459(.A(new_n654), .B1(new_n655), .B2(new_n657), .C1(new_n659), .C2(new_n660), .ZN(G1325gat));
  OAI21_X1  g460(.A(G15gat), .B1(new_n651), .B2(new_n537), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n533), .A2(G15gat), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n651), .B2(new_n663), .ZN(G1326gat));
  INV_X1    g463(.A(new_n488), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n556), .A2(new_n665), .A3(new_n650), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n621), .A2(new_n647), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n252), .A2(new_n253), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n535), .A2(new_n555), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n535), .A2(new_n555), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n592), .A2(KEYINPUT44), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n677), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n592), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT44), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n675), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G29gat), .B1(new_n686), .B2(new_n347), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n592), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n556), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n347), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n218), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT45), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n687), .A2(new_n692), .ZN(G1328gat));
  OAI21_X1  g492(.A(G36gat), .B1(new_n686), .B2(new_n512), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n689), .A2(new_n219), .A3(new_n511), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT103), .B(KEYINPUT46), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(G1329gat));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n702));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  INV_X1    g502(.A(new_n537), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n685), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n533), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n556), .A2(new_n703), .A3(new_n706), .A4(new_n688), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n701), .B(new_n702), .C1(new_n705), .C2(new_n709), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n535), .A2(new_n678), .A3(new_n555), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n678), .B1(new_n535), .B2(new_n555), .ZN(new_n712));
  INV_X1    g511(.A(new_n680), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n592), .B1(new_n535), .B2(new_n555), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n704), .B(new_n674), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G43gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n707), .B(KEYINPUT104), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n719), .A2(new_n699), .A3(new_n700), .A4(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n710), .A2(new_n721), .ZN(G1330gat));
  AND2_X1   g521(.A1(new_n665), .A2(G50gat), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n685), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(G50gat), .B1(new_n689), .B2(new_n665), .ZN(new_n725));
  OR3_X1    g524(.A1(new_n724), .A2(KEYINPUT48), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT48), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1331gat));
  NOR2_X1   g527(.A1(new_n711), .A2(new_n712), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n682), .A2(new_n648), .A3(new_n672), .A4(new_n620), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n690), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g533(.A(new_n512), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n731), .A2(KEYINPUT106), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT106), .B1(new_n731), .B2(new_n736), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(G1333gat));
  OR3_X1    g541(.A1(new_n731), .A2(G71gat), .A3(new_n533), .ZN(new_n743));
  OAI21_X1  g542(.A(G71gat), .B1(new_n731), .B2(new_n537), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n743), .A2(KEYINPUT50), .A3(new_n744), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n665), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n673), .A2(new_n620), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT107), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n715), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(new_n558), .A3(new_n690), .A4(new_n647), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n647), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n681), .B2(new_n684), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n759), .A2(new_n690), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n757), .B1(new_n760), .B2(new_n558), .ZN(G1336gat));
  NOR3_X1   g560(.A1(new_n648), .A2(G92gat), .A3(new_n512), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n762), .B(KEYINPUT108), .Z(new_n763));
  AND2_X1   g562(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n559), .B1(new_n759), .B2(new_n511), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n756), .A2(new_n762), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT109), .B(KEYINPUT52), .Z(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n766), .B1(new_n765), .B2(new_n769), .ZN(G1337gat));
  INV_X1    g569(.A(G99gat), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n756), .A2(new_n771), .A3(new_n706), .A4(new_n647), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n759), .A2(new_n704), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n771), .ZN(G1338gat));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n665), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n648), .A2(G106gat), .A3(new_n488), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT110), .Z(new_n778));
  AOI22_X1  g577(.A1(new_n776), .A2(G106gat), .B1(new_n756), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n776), .A2(G106gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n756), .A2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n775), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n775), .A2(new_n779), .B1(new_n780), .B2(new_n782), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n649), .A2(new_n672), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(new_n622), .C1(new_n631), .C2(new_n637), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n788), .A2(new_n789), .A3(new_n644), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n788), .B2(new_n644), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n638), .A2(KEYINPUT54), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n635), .A2(new_n636), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n639), .A2(new_n623), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n797), .B2(new_n622), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n631), .A2(new_n637), .ZN(new_n799));
  INV_X1    g598(.A(new_n622), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(KEYINPUT111), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n793), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n786), .B1(new_n792), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n787), .B1(new_n797), .B2(new_n622), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT111), .B1(new_n799), .B2(new_n800), .ZN(new_n805));
  NOR4_X1   g604(.A1(new_n631), .A2(new_n637), .A3(new_n794), .A4(new_n622), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n807), .B(KEYINPUT55), .C1(new_n790), .C2(new_n791), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(new_n645), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n242), .A2(new_n243), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n235), .B1(new_n234), .B2(new_n237), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n249), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n253), .A3(new_n814), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n809), .A2(new_n592), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n803), .A2(new_n672), .A3(new_n645), .A4(new_n808), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n813), .A2(new_n647), .A3(new_n253), .A4(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n682), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(KEYINPUT114), .A3(new_n818), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n816), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n785), .B1(new_n823), .B2(new_n621), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n347), .A2(new_n511), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n824), .A2(new_n488), .A3(new_n706), .A4(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n826), .A2(new_n277), .A3(new_n257), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n824), .A2(new_n690), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n494), .A2(new_n512), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n672), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n827), .B1(new_n277), .B2(new_n830), .ZN(G1340gat));
  OAI21_X1  g630(.A(G120gat), .B1(new_n826), .B2(new_n648), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n647), .A2(new_n275), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT115), .Z(new_n834));
  NAND3_X1  g633(.A1(new_n828), .A2(new_n829), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT116), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n826), .B2(new_n620), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n828), .A2(new_n829), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n621), .A2(new_n270), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(G1342gat));
  NAND2_X1  g640(.A1(new_n682), .A2(new_n268), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n839), .A2(KEYINPUT56), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n826), .B2(new_n592), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT56), .B1(new_n839), .B2(new_n842), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n847), .A3(new_n665), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n537), .A2(new_n825), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n808), .A2(new_n645), .ZN(new_n850));
  INV_X1    g649(.A(new_n791), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n788), .A2(new_n789), .A3(new_n644), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n853), .B2(new_n807), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT117), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n803), .A2(new_n856), .A3(new_n645), .A4(new_n808), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n855), .A2(new_n256), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n682), .B1(new_n858), .B2(new_n818), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n620), .B1(new_n859), .B2(new_n816), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n488), .B1(new_n860), .B2(new_n785), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n848), .B(new_n849), .C1(new_n847), .C2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n257), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n704), .A2(new_n488), .A3(new_n511), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n257), .A2(G141gat), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n824), .A2(new_n690), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n866), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n866), .A2(new_n871), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n872), .A2(new_n873), .A3(new_n870), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n862), .B2(new_n673), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n869), .A2(new_n870), .B1(new_n874), .B2(new_n875), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n828), .A2(new_n864), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n877), .A2(G148gat), .A3(new_n648), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n819), .A2(new_n820), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(new_n592), .A3(new_n822), .ZN(new_n881));
  INV_X1    g680(.A(new_n816), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n621), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n665), .B1(new_n883), .B2(new_n784), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n650), .A2(new_n257), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n860), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n488), .A2(KEYINPUT57), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n884), .A2(KEYINPUT57), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n648), .B1(new_n849), .B2(KEYINPUT120), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n888), .B(new_n889), .C1(KEYINPUT120), .C2(new_n849), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n879), .B1(new_n890), .B2(G148gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n879), .A2(G148gat), .ZN(new_n892));
  INV_X1    g691(.A(new_n862), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n647), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n878), .B1(new_n891), .B2(new_n894), .ZN(G1345gat));
  OAI21_X1  g694(.A(KEYINPUT121), .B1(new_n877), .B2(new_n620), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n828), .A2(new_n897), .A3(new_n621), .A4(new_n864), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n301), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n621), .A2(new_n301), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT122), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n862), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n899), .A2(new_n902), .ZN(G1346gat));
  OAI21_X1  g702(.A(G162gat), .B1(new_n862), .B2(new_n592), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n682), .A2(new_n289), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n877), .B2(new_n905), .ZN(G1347gat));
  AND2_X1   g705(.A1(new_n824), .A2(new_n488), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n690), .A2(new_n533), .A3(new_n512), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n257), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n494), .A2(new_n511), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT123), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n824), .A2(new_n347), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n388), .A3(new_n672), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT124), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n910), .A2(new_n918), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1348gat));
  OAI21_X1  g719(.A(G176gat), .B1(new_n909), .B2(new_n648), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n914), .A2(new_n373), .A3(new_n647), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n621), .A3(new_n908), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(G183gat), .ZN(new_n925));
  INV_X1    g724(.A(new_n383), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n620), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT125), .B1(new_n914), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NOR4_X1   g728(.A1(new_n913), .A2(new_n929), .A3(new_n926), .A4(new_n620), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n925), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT60), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT60), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n925), .B(new_n933), .C1(new_n928), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n914), .A2(new_n361), .A3(new_n682), .ZN(new_n936));
  OAI21_X1  g735(.A(G190gat), .B1(new_n909), .B2(new_n592), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(G1351gat));
  AND2_X1   g739(.A1(new_n824), .A2(new_n347), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n704), .A2(new_n488), .A3(new_n512), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n672), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n847), .B1(new_n824), .B2(new_n665), .ZN(new_n946));
  INV_X1    g745(.A(new_n887), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n860), .B2(new_n885), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n537), .A2(new_n347), .A3(new_n511), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n256), .A2(G197gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n647), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n648), .A2(G204gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n941), .A2(new_n942), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(KEYINPUT62), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n956), .A2(new_n960), .A3(KEYINPUT62), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n954), .B(new_n957), .C1(new_n959), .C2(new_n961), .ZN(G1353gat));
  NAND3_X1  g761(.A1(new_n944), .A2(new_n444), .A3(new_n621), .ZN(new_n963));
  INV_X1    g762(.A(new_n949), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n888), .A2(new_n621), .A3(new_n964), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  NAND3_X1  g767(.A1(new_n944), .A2(new_n435), .A3(new_n682), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n888), .B2(new_n964), .ZN(new_n971));
  NOR4_X1   g770(.A1(new_n946), .A2(new_n948), .A3(KEYINPUT127), .A4(new_n949), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n971), .A2(new_n972), .A3(new_n592), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n973), .B2(new_n435), .ZN(G1355gat));
endmodule


