//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990;
  INV_X1    g000(.A(KEYINPUT83), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G211gat), .A2(G218gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209));
  AND2_X1   g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n214), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT73), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT73), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n221));
  NAND2_X1  g020(.A1(G226gat), .A2(G233gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT23), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT23), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n225), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n226), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234));
  AND2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(KEYINPUT24), .ZN(new_n236));
  NAND2_X1  g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n237), .A2(KEYINPUT64), .A3(new_n238), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(new_n239), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT25), .B(new_n224), .C1(new_n225), .C2(KEYINPUT23), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n225), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n247), .B1(new_n251), .B2(KEYINPUT23), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n244), .A2(new_n245), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G190gat), .ZN(new_n254));
  AND2_X1   g053(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT28), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n259), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n237), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT26), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n251), .A2(KEYINPUT67), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n224), .B1(new_n225), .B2(new_n262), .ZN(new_n264));
  INV_X1    g063(.A(new_n250), .ZN(new_n265));
  NOR3_X1   g064(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n261), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n223), .B1(new_n253), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n253), .B2(new_n270), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n221), .A2(new_n271), .B1(new_n273), .B2(new_n222), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n236), .A2(new_n241), .A3(new_n242), .ZN(new_n275));
  AND2_X1   g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n227), .A2(new_n228), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT23), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n229), .A2(new_n230), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT65), .B1(new_n225), .B2(KEYINPUT23), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n245), .B1(new_n275), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n252), .A2(new_n246), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n263), .ZN(new_n286));
  INV_X1    g085(.A(new_n261), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(KEYINPUT75), .A3(new_n223), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n220), .B1(new_n274), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT29), .B1(new_n285), .B2(new_n288), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n220), .B(new_n271), .C1(new_n292), .C2(new_n223), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n205), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n222), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n271), .A2(new_n221), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n290), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n219), .ZN(new_n299));
  INV_X1    g098(.A(new_n205), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(new_n293), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(KEYINPUT30), .A3(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n291), .A2(new_n294), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n300), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308));
  INV_X1    g107(.A(G85gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT0), .B(G57gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G141gat), .B(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OR2_X1    g114(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n316));
  INV_X1    g115(.A(G155gat), .ZN(new_n317));
  INV_X1    g116(.A(G162gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(G155gat), .B2(G162gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n315), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n328), .B(new_n316), .C1(new_n314), .C2(new_n323), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331));
  INV_X1    g130(.A(G127gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(G134gat), .ZN(new_n333));
  INV_X1    g132(.A(G134gat), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n333), .B1(G127gat), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(G127gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(new_n331), .ZN(new_n337));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338));
  OAI22_X1  g137(.A1(new_n335), .A2(new_n337), .B1(KEYINPUT1), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(KEYINPUT69), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(G120gat), .ZN(new_n343));
  INV_X1    g142(.A(G120gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n344), .A2(G113gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n341), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT1), .B1(new_n332), .B2(G134gat), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n340), .A2(new_n346), .A3(new_n336), .A4(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n339), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT4), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n339), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n325), .A2(new_n329), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n351), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n325), .A2(new_n329), .A3(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(KEYINPUT3), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT5), .A2(new_n354), .A3(new_n355), .A4(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT5), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n351), .A2(new_n352), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n349), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n355), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n350), .A2(new_n353), .B1(new_n359), .B2(new_n358), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n313), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(new_n360), .ZN(new_n371));
  INV_X1    g170(.A(new_n366), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n367), .A2(KEYINPUT5), .A3(new_n355), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n312), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n369), .A2(new_n370), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT6), .A4(new_n312), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n306), .A2(new_n307), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n351), .B1(new_n253), .B2(new_n270), .ZN(new_n380));
  INV_X1    g179(.A(new_n351), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n285), .A2(new_n288), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G227gat), .ZN(new_n383));
  INV_X1    g182(.A(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n380), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT70), .B(G15gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G43gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  AOI21_X1  g190(.A(new_n386), .B1(new_n380), .B2(new_n382), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n387), .B(new_n391), .C1(new_n392), .C2(KEYINPUT33), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n253), .A2(new_n270), .A3(new_n351), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n381), .B1(new_n285), .B2(new_n288), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  INV_X1    g196(.A(new_n391), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n396), .B(new_n386), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n385), .B1(new_n394), .B2(new_n395), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT34), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(KEYINPUT32), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT34), .B1(new_n392), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n213), .A2(new_n215), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n352), .A2(new_n408), .A3(new_n272), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n359), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT78), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT78), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n412), .A3(new_n359), .ZN(new_n413));
  AND2_X1   g212(.A1(G228gat), .A2(G233gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n357), .A2(new_n272), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n415), .B2(new_n219), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n217), .A2(new_n418), .A3(new_n218), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n330), .B1(new_n419), .B2(new_n356), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n357), .A2(new_n272), .B1(new_n217), .B2(new_n218), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n424), .B(KEYINPUT31), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G22gat), .B(G50gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT79), .ZN(new_n428));
  INV_X1    g227(.A(new_n425), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n417), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n428), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n417), .A2(new_n422), .A3(new_n429), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n417), .B2(new_n422), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n393), .A2(new_n399), .A3(new_n403), .A4(new_n405), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n407), .A2(new_n431), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n435), .A2(new_n431), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(KEYINPUT82), .A3(new_n436), .A4(new_n407), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n307), .B1(new_n306), .B2(new_n378), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n379), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT35), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n202), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n439), .A2(new_n441), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n306), .A2(new_n378), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT77), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n306), .A2(new_n307), .A3(new_n378), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(KEYINPUT83), .A3(KEYINPUT35), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n407), .A2(new_n436), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n445), .A3(new_n440), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(new_n448), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n446), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n367), .A2(new_n355), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT39), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n312), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n364), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n460), .B1(new_n462), .B2(new_n355), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n367), .B2(new_n355), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n461), .A2(KEYINPUT40), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n375), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT40), .B1(new_n461), .B2(new_n464), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n440), .B1(new_n468), .B2(new_n306), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT38), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n300), .B1(new_n303), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n291), .B2(new_n294), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n376), .A2(new_n377), .A3(new_n301), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n296), .A2(new_n297), .A3(new_n290), .A4(new_n220), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n292), .A2(new_n223), .ZN(new_n478));
  INV_X1    g277(.A(new_n271), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n219), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(new_n476), .B2(KEYINPUT80), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT37), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n472), .A2(new_n470), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n475), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n474), .B1(new_n484), .B2(KEYINPUT81), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT81), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n475), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n469), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n440), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n379), .B2(new_n443), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n407), .A2(KEYINPUT36), .A3(new_n436), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(KEYINPUT71), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n453), .B2(new_n495), .ZN(new_n496));
  AOI211_X1 g295(.A(KEYINPUT72), .B(KEYINPUT36), .C1(new_n407), .C2(new_n436), .ZN(new_n497));
  OAI22_X1  g296(.A1(new_n492), .A2(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n488), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n458), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g300(.A1(G29gat), .A2(G36gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n502), .B(KEYINPUT14), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT86), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n502), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT86), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509));
  OR2_X1    g308(.A1(G43gat), .A2(G50gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(G43gat), .A2(G50gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(KEYINPUT85), .B(G50gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n509), .B(new_n511), .C1(new_n517), .C2(G43gat), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n505), .A2(new_n508), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n512), .B1(new_n503), .B2(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n523), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  INV_X1    g325(.A(G92gat), .ZN(new_n527));
  AOI22_X1  g326(.A1(KEYINPUT8), .A2(new_n526), .B1(new_n309), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529));
  OAI22_X1  g328(.A1(new_n309), .A2(new_n527), .B1(new_n529), .B2(KEYINPUT89), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n531), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  XOR2_X1   g332(.A(G99gat), .B(G106gat), .Z(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT90), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n525), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(G134gat), .B(G162gat), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n520), .B2(new_n519), .ZN(new_n542));
  AND2_X1   g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(KEYINPUT41), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n539), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(new_n539), .B2(new_n544), .ZN(new_n546));
  XOR2_X1   g345(.A(G190gat), .B(G218gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT91), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n543), .A2(KEYINPUT41), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  OR3_X1    g350(.A1(new_n545), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n545), .B2(new_n546), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT16), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(G1gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(G1gat), .B2(new_n556), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G8gat), .ZN(new_n560));
  XOR2_X1   g359(.A(G57gat), .B(G64gat), .Z(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n561), .A2(new_n567), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n560), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n571), .B(KEYINPUT21), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(new_n560), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT88), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G183gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(G211gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n576), .B(new_n580), .Z(new_n581));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n581), .A2(new_n584), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n555), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n560), .B1(new_n522), .B2(new_n524), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n560), .A2(new_n521), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT18), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n560), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n525), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n593), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(new_n591), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT18), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(KEYINPUT87), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n560), .B(new_n521), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n591), .B(KEYINPUT13), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n596), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G169gat), .B(G197gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G113gat), .B(G141gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT84), .B(KEYINPUT11), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n596), .A2(new_n602), .A3(new_n613), .A4(new_n606), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n537), .A2(new_n571), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n535), .A2(new_n570), .A3(new_n569), .A4(new_n536), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n621), .A2(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n621), .ZN(new_n627));
  INV_X1    g426(.A(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n626), .A2(new_n629), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT92), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n626), .A2(KEYINPUT92), .A3(new_n629), .A4(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n626), .A2(new_n629), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n632), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n618), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n501), .A2(new_n589), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n378), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G1gat), .ZN(G1324gat));
  INV_X1    g445(.A(new_n306), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G8gat), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT42), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n557), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  MUX2_X1   g452(.A(KEYINPUT42), .B(new_n650), .S(new_n653), .Z(G1325gat));
  AOI21_X1  g453(.A(G15gat), .B1(new_n643), .B2(new_n454), .ZN(new_n655));
  INV_X1    g454(.A(new_n498), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n656), .A2(G15gat), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n643), .B2(new_n657), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n489), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT43), .B(G22gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1327gat));
  NOR2_X1   g460(.A1(new_n488), .A2(new_n499), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n456), .B1(new_n663), .B2(new_n202), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n664), .B2(new_n452), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n585), .A2(new_n586), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n642), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n665), .A2(new_n555), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n513), .A3(new_n644), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT93), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT93), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n668), .A2(new_n671), .A3(new_n513), .A4(new_n644), .ZN(new_n672));
  AND3_X1   g471(.A1(new_n670), .A2(new_n672), .A3(KEYINPUT45), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT45), .B1(new_n670), .B2(new_n672), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n666), .B(KEYINPUT94), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n641), .B(KEYINPUT95), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n617), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT96), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n555), .B1(new_n458), .B2(new_n500), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n680), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OAI211_X1 g482(.A(KEYINPUT96), .B(KEYINPUT44), .C1(new_n665), .C2(new_n555), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT97), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n458), .A2(new_n686), .A3(new_n500), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n458), .B2(new_n500), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n682), .B(new_n554), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n679), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n644), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G29gat), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n690), .B2(new_n644), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n675), .B1(new_n693), .B2(new_n694), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n668), .A2(new_n514), .A3(new_n647), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(KEYINPUT46), .Z(new_n697));
  INV_X1    g496(.A(KEYINPUT99), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n690), .A2(new_n698), .A3(new_n647), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G36gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n690), .B2(new_n647), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n668), .A2(new_n703), .A3(new_n454), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n498), .B(new_n679), .C1(new_n685), .C2(new_n689), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n703), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT47), .B(new_n704), .C1(new_n705), .C2(new_n703), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1330gat));
  INV_X1    g509(.A(new_n517), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n668), .A2(new_n489), .A3(new_n711), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n440), .B(new_n679), .C1(new_n685), .C2(new_n689), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n713), .B2(new_n711), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g515(.A(KEYINPUT48), .B(new_n712), .C1(new_n713), .C2(new_n711), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n588), .A2(new_n617), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n677), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT100), .Z(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n687), .B2(new_n688), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n644), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT101), .B(G57gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1332gat));
  XNOR2_X1  g525(.A(new_n306), .B(KEYINPUT103), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(KEYINPUT102), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n729), .B(new_n721), .C1(new_n687), .C2(new_n688), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n727), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n732));
  AND2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n734), .B1(new_n731), .B2(new_n732), .ZN(G1333gat));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n501), .A2(KEYINPUT97), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n458), .A2(new_n500), .A3(new_n686), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n729), .B1(new_n739), .B2(new_n721), .ZN(new_n740));
  INV_X1    g539(.A(new_n730), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n656), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G71gat), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n723), .A2(new_n563), .A3(new_n454), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n736), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n498), .B1(new_n728), .B2(new_n730), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n744), .B(new_n736), .C1(new_n746), .C2(new_n563), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n745), .A2(new_n748), .ZN(G1334gat));
  AOI21_X1  g548(.A(new_n440), .B1(new_n728), .B2(new_n730), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(new_n564), .ZN(G1335gat));
  NAND3_X1  g550(.A1(new_n618), .A2(new_n666), .A3(new_n641), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n752), .B1(new_n685), .B2(new_n689), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n378), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT104), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n617), .A2(new_n587), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n501), .A2(new_n554), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n756), .A3(KEYINPUT51), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(KEYINPUT51), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n681), .A2(new_n761), .A3(new_n758), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n641), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n644), .A2(new_n309), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n755), .B1(new_n763), .B2(new_n764), .ZN(G1336gat));
  AOI21_X1  g564(.A(new_n527), .B1(new_n753), .B2(new_n647), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n727), .A2(G92gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n760), .A2(new_n677), .A3(new_n762), .A4(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(KEYINPUT52), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n771));
  INV_X1    g570(.A(new_n727), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n527), .B1(new_n753), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n768), .A2(new_n774), .ZN(new_n777));
  AOI211_X1 g576(.A(new_n727), .B(new_n752), .C1(new_n685), .C2(new_n689), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n777), .B(KEYINPUT105), .C1(new_n778), .C2(new_n527), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n770), .A2(new_n776), .A3(new_n779), .ZN(G1337gat));
  NOR2_X1   g579(.A1(new_n754), .A2(new_n498), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT106), .B(G99gat), .Z(new_n782));
  NAND2_X1  g581(.A1(new_n454), .A2(new_n782), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n781), .A2(new_n782), .B1(new_n763), .B2(new_n783), .ZN(G1338gat));
  NOR2_X1   g583(.A1(new_n440), .A2(G106gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n760), .A2(new_n677), .A3(new_n762), .A4(new_n785), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n440), .B(new_n752), .C1(new_n685), .C2(new_n689), .ZN(new_n787));
  INV_X1    g586(.A(G106gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1339gat));
  INV_X1    g592(.A(new_n676), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n591), .B1(new_n598), .B2(new_n599), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n603), .A2(new_n605), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n612), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT108), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(KEYINPUT108), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n641), .A2(new_n798), .A3(new_n616), .A4(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n626), .A2(KEYINPUT54), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n628), .B1(new_n622), .B2(new_n623), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n633), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n804), .B1(new_n803), .B2(new_n807), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n638), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n615), .B2(new_n616), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n801), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n803), .A2(new_n807), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT55), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n814), .A2(new_n815), .B1(new_n636), .B2(new_n637), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n617), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n817), .A2(new_n818), .A3(new_n800), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n812), .A2(new_n555), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n816), .A2(new_n554), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n798), .A2(new_n616), .A3(new_n799), .ZN(new_n822));
  OR3_X1    g621(.A1(new_n821), .A2(KEYINPUT109), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT109), .B1(new_n821), .B2(new_n822), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n794), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n641), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n589), .A2(new_n827), .A3(new_n618), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT107), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n719), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n440), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n826), .A2(new_n832), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT111), .B1(new_n836), .B2(new_n489), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n453), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n644), .A3(new_n727), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n618), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n836), .A2(new_n378), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n447), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n772), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n342), .A3(new_n617), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(G1340gat));
  OAI21_X1  g644(.A(G120gat), .B1(new_n839), .B2(new_n678), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n344), .A3(new_n641), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1341gat));
  NOR3_X1   g647(.A1(new_n839), .A2(new_n332), .A3(new_n676), .ZN(new_n849));
  AOI21_X1  g648(.A(G127gat), .B1(new_n843), .B2(new_n587), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(G1342gat));
  OAI21_X1  g650(.A(G134gat), .B1(new_n839), .B2(new_n555), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n647), .A2(new_n555), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n334), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT56), .B1(new_n842), .B2(new_n854), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n842), .A2(KEYINPUT56), .A3(new_n854), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(G1343gat));
  OAI21_X1  g656(.A(new_n555), .B1(new_n801), .B2(new_n811), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT112), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n554), .B1(new_n817), .B2(new_n800), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n825), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n832), .B1(new_n863), .B2(new_n666), .ZN(new_n864));
  OAI21_X1  g663(.A(KEYINPUT57), .B1(new_n864), .B2(new_n440), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n727), .A2(new_n644), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n656), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n868), .B(new_n489), .C1(new_n826), .C2(new_n832), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G141gat), .B1(new_n870), .B2(new_n618), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n498), .A2(new_n489), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT113), .Z(new_n873));
  AND4_X1   g672(.A1(new_n644), .A2(new_n833), .A3(new_n727), .A4(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(G141gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n874), .A2(new_n875), .A3(new_n617), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n871), .B2(new_n876), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n871), .A2(new_n881), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n879), .A2(new_n880), .B1(new_n882), .B2(KEYINPUT58), .ZN(new_n883));
  INV_X1    g682(.A(new_n880), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT58), .B1(new_n871), .B2(new_n881), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n885), .A3(new_n878), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(G1344gat));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n865), .A2(new_n869), .A3(new_n641), .A4(new_n867), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  INV_X1    g689(.A(G148gat), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n891), .A2(KEYINPUT59), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n836), .B2(new_n440), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n821), .A2(new_n822), .ZN(new_n896));
  OR3_X1    g695(.A1(new_n860), .A2(KEYINPUT118), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT118), .B1(new_n860), .B2(new_n896), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n666), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n828), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n868), .A3(new_n489), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n895), .A2(new_n901), .A3(new_n641), .A4(new_n867), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n894), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n890), .B1(new_n889), .B2(new_n892), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n893), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n841), .A2(new_n727), .A3(new_n873), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n641), .A2(new_n891), .ZN(new_n907));
  OR3_X1    g706(.A1(new_n906), .A2(KEYINPUT116), .A3(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT116), .B1(new_n906), .B2(new_n907), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n888), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n889), .A2(new_n892), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT117), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n902), .A2(G148gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n894), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT119), .B(new_n912), .C1(new_n916), .C2(new_n893), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n917), .ZN(G1345gat));
  NOR3_X1   g717(.A1(new_n870), .A2(new_n317), .A3(new_n676), .ZN(new_n919));
  AOI21_X1  g718(.A(G155gat), .B1(new_n874), .B2(new_n587), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(G1346gat));
  OAI21_X1  g720(.A(G162gat), .B1(new_n870), .B2(new_n555), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n841), .A2(new_n318), .A3(new_n853), .A4(new_n873), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n924), .B(KEYINPUT120), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n644), .A2(new_n306), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n838), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n618), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n836), .A2(new_n644), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n727), .A2(new_n442), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n227), .A3(new_n617), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n933), .ZN(G1348gat));
  OAI21_X1  g733(.A(new_n228), .B1(new_n931), .B2(new_n827), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT121), .Z(new_n936));
  NOR3_X1   g735(.A1(new_n927), .A2(new_n228), .A3(new_n678), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n927), .B2(new_n676), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n932), .B(new_n587), .C1(new_n256), .C2(new_n255), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT60), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n254), .A3(new_n554), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n838), .A2(new_n554), .A3(new_n926), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n947), .A2(new_n948), .A3(G190gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n947), .B2(G190gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(G1351gat));
  NOR2_X1   g750(.A1(new_n872), .A2(new_n727), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n929), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n618), .A2(G197gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n895), .A2(new_n901), .A3(new_n498), .A4(new_n926), .ZN(new_n958));
  OAI21_X1  g757(.A(G197gat), .B1(new_n958), .B2(new_n618), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT123), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT123), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1352gat));
  OR2_X1    g763(.A1(new_n958), .A2(new_n678), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n827), .A2(G204gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n929), .A2(new_n952), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  OR3_X1    g768(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT62), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n968), .B2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(KEYINPUT62), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n966), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT125), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n966), .A2(new_n973), .A3(new_n976), .A4(new_n970), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n975), .A2(new_n977), .ZN(G1353gat));
  OR3_X1    g777(.A1(new_n953), .A2(G211gat), .A3(new_n666), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n958), .A2(new_n666), .ZN(new_n980));
  AND3_X1   g779(.A1(new_n980), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n981));
  AOI21_X1  g780(.A(KEYINPUT63), .B1(new_n980), .B2(G211gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  INV_X1    g782(.A(G218gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n984), .B1(new_n953), .B2(new_n555), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987));
  OAI211_X1 g786(.A(new_n987), .B(new_n984), .C1(new_n953), .C2(new_n555), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n554), .A2(G218gat), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n986), .B(new_n988), .C1(new_n958), .C2(new_n989), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


