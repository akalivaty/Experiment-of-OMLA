

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U325 ( .A(n424), .B(n309), .Z(n525) );
  XNOR2_X1 U326 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U327 ( .A(n351), .B(n350), .ZN(n354) );
  XNOR2_X1 U328 ( .A(n363), .B(KEYINPUT65), .ZN(n364) );
  XNOR2_X1 U329 ( .A(n573), .B(n364), .ZN(n452) );
  XNOR2_X1 U330 ( .A(n457), .B(G190GAT), .ZN(n458) );
  XNOR2_X1 U331 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT86), .B(KEYINPUT17), .Z(n294) );
  XNOR2_X1 U333 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U335 ( .A(G169GAT), .B(n295), .ZN(n424) );
  XOR2_X1 U336 ( .A(G15GAT), .B(G127GAT), .Z(n386) );
  XOR2_X1 U337 ( .A(G120GAT), .B(KEYINPUT0), .Z(n297) );
  XNOR2_X1 U338 ( .A(G113GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n297), .B(n296), .ZN(n445) );
  XOR2_X1 U340 ( .A(n386), .B(n445), .Z(n299) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U342 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U343 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n301) );
  NAND2_X1 U344 ( .A1(G227GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U346 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U347 ( .A(G183GAT), .B(KEYINPUT85), .Z(n305) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G71GAT), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n306), .B(G176GAT), .ZN(n307) );
  XNOR2_X1 U351 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U352 ( .A(G211GAT), .B(KEYINPUT22), .Z(n311) );
  XNOR2_X1 U353 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n324) );
  XOR2_X1 U355 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n313) );
  NAND2_X1 U356 ( .A1(G228GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U358 ( .A(n314), .B(G204GAT), .Z(n318) );
  XNOR2_X1 U359 ( .A(G22GAT), .B(G155GAT), .ZN(n315) );
  XNOR2_X1 U360 ( .A(n315), .B(G78GAT), .ZN(n395) );
  XNOR2_X1 U361 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n316), .B(KEYINPUT2), .ZN(n444) );
  XNOR2_X1 U363 ( .A(n395), .B(n444), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n318), .B(n317), .ZN(n320) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n319), .B(G148GAT), .ZN(n358) );
  XOR2_X1 U367 ( .A(n320), .B(n358), .Z(n322) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n335) );
  XOR2_X1 U369 ( .A(G197GAT), .B(KEYINPUT21), .Z(n415) );
  XNOR2_X1 U370 ( .A(n335), .B(n415), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n466) );
  XOR2_X1 U373 ( .A(KEYINPUT78), .B(G92GAT), .Z(n326) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(KEYINPUT80), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n343) );
  XOR2_X1 U376 ( .A(KEYINPUT9), .B(KEYINPUT79), .Z(n328) );
  NAND2_X1 U377 ( .A1(G232GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U379 ( .A(n329), .B(KEYINPUT11), .Z(n334) );
  XOR2_X1 U380 ( .A(G29GAT), .B(G43GAT), .Z(n331) );
  XNOR2_X1 U381 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n331), .B(n330), .ZN(n367) );
  XNOR2_X1 U383 ( .A(G36GAT), .B(G190GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n332), .B(G218GAT), .ZN(n421) );
  XNOR2_X1 U385 ( .A(n367), .B(n421), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U387 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n337) );
  XOR2_X1 U388 ( .A(G99GAT), .B(G85GAT), .Z(n349) );
  XNOR2_X1 U389 ( .A(n335), .B(n349), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n341) );
  XNOR2_X1 U392 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U394 ( .A(n343), .B(n342), .Z(n542) );
  INV_X1 U395 ( .A(n542), .ZN(n557) );
  XOR2_X1 U396 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n345) );
  XNOR2_X1 U397 ( .A(KEYINPUT76), .B(KEYINPUT75), .ZN(n344) );
  XOR2_X1 U398 ( .A(n345), .B(n344), .Z(n362) );
  XOR2_X1 U399 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n347) );
  XNOR2_X1 U400 ( .A(G120GAT), .B(G78GAT), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n351) );
  NAND2_X1 U402 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XOR2_X1 U403 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n353) );
  XNOR2_X1 U404 ( .A(G71GAT), .B(G57GAT), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n399) );
  XNOR2_X1 U406 ( .A(n354), .B(n399), .ZN(n360) );
  XOR2_X1 U407 ( .A(G64GAT), .B(KEYINPUT77), .Z(n356) );
  XNOR2_X1 U408 ( .A(G204GAT), .B(G92GAT), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U410 ( .A(G176GAT), .B(n357), .Z(n420) );
  XNOR2_X1 U411 ( .A(n358), .B(n420), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U413 ( .A(n362), .B(n361), .ZN(n573) );
  INV_X1 U414 ( .A(KEYINPUT41), .ZN(n363) );
  XOR2_X1 U415 ( .A(G141GAT), .B(G197GAT), .Z(n366) );
  XNOR2_X1 U416 ( .A(G169GAT), .B(G22GAT), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n366), .B(n365), .ZN(n380) );
  XOR2_X1 U418 ( .A(KEYINPUT71), .B(G1GAT), .Z(n387) );
  XOR2_X1 U419 ( .A(n387), .B(n367), .Z(n369) );
  XNOR2_X1 U420 ( .A(G50GAT), .B(G36GAT), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U422 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n371) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U425 ( .A(n373), .B(n372), .Z(n378) );
  XOR2_X1 U426 ( .A(KEYINPUT29), .B(G8GAT), .Z(n375) );
  XNOR2_X1 U427 ( .A(G113GAT), .B(G15GAT), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n376), .B(KEYINPUT30), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U431 ( .A(n380), .B(n379), .Z(n545) );
  OR2_X1 U432 ( .A1(n452), .A2(n545), .ZN(n382) );
  XOR2_X1 U433 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n381) );
  XNOR2_X1 U434 ( .A(n382), .B(n381), .ZN(n383) );
  NOR2_X1 U435 ( .A1(n557), .A2(n383), .ZN(n402) );
  XOR2_X1 U436 ( .A(KEYINPUT84), .B(KEYINPUT81), .Z(n385) );
  XNOR2_X1 U437 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n391) );
  XOR2_X1 U439 ( .A(KEYINPUT82), .B(G64GAT), .Z(n389) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U441 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U442 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U443 ( .A1(G231GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U445 ( .A(n394), .B(KEYINPUT14), .Z(n397) );
  XNOR2_X1 U446 ( .A(n395), .B(KEYINPUT83), .ZN(n396) );
  XNOR2_X1 U447 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U448 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U449 ( .A(G8GAT), .B(G183GAT), .Z(n400) );
  XOR2_X1 U450 ( .A(G211GAT), .B(n400), .Z(n418) );
  XNOR2_X1 U451 ( .A(n401), .B(n418), .ZN(n405) );
  XOR2_X1 U452 ( .A(KEYINPUT111), .B(n405), .Z(n564) );
  NAND2_X1 U453 ( .A1(n402), .A2(n564), .ZN(n403) );
  XNOR2_X1 U454 ( .A(n403), .B(KEYINPUT47), .ZN(n404) );
  XNOR2_X1 U455 ( .A(n404), .B(KEYINPUT113), .ZN(n411) );
  INV_X1 U456 ( .A(n405), .ZN(n576) );
  INV_X1 U457 ( .A(n576), .ZN(n490) );
  XNOR2_X1 U458 ( .A(KEYINPUT36), .B(KEYINPUT101), .ZN(n406) );
  XOR2_X1 U459 ( .A(n406), .B(n542), .Z(n579) );
  NOR2_X1 U460 ( .A1(n490), .A2(n579), .ZN(n407) );
  XOR2_X1 U461 ( .A(KEYINPUT45), .B(n407), .Z(n408) );
  NOR2_X1 U462 ( .A1(n573), .A2(n408), .ZN(n409) );
  NAND2_X1 U463 ( .A1(n409), .A2(n545), .ZN(n410) );
  NAND2_X1 U464 ( .A1(n411), .A2(n410), .ZN(n414) );
  XOR2_X1 U465 ( .A(KEYINPUT64), .B(KEYINPUT114), .Z(n412) );
  XNOR2_X1 U466 ( .A(KEYINPUT48), .B(n412), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n414), .B(n413), .ZN(n546) );
  XOR2_X1 U468 ( .A(KEYINPUT92), .B(n415), .Z(n417) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U471 ( .A(n419), .B(n418), .Z(n423) );
  XNOR2_X1 U472 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U473 ( .A(n423), .B(n422), .ZN(n426) );
  INV_X1 U474 ( .A(n424), .ZN(n425) );
  XOR2_X1 U475 ( .A(n426), .B(n425), .Z(n523) );
  XNOR2_X1 U476 ( .A(n523), .B(KEYINPUT120), .ZN(n427) );
  NOR2_X1 U477 ( .A1(n546), .A2(n427), .ZN(n428) );
  XNOR2_X1 U478 ( .A(n428), .B(KEYINPUT54), .ZN(n448) );
  XOR2_X1 U479 ( .A(G85GAT), .B(G162GAT), .Z(n430) );
  XNOR2_X1 U480 ( .A(G29GAT), .B(G155GAT), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U482 ( .A(G57GAT), .B(G148GAT), .Z(n432) );
  XNOR2_X1 U483 ( .A(G1GAT), .B(G127GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U485 ( .A(n434), .B(n433), .Z(n439) );
  XOR2_X1 U486 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n436) );
  NAND2_X1 U487 ( .A1(G225GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U489 ( .A(KEYINPUT6), .B(n437), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U491 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n441) );
  XNOR2_X1 U492 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U496 ( .A(n447), .B(n446), .Z(n473) );
  INV_X1 U497 ( .A(n473), .ZN(n521) );
  NAND2_X1 U498 ( .A1(n448), .A2(n521), .ZN(n567) );
  NOR2_X1 U499 ( .A1(n466), .A2(n567), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n449), .B(KEYINPUT55), .ZN(n450) );
  NOR2_X1 U501 ( .A1(n525), .A2(n450), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n451), .B(KEYINPUT121), .ZN(n563) );
  INV_X1 U503 ( .A(n563), .ZN(n561) );
  INV_X1 U504 ( .A(n452), .ZN(n552) );
  NAND2_X1 U505 ( .A1(n561), .A2(n552), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n454) );
  XNOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n453) );
  XNOR2_X1 U508 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(G1349GAT) );
  NAND2_X1 U510 ( .A1(n561), .A2(n557), .ZN(n459) );
  XOR2_X1 U511 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n457) );
  NOR2_X1 U512 ( .A1(n545), .A2(n573), .ZN(n495) );
  INV_X1 U513 ( .A(n525), .ZN(n533) );
  XNOR2_X1 U514 ( .A(n523), .B(KEYINPUT27), .ZN(n470) );
  NOR2_X1 U515 ( .A1(n521), .A2(n470), .ZN(n548) );
  XOR2_X1 U516 ( .A(KEYINPUT28), .B(KEYINPUT68), .Z(n460) );
  XNOR2_X1 U517 ( .A(n466), .B(n460), .ZN(n528) );
  NAND2_X1 U518 ( .A1(n548), .A2(n528), .ZN(n531) );
  XOR2_X1 U519 ( .A(KEYINPUT93), .B(n531), .Z(n461) );
  NOR2_X1 U520 ( .A1(n533), .A2(n461), .ZN(n476) );
  XNOR2_X1 U521 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT96), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n523), .A2(n525), .ZN(n463) );
  NOR2_X1 U524 ( .A1(n466), .A2(n463), .ZN(n464) );
  XNOR2_X1 U525 ( .A(n465), .B(n464), .ZN(n472) );
  XOR2_X1 U526 ( .A(KEYINPUT95), .B(KEYINPUT26), .Z(n468) );
  NAND2_X1 U527 ( .A1(n466), .A2(n525), .ZN(n467) );
  XNOR2_X1 U528 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U529 ( .A(KEYINPUT94), .B(n469), .ZN(n566) );
  NOR2_X1 U530 ( .A1(n566), .A2(n470), .ZN(n471) );
  NOR2_X1 U531 ( .A1(n472), .A2(n471), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n489) );
  NOR2_X1 U534 ( .A1(n490), .A2(n557), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U536 ( .A1(n489), .A2(n478), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT98), .B(n479), .ZN(n507) );
  NAND2_X1 U538 ( .A1(n495), .A2(n507), .ZN(n487) );
  NOR2_X1 U539 ( .A1(n521), .A2(n487), .ZN(n481) );
  XNOR2_X1 U540 ( .A(KEYINPUT34), .B(KEYINPUT99), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n523), .A2(n487), .ZN(n483) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n483), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n525), .A2(n487), .ZN(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n486), .ZN(G1326GAT) );
  NOR2_X1 U549 ( .A1(n528), .A2(n487), .ZN(n488) );
  XOR2_X1 U550 ( .A(G22GAT), .B(n488), .Z(G1327GAT) );
  NOR2_X1 U551 ( .A1(n489), .A2(n579), .ZN(n491) );
  NAND2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT103), .B(KEYINPUT37), .Z(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(n492), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n519) );
  NAND2_X1 U556 ( .A1(n519), .A2(n495), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(KEYINPUT38), .ZN(n503) );
  NOR2_X1 U558 ( .A1(n503), .A2(n521), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(n498), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n523), .A2(n503), .ZN(n499) );
  XOR2_X1 U562 ( .A(KEYINPUT104), .B(n499), .Z(n500) );
  XNOR2_X1 U563 ( .A(G36GAT), .B(n500), .ZN(G1329GAT) );
  NOR2_X1 U564 ( .A1(n503), .A2(n525), .ZN(n501) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(n501), .Z(n502) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n502), .ZN(G1330GAT) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n505) );
  NOR2_X1 U568 ( .A1(n528), .A2(n503), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  NAND2_X1 U570 ( .A1(n552), .A2(n545), .ZN(n506) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT107), .ZN(n520) );
  NAND2_X1 U572 ( .A1(n520), .A2(n507), .ZN(n515) );
  NOR2_X1 U573 ( .A1(n521), .A2(n515), .ZN(n511) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n509) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT108), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U578 ( .A1(n523), .A2(n515), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NOR2_X1 U581 ( .A1(n525), .A2(n515), .ZN(n514) );
  XOR2_X1 U582 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U583 ( .A1(n528), .A2(n515), .ZN(n517) );
  XNOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U586 ( .A(G78GAT), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n527) );
  NOR2_X1 U588 ( .A1(n521), .A2(n527), .ZN(n522) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U591 ( .A(G92GAT), .B(n524), .Z(G1337GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n527), .ZN(n526) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n546), .A2(n531), .ZN(n532) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n541) );
  NOR2_X1 U599 ( .A1(n545), .A2(n541), .ZN(n534) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n534), .Z(G1340GAT) );
  NOR2_X1 U601 ( .A1(n452), .A2(n541), .ZN(n536) );
  XNOR2_X1 U602 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  NOR2_X1 U605 ( .A1(n564), .A2(n541), .ZN(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  INV_X1 U612 ( .A(n545), .ZN(n569) );
  NOR2_X1 U613 ( .A1(n546), .A2(n566), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(KEYINPUT117), .B(n549), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n569), .A2(n558), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n550), .B(KEYINPUT118), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U620 ( .A1(n558), .A2(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n576), .A2(n558), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT119), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n569), .A2(n561), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(n568), .Z(n580) );
  INV_X1 U635 ( .A(n580), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n577), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(n577), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n585) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(KEYINPUT125), .B(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1355GAT) );
endmodule

