

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733;

  NAND2_X1 U363 ( .A1(n429), .A2(n612), .ZN(n426) );
  NAND2_X1 U364 ( .A1(n714), .A2(n438), .ZN(n437) );
  NOR2_X1 U365 ( .A1(n590), .A2(n440), .ZN(n587) );
  XNOR2_X1 U366 ( .A(n432), .B(KEYINPUT33), .ZN(n677) );
  AND2_X1 U367 ( .A1(n586), .A2(n646), .ZN(n402) );
  XNOR2_X1 U368 ( .A(n564), .B(KEYINPUT1), .ZN(n643) );
  XNOR2_X1 U369 ( .A(n487), .B(n475), .ZN(n692) );
  INV_X1 U370 ( .A(KEYINPUT3), .ZN(n396) );
  INV_X1 U371 ( .A(G953), .ZN(n722) );
  NAND2_X2 U372 ( .A1(n579), .A2(n580), .ZN(n385) );
  XNOR2_X2 U373 ( .A(n372), .B(n469), .ZN(n719) );
  XNOR2_X1 U374 ( .A(G119), .B(G128), .ZN(n479) );
  INV_X1 U375 ( .A(n599), .ZN(n650) );
  NOR2_X1 U376 ( .A1(n650), .A2(n588), .ZN(n624) );
  XNOR2_X2 U377 ( .A(n385), .B(KEYINPUT0), .ZN(n600) );
  XNOR2_X2 U378 ( .A(n518), .B(n466), .ZN(n372) );
  XNOR2_X1 U379 ( .A(n650), .B(n566), .ZN(n589) );
  NAND2_X1 U380 ( .A1(n364), .A2(n363), .ZN(n568) );
  NOR2_X1 U381 ( .A1(n590), .A2(n589), .ZN(n595) );
  XNOR2_X1 U382 ( .A(n402), .B(n401), .ZN(n590) );
  XNOR2_X1 U383 ( .A(n371), .B(KEYINPUT41), .ZN(n676) );
  XNOR2_X1 U384 ( .A(n436), .B(n433), .ZN(n591) );
  XNOR2_X1 U385 ( .A(n445), .B(n444), .ZN(n538) );
  XNOR2_X1 U386 ( .A(n506), .B(n505), .ZN(n707) );
  XNOR2_X1 U387 ( .A(G107), .B(G110), .ZN(n453) );
  XNOR2_X1 U388 ( .A(n452), .B(n451), .ZN(n392) );
  INV_X1 U389 ( .A(n538), .ZN(n558) );
  NOR2_X1 U390 ( .A1(n567), .A2(n416), .ZN(n413) );
  NAND2_X1 U391 ( .A1(n415), .A2(n362), .ZN(n410) );
  NAND2_X1 U392 ( .A1(n567), .A2(n416), .ZN(n415) );
  NAND2_X1 U393 ( .A1(n568), .A2(n416), .ZN(n362) );
  NAND2_X1 U394 ( .A1(n343), .A2(n380), .ZN(n611) );
  XNOR2_X1 U395 ( .A(G131), .B(KEYINPUT66), .ZN(n467) );
  XOR2_X1 U396 ( .A(G134), .B(G137), .Z(n468) );
  INV_X1 U397 ( .A(n568), .ZN(n414) );
  NAND2_X1 U398 ( .A1(n591), .A2(n359), .ZN(n565) );
  NOR2_X1 U399 ( .A1(n585), .A2(n360), .ZN(n359) );
  INV_X1 U400 ( .A(n543), .ZN(n360) );
  NOR2_X1 U401 ( .A1(n616), .A2(G902), .ZN(n493) );
  NAND2_X1 U402 ( .A1(n659), .A2(n559), .ZN(n371) );
  NAND2_X1 U403 ( .A1(n417), .A2(n420), .ZN(n419) );
  AND2_X1 U404 ( .A1(n424), .A2(n422), .ZN(n420) );
  XNOR2_X1 U405 ( .A(n553), .B(KEYINPUT69), .ZN(n363) );
  XNOR2_X1 U406 ( .A(n370), .B(n563), .ZN(n364) );
  NOR2_X1 U407 ( .A1(n614), .A2(n412), .ZN(n411) );
  INV_X1 U408 ( .A(n642), .ZN(n412) );
  OR2_X1 U409 ( .A1(n612), .A2(n641), .ZN(n613) );
  XNOR2_X1 U410 ( .A(n492), .B(n491), .ZN(n506) );
  XNOR2_X1 U411 ( .A(G116), .B(G119), .ZN(n491) );
  INV_X1 U412 ( .A(KEYINPUT4), .ZN(n466) );
  XOR2_X1 U413 ( .A(G146), .B(G125), .Z(n507) );
  AND2_X1 U414 ( .A1(n411), .A2(n413), .ZN(n408) );
  NAND2_X1 U415 ( .A1(n410), .A2(n411), .ZN(n409) );
  NOR2_X1 U416 ( .A1(n605), .A2(n425), .ZN(n424) );
  NAND2_X2 U417 ( .A1(n377), .A2(n373), .ZN(n564) );
  AND2_X1 U418 ( .A1(n379), .A2(n378), .ZN(n377) );
  NAND2_X1 U419 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U420 ( .A(KEYINPUT6), .ZN(n566) );
  AND2_X1 U421 ( .A1(n404), .A2(n348), .ZN(n721) );
  NAND2_X1 U422 ( .A1(n406), .A2(n405), .ZN(n404) );
  INV_X1 U423 ( .A(n641), .ZN(n391) );
  NAND2_X1 U424 ( .A1(n392), .A2(n342), .ZN(n450) );
  XNOR2_X1 U425 ( .A(n481), .B(n341), .ZN(n384) );
  XNOR2_X1 U426 ( .A(n361), .B(KEYINPUT90), .ZN(n481) );
  INV_X1 U427 ( .A(KEYINPUT23), .ZN(n361) );
  XNOR2_X1 U428 ( .A(G113), .B(G143), .ZN(n528) );
  XNOR2_X1 U429 ( .A(n525), .B(n347), .ZN(n403) );
  XNOR2_X1 U430 ( .A(n507), .B(n357), .ZN(n720) );
  XNOR2_X1 U431 ( .A(KEYINPUT10), .B(G140), .ZN(n357) );
  XNOR2_X1 U432 ( .A(G101), .B(G104), .ZN(n470) );
  XOR2_X1 U433 ( .A(KEYINPUT75), .B(G140), .Z(n471) );
  OR2_X1 U434 ( .A1(n424), .A2(n422), .ZN(n421) );
  NOR2_X1 U435 ( .A1(n677), .A2(n603), .ZN(n582) );
  NAND2_X1 U436 ( .A1(n389), .A2(n543), .ZN(n503) );
  XNOR2_X1 U437 ( .A(n496), .B(n390), .ZN(n389) );
  INV_X1 U438 ( .A(KEYINPUT30), .ZN(n390) );
  XNOR2_X1 U439 ( .A(n486), .B(n434), .ZN(n433) );
  NOR2_X1 U440 ( .A1(n704), .A2(G902), .ZN(n436) );
  XNOR2_X1 U441 ( .A(n484), .B(n435), .ZN(n434) );
  INV_X1 U442 ( .A(KEYINPUT22), .ZN(n401) );
  INV_X1 U443 ( .A(n594), .ZN(n440) );
  XNOR2_X1 U444 ( .A(n537), .B(n536), .ZN(n557) );
  INV_X1 U445 ( .A(G475), .ZN(n534) );
  NAND2_X1 U446 ( .A1(n696), .A2(G472), .ZN(n457) );
  NOR2_X1 U447 ( .A1(G952), .A2(n722), .ZN(n706) );
  XNOR2_X1 U448 ( .A(n639), .B(KEYINPUT82), .ZN(n567) );
  INV_X1 U449 ( .A(KEYINPUT48), .ZN(n416) );
  XNOR2_X1 U450 ( .A(n396), .B(G101), .ZN(n489) );
  INV_X1 U451 ( .A(G902), .ZN(n375) );
  INV_X1 U452 ( .A(G469), .ZN(n376) );
  NAND2_X1 U453 ( .A1(G902), .A2(G469), .ZN(n378) );
  INV_X1 U454 ( .A(n410), .ZN(n406) );
  NAND2_X1 U455 ( .A1(n414), .A2(n413), .ZN(n405) );
  INV_X1 U456 ( .A(KEYINPUT84), .ZN(n451) );
  XNOR2_X1 U457 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n447) );
  XNOR2_X1 U458 ( .A(n556), .B(n395), .ZN(n659) );
  INV_X1 U459 ( .A(KEYINPUT110), .ZN(n395) );
  INV_X1 U460 ( .A(KEYINPUT71), .ZN(n382) );
  NOR2_X1 U461 ( .A1(G237), .A2(G902), .ZN(n494) );
  INV_X1 U462 ( .A(KEYINPUT93), .ZN(n435) );
  NOR2_X1 U463 ( .A1(n585), .A2(n591), .ZN(n644) );
  XNOR2_X1 U464 ( .A(n487), .B(n365), .ZN(n616) );
  XNOR2_X1 U465 ( .A(n506), .B(n366), .ZN(n365) );
  XNOR2_X1 U466 ( .A(n346), .B(n461), .ZN(n366) );
  XNOR2_X1 U467 ( .A(n448), .B(n446), .ZN(n520) );
  XNOR2_X1 U468 ( .A(n517), .B(n447), .ZN(n446) );
  XNOR2_X1 U469 ( .A(n516), .B(n515), .ZN(n448) );
  XNOR2_X1 U470 ( .A(G107), .B(G122), .ZN(n517) );
  XNOR2_X1 U471 ( .A(G902), .B(KEYINPUT15), .ZN(n464) );
  XNOR2_X1 U472 ( .A(n707), .B(n458), .ZN(n687) );
  XNOR2_X1 U473 ( .A(n510), .B(n460), .ZN(n459) );
  INV_X1 U474 ( .A(n507), .ZN(n460) );
  NAND2_X1 U475 ( .A1(n408), .A2(n414), .ZN(n407) );
  NAND2_X1 U476 ( .A1(n421), .A2(n634), .ZN(n394) );
  XNOR2_X1 U477 ( .A(n368), .B(n367), .ZN(n569) );
  INV_X1 U478 ( .A(KEYINPUT107), .ZN(n367) );
  NOR2_X1 U479 ( .A1(n631), .A2(n565), .ZN(n369) );
  XNOR2_X1 U480 ( .A(KEYINPUT104), .B(G478), .ZN(n444) );
  OR2_X1 U481 ( .A1(n701), .A2(G902), .ZN(n445) );
  XNOR2_X1 U482 ( .A(n356), .B(n355), .ZN(n704) );
  XNOR2_X1 U483 ( .A(n384), .B(n482), .ZN(n355) );
  XNOR2_X1 U484 ( .A(n358), .B(n720), .ZN(n356) );
  XNOR2_X1 U485 ( .A(n533), .B(n532), .ZN(n698) );
  XNOR2_X1 U486 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U487 ( .A(n720), .B(n403), .ZN(n533) );
  XNOR2_X1 U488 ( .A(n453), .B(n472), .ZN(n474) );
  XNOR2_X1 U489 ( .A(n562), .B(n561), .ZN(n733) );
  NOR2_X1 U490 ( .A1(n554), .A2(n539), .ZN(n641) );
  XNOR2_X1 U491 ( .A(n555), .B(n388), .ZN(n731) );
  INV_X1 U492 ( .A(KEYINPUT40), .ZN(n388) );
  AND2_X1 U493 ( .A1(n418), .A2(n419), .ZN(n555) );
  NOR2_X1 U494 ( .A1(n394), .A2(n393), .ZN(n418) );
  AND2_X1 U495 ( .A1(n441), .A2(n440), .ZN(n639) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n441) );
  INV_X1 U497 ( .A(KEYINPUT36), .ZN(n442) );
  OR2_X1 U498 ( .A1(n569), .A2(n449), .ZN(n443) );
  INV_X1 U499 ( .A(KEYINPUT35), .ZN(n381) );
  XNOR2_X1 U500 ( .A(n399), .B(n397), .ZN(n730) );
  XNOR2_X1 U501 ( .A(n593), .B(KEYINPUT32), .ZN(n397) );
  INV_X1 U502 ( .A(KEYINPUT77), .ZN(n593) );
  INV_X1 U503 ( .A(n706), .ZN(n455) );
  XNOR2_X1 U504 ( .A(n457), .B(n351), .ZN(n456) );
  XOR2_X1 U505 ( .A(KEYINPUT74), .B(KEYINPUT24), .Z(n341) );
  OR2_X1 U506 ( .A1(n611), .A2(KEYINPUT44), .ZN(n342) );
  AND2_X1 U507 ( .A1(n730), .A2(n430), .ZN(n343) );
  NOR2_X1 U508 ( .A1(n538), .A2(n557), .ZN(n634) );
  AND2_X1 U509 ( .A1(n511), .A2(G210), .ZN(n344) );
  AND2_X1 U510 ( .A1(n423), .A2(n421), .ZN(n345) );
  XOR2_X1 U511 ( .A(n488), .B(KEYINPUT94), .Z(n346) );
  AND2_X1 U512 ( .A1(G214), .A2(n526), .ZN(n347) );
  AND2_X1 U513 ( .A1(n642), .A2(n391), .ZN(n348) );
  AND2_X1 U514 ( .A1(n540), .A2(n663), .ZN(n349) );
  XOR2_X1 U515 ( .A(KEYINPUT68), .B(KEYINPUT39), .Z(n350) );
  XOR2_X1 U516 ( .A(n617), .B(KEYINPUT62), .Z(n351) );
  XNOR2_X1 U517 ( .A(n687), .B(n462), .ZN(n352) );
  XNOR2_X1 U518 ( .A(n698), .B(n697), .ZN(n353) );
  XOR2_X1 U519 ( .A(KEYINPUT45), .B(KEYINPUT79), .Z(n354) );
  NAND2_X1 U520 ( .A1(n611), .A2(KEYINPUT44), .ZN(n610) );
  NAND2_X1 U521 ( .A1(n514), .A2(G221), .ZN(n358) );
  NOR2_X1 U522 ( .A1(n599), .A2(n565), .ZN(n544) );
  XNOR2_X2 U523 ( .A(n719), .B(G146), .ZN(n487) );
  INV_X1 U524 ( .A(n589), .ZN(n581) );
  NAND2_X1 U525 ( .A1(n589), .A2(n369), .ZN(n368) );
  INV_X1 U526 ( .A(n549), .ZN(n572) );
  XNOR2_X2 U527 ( .A(n512), .B(n344), .ZN(n549) );
  NAND2_X1 U528 ( .A1(n549), .A2(n349), .ZN(n541) );
  NAND2_X1 U529 ( .A1(n733), .A2(n731), .ZN(n370) );
  NAND2_X1 U530 ( .A1(n560), .A2(n676), .ZN(n561) );
  XNOR2_X1 U531 ( .A(n459), .B(n372), .ZN(n458) );
  NAND2_X1 U532 ( .A1(n692), .A2(G469), .ZN(n379) );
  OR2_X1 U533 ( .A1(n692), .A2(n374), .ZN(n373) );
  XNOR2_X1 U534 ( .A(n380), .B(G122), .ZN(G24) );
  XNOR2_X2 U535 ( .A(n431), .B(n381), .ZN(n380) );
  NAND2_X1 U536 ( .A1(n696), .A2(G210), .ZN(n387) );
  AND2_X4 U537 ( .A1(n427), .A2(n426), .ZN(n696) );
  XNOR2_X1 U538 ( .A(n387), .B(n352), .ZN(n688) );
  XNOR2_X2 U539 ( .A(n450), .B(n354), .ZN(n714) );
  NOR2_X2 U540 ( .A1(n598), .A2(n581), .ZN(n432) );
  XNOR2_X2 U541 ( .A(n383), .B(n382), .ZN(n598) );
  NAND2_X1 U542 ( .A1(n643), .A2(n644), .ZN(n383) );
  NAND2_X1 U543 ( .A1(n456), .A2(n455), .ZN(n454) );
  XNOR2_X1 U544 ( .A(n386), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U545 ( .A1(n699), .A2(n706), .ZN(n386) );
  XNOR2_X2 U546 ( .A(n493), .B(G472), .ZN(n599) );
  XNOR2_X1 U547 ( .A(n400), .B(n353), .ZN(n699) );
  NAND2_X1 U548 ( .A1(n409), .A2(n407), .ZN(n439) );
  INV_X1 U549 ( .A(n423), .ZN(n393) );
  NAND2_X1 U550 ( .A1(n714), .A2(n721), .ZN(n429) );
  INV_X1 U551 ( .A(n662), .ZN(n425) );
  XNOR2_X1 U552 ( .A(n453), .B(KEYINPUT16), .ZN(n504) );
  INV_X1 U553 ( .A(n624), .ZN(n430) );
  NAND2_X1 U554 ( .A1(n549), .A2(n663), .ZN(n449) );
  XNOR2_X1 U555 ( .A(n398), .B(n689), .ZN(G51) );
  NOR2_X2 U556 ( .A1(n688), .A2(n706), .ZN(n398) );
  NAND2_X1 U557 ( .A1(n595), .A2(n592), .ZN(n399) );
  NAND2_X1 U558 ( .A1(n696), .A2(G475), .ZN(n400) );
  INV_X1 U559 ( .A(n503), .ZN(n417) );
  NAND2_X1 U560 ( .A1(n503), .A2(n350), .ZN(n423) );
  NAND2_X1 U561 ( .A1(n345), .A2(n419), .ZN(n554) );
  INV_X1 U562 ( .A(n350), .ZN(n422) );
  NOR2_X1 U563 ( .A1(n503), .A2(n605), .ZN(n548) );
  NAND2_X1 U564 ( .A1(n426), .A2(n437), .ZN(n681) );
  AND2_X2 U565 ( .A1(n437), .A2(n428), .ZN(n427) );
  INV_X1 U566 ( .A(n615), .ZN(n428) );
  NAND2_X1 U567 ( .A1(n583), .A2(n584), .ZN(n431) );
  XNOR2_X1 U568 ( .A(n439), .B(KEYINPUT80), .ZN(n438) );
  NAND2_X1 U569 ( .A1(n449), .A2(KEYINPUT19), .ZN(n542) );
  NAND2_X1 U570 ( .A1(n610), .A2(n609), .ZN(n452) );
  XNOR2_X1 U571 ( .A(n454), .B(KEYINPUT63), .ZN(G57) );
  AND2_X1 U572 ( .A1(n526), .A2(G210), .ZN(n461) );
  XNOR2_X1 U573 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n462) );
  XOR2_X1 U574 ( .A(n691), .B(n690), .Z(n463) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n489), .B(n490), .ZN(n492) );
  XNOR2_X1 U577 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U578 ( .A(n692), .B(n463), .ZN(n693) );
  XNOR2_X1 U579 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U580 ( .A(n464), .B(KEYINPUT86), .ZN(n615) );
  XNOR2_X2 U581 ( .A(G128), .B(KEYINPUT65), .ZN(n465) );
  XNOR2_X2 U582 ( .A(n465), .B(G143), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U585 ( .A1(G227), .A2(n722), .ZN(n473) );
  XNOR2_X1 U586 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U587 ( .A1(G234), .A2(n615), .ZN(n477) );
  XNOR2_X1 U588 ( .A(KEYINPUT20), .B(KEYINPUT92), .ZN(n476) );
  XNOR2_X1 U589 ( .A(n477), .B(n476), .ZN(n485) );
  NAND2_X1 U590 ( .A1(G221), .A2(n485), .ZN(n478) );
  XNOR2_X1 U591 ( .A(KEYINPUT21), .B(n478), .ZN(n585) );
  XOR2_X1 U592 ( .A(G110), .B(G137), .Z(n480) );
  XNOR2_X1 U593 ( .A(n480), .B(n479), .ZN(n482) );
  NAND2_X1 U594 ( .A1(G234), .A2(n722), .ZN(n483) );
  XOR2_X1 U595 ( .A(KEYINPUT8), .B(n483), .Z(n514) );
  XNOR2_X1 U596 ( .A(KEYINPUT25), .B(KEYINPUT91), .ZN(n484) );
  NAND2_X1 U597 ( .A1(G217), .A2(n485), .ZN(n486) );
  NAND2_X1 U598 ( .A1(n564), .A2(n644), .ZN(n605) );
  XNOR2_X1 U599 ( .A(KEYINPUT73), .B(KEYINPUT5), .ZN(n488) );
  XNOR2_X1 U600 ( .A(G113), .B(KEYINPUT67), .ZN(n490) );
  NOR2_X1 U601 ( .A1(G953), .A2(G237), .ZN(n526) );
  XOR2_X1 U602 ( .A(KEYINPUT72), .B(n494), .Z(n511) );
  NAND2_X1 U603 ( .A1(G214), .A2(n511), .ZN(n663) );
  INV_X1 U604 ( .A(n663), .ZN(n495) );
  OR2_X1 U605 ( .A1(n599), .A2(n495), .ZN(n496) );
  XOR2_X1 U606 ( .A(KEYINPUT14), .B(KEYINPUT87), .Z(n498) );
  NAND2_X1 U607 ( .A1(G234), .A2(G237), .ZN(n497) );
  XNOR2_X1 U608 ( .A(n498), .B(n497), .ZN(n500) );
  NAND2_X1 U609 ( .A1(G952), .A2(n500), .ZN(n675) );
  NOR2_X1 U610 ( .A1(G953), .A2(n675), .ZN(n499) );
  XOR2_X1 U611 ( .A(KEYINPUT88), .B(n499), .Z(n577) );
  NAND2_X1 U612 ( .A1(G902), .A2(n500), .ZN(n575) );
  NOR2_X1 U613 ( .A1(G900), .A2(n575), .ZN(n501) );
  NAND2_X1 U614 ( .A1(G953), .A2(n501), .ZN(n502) );
  NAND2_X1 U615 ( .A1(n577), .A2(n502), .ZN(n543) );
  XOR2_X1 U616 ( .A(G122), .B(G104), .Z(n527) );
  XNOR2_X1 U617 ( .A(n504), .B(n527), .ZN(n505) );
  NAND2_X1 U618 ( .A1(G224), .A2(n722), .ZN(n509) );
  XNOR2_X1 U619 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n508) );
  NAND2_X1 U620 ( .A1(n687), .A2(n615), .ZN(n512) );
  XNOR2_X1 U621 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n513) );
  XNOR2_X1 U622 ( .A(n572), .B(n513), .ZN(n662) );
  NAND2_X1 U623 ( .A1(n514), .A2(G217), .ZN(n522) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n516) );
  XNOR2_X1 U625 ( .A(G116), .B(KEYINPUT102), .ZN(n515) );
  XNOR2_X1 U626 ( .A(n518), .B(G134), .ZN(n519) );
  XNOR2_X1 U627 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U628 ( .A(n522), .B(n521), .ZN(n701) );
  XOR2_X1 U629 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n524) );
  XNOR2_X1 U630 ( .A(G131), .B(KEYINPUT98), .ZN(n523) );
  XNOR2_X1 U631 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U632 ( .A(n527), .B(KEYINPUT11), .ZN(n531) );
  XOR2_X1 U633 ( .A(KEYINPUT99), .B(KEYINPUT96), .Z(n529) );
  XNOR2_X1 U634 ( .A(n529), .B(n528), .ZN(n530) );
  NOR2_X1 U635 ( .A1(G902), .A2(n698), .ZN(n537) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n535) );
  NAND2_X1 U637 ( .A1(n538), .A2(n557), .ZN(n625) );
  INV_X1 U638 ( .A(n625), .ZN(n636) );
  XNOR2_X1 U639 ( .A(KEYINPUT105), .B(n636), .ZN(n539) );
  INV_X1 U640 ( .A(n634), .ZN(n631) );
  NAND2_X1 U641 ( .A1(n631), .A2(n539), .ZN(n660) );
  INV_X1 U642 ( .A(n660), .ZN(n607) );
  INV_X1 U643 ( .A(KEYINPUT19), .ZN(n540) );
  NAND2_X1 U644 ( .A1(n542), .A2(n541), .ZN(n579) );
  XOR2_X1 U645 ( .A(KEYINPUT28), .B(n544), .Z(n546) );
  XNOR2_X1 U646 ( .A(n564), .B(KEYINPUT109), .ZN(n545) );
  NOR2_X1 U647 ( .A1(n546), .A2(n545), .ZN(n560) );
  NAND2_X1 U648 ( .A1(n579), .A2(n560), .ZN(n630) );
  NOR2_X1 U649 ( .A1(n607), .A2(n630), .ZN(n547) );
  XNOR2_X1 U650 ( .A(n547), .B(KEYINPUT47), .ZN(n552) );
  AND2_X1 U651 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U652 ( .A(KEYINPUT108), .B(n550), .ZN(n551) );
  NOR2_X1 U653 ( .A1(n558), .A2(n557), .ZN(n574) );
  NAND2_X1 U654 ( .A1(n551), .A2(n574), .ZN(n629) );
  NAND2_X1 U655 ( .A1(n552), .A2(n629), .ZN(n553) );
  XOR2_X1 U656 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n563) );
  XOR2_X1 U657 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n562) );
  NAND2_X1 U658 ( .A1(n662), .A2(n663), .ZN(n556) );
  NAND2_X1 U659 ( .A1(n558), .A2(n557), .ZN(n665) );
  INV_X1 U660 ( .A(n665), .ZN(n559) );
  INV_X1 U661 ( .A(n643), .ZN(n594) );
  NOR2_X1 U662 ( .A1(n440), .A2(n569), .ZN(n570) );
  NAND2_X1 U663 ( .A1(n570), .A2(n663), .ZN(n571) );
  XNOR2_X1 U664 ( .A(n571), .B(KEYINPUT43), .ZN(n573) );
  NAND2_X1 U665 ( .A1(n573), .A2(n572), .ZN(n642) );
  XNOR2_X1 U666 ( .A(KEYINPUT76), .B(n574), .ZN(n584) );
  NOR2_X1 U667 ( .A1(G898), .A2(n722), .ZN(n709) );
  INV_X1 U668 ( .A(n575), .ZN(n576) );
  NAND2_X1 U669 ( .A1(n709), .A2(n576), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U671 ( .A(n600), .B(KEYINPUT89), .Z(n603) );
  XNOR2_X1 U672 ( .A(n582), .B(KEYINPUT34), .ZN(n583) );
  NOR2_X1 U673 ( .A1(n600), .A2(n665), .ZN(n586) );
  INV_X1 U674 ( .A(n585), .ZN(n646) );
  NAND2_X1 U675 ( .A1(n591), .A2(n587), .ZN(n588) );
  XOR2_X1 U676 ( .A(n591), .B(KEYINPUT106), .Z(n647) );
  NOR2_X1 U677 ( .A1(n594), .A2(n647), .ZN(n592) );
  NAND2_X1 U678 ( .A1(n594), .A2(n647), .ZN(n597) );
  XNOR2_X1 U679 ( .A(KEYINPUT83), .B(n595), .ZN(n596) );
  NOR2_X1 U680 ( .A1(n597), .A2(n596), .ZN(n618) );
  OR2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n654) );
  NOR2_X1 U682 ( .A1(n600), .A2(n654), .ZN(n602) );
  XNOR2_X1 U683 ( .A(KEYINPUT95), .B(KEYINPUT31), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n602), .B(n601), .ZN(n637) );
  OR2_X1 U685 ( .A1(n650), .A2(n603), .ZN(n604) );
  NOR2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n620) );
  NOR2_X1 U687 ( .A1(n637), .A2(n620), .ZN(n606) );
  NOR2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U689 ( .A1(n618), .A2(n608), .ZN(n609) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n612) );
  XNOR2_X1 U691 ( .A(KEYINPUT78), .B(n613), .ZN(n614) );
  XOR2_X1 U692 ( .A(n616), .B(KEYINPUT85), .Z(n617) );
  XOR2_X1 U693 ( .A(G101), .B(n618), .Z(G3) );
  NAND2_X1 U694 ( .A1(n620), .A2(n634), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n619), .B(G104), .ZN(G6) );
  XOR2_X1 U696 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n622) );
  NAND2_X1 U697 ( .A1(n620), .A2(n636), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U699 ( .A(G107), .B(n623), .ZN(G9) );
  XOR2_X1 U700 ( .A(n624), .B(G110), .Z(G12) );
  NOR2_X1 U701 ( .A1(n625), .A2(n630), .ZN(n627) );
  XNOR2_X1 U702 ( .A(KEYINPUT29), .B(KEYINPUT112), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U704 ( .A(G128), .B(n628), .ZN(G30) );
  XNOR2_X1 U705 ( .A(G143), .B(n629), .ZN(G45) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n633) );
  XNOR2_X1 U707 ( .A(G146), .B(KEYINPUT113), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n633), .B(n632), .ZN(G48) );
  NAND2_X1 U709 ( .A1(n637), .A2(n634), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n635), .B(G113), .ZN(G15) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n638), .B(G116), .ZN(G18) );
  XNOR2_X1 U713 ( .A(G125), .B(n639), .ZN(n640) );
  XNOR2_X1 U714 ( .A(n640), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U715 ( .A(G134), .B(n641), .Z(G36) );
  XNOR2_X1 U716 ( .A(G140), .B(n642), .ZN(G42) );
  NOR2_X1 U717 ( .A1(n644), .A2(n440), .ZN(n645) );
  XOR2_X1 U718 ( .A(KEYINPUT50), .B(n645), .Z(n653) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U720 ( .A(KEYINPUT49), .B(n648), .Z(n649) );
  NOR2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U722 ( .A(KEYINPUT114), .B(n651), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n656), .B(KEYINPUT115), .ZN(n657) );
  XNOR2_X1 U726 ( .A(KEYINPUT51), .B(n657), .ZN(n658) );
  NAND2_X1 U727 ( .A1(n658), .A2(n676), .ZN(n672) );
  NAND2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U729 ( .A(KEYINPUT117), .B(n661), .ZN(n668) );
  NOR2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U731 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U732 ( .A(n666), .B(KEYINPUT116), .ZN(n667) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U734 ( .A1(n669), .A2(n677), .ZN(n670) );
  XOR2_X1 U735 ( .A(KEYINPUT118), .B(n670), .Z(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U737 ( .A(KEYINPUT52), .B(n673), .Z(n674) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n680) );
  INV_X1 U739 ( .A(n676), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U743 ( .A1(G953), .A2(n683), .ZN(n685) );
  XNOR2_X1 U744 ( .A(KEYINPUT53), .B(KEYINPUT119), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n685), .B(n684), .ZN(n686) );
  XOR2_X1 U746 ( .A(KEYINPUT120), .B(n686), .Z(G75) );
  XOR2_X1 U747 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n689) );
  NAND2_X1 U748 ( .A1(n696), .A2(G469), .ZN(n694) );
  XOR2_X1 U749 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n691) );
  XNOR2_X1 U750 ( .A(KEYINPUT122), .B(KEYINPUT121), .ZN(n690) );
  NOR2_X1 U751 ( .A1(n706), .A2(n695), .ZN(G54) );
  INV_X1 U752 ( .A(KEYINPUT59), .ZN(n697) );
  NAND2_X1 U753 ( .A1(G478), .A2(n696), .ZN(n700) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n706), .A2(n702), .ZN(G63) );
  NAND2_X1 U756 ( .A1(G217), .A2(n696), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n706), .A2(n705), .ZN(G66) );
  XNOR2_X1 U759 ( .A(KEYINPUT125), .B(n707), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(KEYINPUT124), .B(n710), .ZN(n718) );
  XOR2_X1 U762 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n712) );
  NAND2_X1 U763 ( .A1(G224), .A2(G953), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n713), .A2(G898), .ZN(n716) );
  NAND2_X1 U766 ( .A1(n714), .A2(n722), .ZN(n715) );
  NAND2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U769 ( .A(n719), .B(n720), .Z(n724) );
  XOR2_X1 U770 ( .A(n721), .B(n724), .Z(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(n722), .ZN(n728) );
  XNOR2_X1 U772 ( .A(G227), .B(n724), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n725), .A2(G900), .ZN(n726) );
  NAND2_X1 U774 ( .A1(G953), .A2(n726), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U776 ( .A(KEYINPUT126), .B(n729), .ZN(G72) );
  XNOR2_X1 U777 ( .A(n730), .B(G119), .ZN(G21) );
  XOR2_X1 U778 ( .A(G131), .B(n731), .Z(n732) );
  XNOR2_X1 U779 ( .A(KEYINPUT127), .B(n732), .ZN(G33) );
  XNOR2_X1 U780 ( .A(G137), .B(n733), .ZN(G39) );
endmodule

