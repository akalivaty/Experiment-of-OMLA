//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n206), .A2(new_n208), .B1(KEYINPUT2), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211));
  INV_X1    g010(.A(new_n209), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(KEYINPUT79), .A3(new_n209), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n209), .ZN(new_n220));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n209), .A2(KEYINPUT2), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n220), .B(new_n211), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n204), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n219), .A2(new_n223), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(KEYINPUT80), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT74), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(KEYINPUT74), .ZN(new_n234));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(G211gat), .B(G218gat), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n237), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n239), .A2(new_n233), .A3(new_n234), .A4(new_n235), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n231), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT82), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n238), .A2(new_n244), .A3(new_n240), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n230), .B1(new_n240), .B2(new_n244), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n227), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n224), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n203), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n241), .B1(new_n229), .B2(new_n230), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT29), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n241), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n203), .B1(new_n252), .B2(new_n226), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(G22gat), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G22gat), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n231), .A2(new_n242), .B1(new_n224), .B2(new_n247), .ZN(new_n257));
  OAI221_X1 g056(.A(new_n256), .B1(new_n250), .B2(new_n253), .C1(new_n257), .C2(new_n203), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n257), .A2(new_n203), .B1(new_n250), .B2(new_n253), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT83), .B1(new_n260), .B2(G22gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT31), .B(G50gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n259), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n255), .A2(new_n258), .A3(KEYINPUT83), .A4(new_n264), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT24), .ZN(new_n269));
  INV_X1    g068(.A(G183gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G190gat), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G183gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n269), .A2(G183gat), .A3(G190gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT65), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  OR3_X1    g076(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(G169gat), .A2(G176gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(G169gat), .A3(G176gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n278), .A2(new_n279), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n285));
  XNOR2_X1  g084(.A(G183gat), .B(G190gat), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n285), .B(new_n275), .C1(new_n286), .C2(new_n269), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n277), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n276), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n284), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n270), .A2(KEYINPUT27), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n272), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G183gat), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT67), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n294), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n295), .A2(new_n299), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(KEYINPUT28), .A3(new_n272), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n301), .A2(new_n303), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n281), .A2(new_n283), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT68), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n308), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT69), .ZN(new_n311));
  OR3_X1    g110(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n305), .A2(new_n307), .A3(new_n313), .A4(new_n309), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n311), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n304), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n293), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G120gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G113gat), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G120gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT70), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n319), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT1), .B1(new_n324), .B2(KEYINPUT70), .ZN(new_n325));
  NAND2_X1  g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(G127gat), .A2(G134gat), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT71), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n330));
  INV_X1    g129(.A(G127gat), .ZN(new_n331));
  INV_X1    g130(.A(G134gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n330), .B1(new_n333), .B2(new_n326), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n323), .B(new_n325), .C1(new_n329), .C2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n319), .A2(new_n321), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n333), .B(new_n326), .C1(new_n336), .C2(KEYINPUT1), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g138(.A1(G227gat), .A2(G233gat), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n290), .A2(new_n292), .B1(new_n304), .B2(new_n315), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n335), .A2(new_n337), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT33), .ZN(new_n345));
  XNOR2_X1  g144(.A(G15gat), .B(G43gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G71gat), .B(G99gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n344), .B(KEYINPUT32), .C1(new_n345), .C2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n344), .B2(KEYINPUT32), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(new_n351), .A3(new_n345), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n344), .B2(new_n345), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n340), .B1(new_n339), .B2(new_n343), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT34), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n355), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n355), .B2(new_n356), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n268), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT90), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n226), .A2(new_n335), .A3(new_n366), .A4(new_n337), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT81), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT4), .B1(new_n342), .B2(new_n224), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(KEYINPUT81), .B(KEYINPUT4), .C1(new_n342), .C2(new_n224), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n338), .B1(KEYINPUT3), .B2(new_n224), .ZN(new_n372));
  AOI22_X1  g171(.A1(new_n370), .A2(new_n371), .B1(new_n372), .B2(new_n229), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT5), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n229), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n369), .A2(new_n367), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n342), .B(new_n224), .ZN(new_n380));
  INV_X1    g179(.A(new_n375), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT0), .ZN(new_n386));
  XNOR2_X1  g185(.A(G57gat), .B(G85gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n386), .B(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390));
  INV_X1    g189(.A(new_n388), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n383), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n384), .A2(KEYINPUT6), .A3(new_n388), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT75), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n230), .ZN(new_n400));
  OAI211_X1 g199(.A(KEYINPUT77), .B(new_n399), .C1(new_n341), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n398), .B1(new_n317), .B2(new_n230), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT77), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n403), .B1(new_n317), .B2(new_n398), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n401), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n242), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n399), .B1(new_n341), .B2(KEYINPUT29), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n317), .A2(new_n398), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n241), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT78), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n407), .A2(new_n408), .A3(new_n411), .A4(new_n241), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G8gat), .B(G36gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OR3_X1    g216(.A1(new_n413), .A2(KEYINPUT30), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n417), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n406), .A2(new_n416), .A3(new_n410), .A4(new_n412), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(KEYINPUT30), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n396), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n268), .B(KEYINPUT90), .C1(new_n361), .C2(new_n362), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n365), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT35), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n355), .B(new_n360), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT89), .B(KEYINPUT35), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n393), .B2(new_n394), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n268), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n418), .A3(KEYINPUT84), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(new_n418), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT88), .A3(new_n417), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT88), .B1(new_n437), .B2(new_n417), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT38), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n393), .A2(new_n394), .A3(new_n420), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n439), .A2(KEYINPUT38), .A3(new_n416), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n407), .A2(new_n242), .A3(new_n408), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n241), .B2(new_n405), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n448), .B(KEYINPUT87), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n444), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n370), .A2(new_n371), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n377), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n381), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT39), .ZN(new_n455));
  INV_X1    g254(.A(new_n380), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n375), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n373), .A2(KEYINPUT39), .A3(new_n375), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n459), .A2(KEYINPUT85), .A3(new_n388), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n455), .A3(new_n381), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n462), .B2(new_n391), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT40), .B(new_n458), .C1(new_n460), .C2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n389), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT85), .B1(new_n459), .B2(new_n388), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n462), .A2(new_n461), .A3(new_n391), .ZN(new_n467));
  AOI22_X1  g266(.A1(new_n466), .A2(new_n467), .B1(new_n454), .B2(new_n457), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT86), .B1(new_n468), .B2(KEYINPUT40), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n458), .B1(new_n460), .B2(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT40), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n465), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n433), .A2(new_n474), .A3(new_n430), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n451), .A2(new_n475), .A3(new_n268), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n422), .A2(new_n268), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT36), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n426), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n362), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n355), .A2(new_n356), .A3(new_n360), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT36), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n436), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  AND2_X1   g286(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G50gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G43gat), .ZN(new_n496));
  INV_X1    g295(.A(G43gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G50gat), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(KEYINPUT92), .A3(G50gat), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT93), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n496), .A2(new_n498), .A3(KEYINPUT15), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n494), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n505), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n502), .A4(new_n501), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n510), .B2(new_n493), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT17), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(G1gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT16), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G1gat), .B2(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G8gat), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n516), .B(new_n519), .C1(G1gat), .C2(new_n513), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n510), .A2(new_n493), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(new_n505), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n495), .A2(G43gat), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT15), .B1(new_n525), .B2(KEYINPUT92), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n509), .B1(new_n526), .B2(new_n508), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n493), .B1(new_n527), .B2(new_n507), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n522), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n506), .A2(new_n511), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n521), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n524), .A2(new_n528), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n532), .B(KEYINPUT13), .Z(new_n540));
  AOI22_X1  g339(.A1(new_n535), .A2(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n532), .A4(new_n534), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT11), .B(G169gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT12), .Z(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n546), .B2(new_n547), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT95), .B1(new_n486), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n546), .A2(new_n547), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n552), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n554), .ZN(new_n562));
  AOI211_X1 g361(.A(new_n559), .B(new_n562), .C1(new_n436), .C2(new_n485), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n558), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT98), .ZN(new_n565));
  AND2_X1   g364(.A1(G57gat), .A2(G64gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(G57gat), .A2(G64gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT97), .ZN(new_n569));
  NAND2_X1  g368(.A1(G71gat), .A2(G78gat), .ZN(new_n570));
  OR2_X1    g369(.A1(G71gat), .A2(G78gat), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n568), .A2(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT9), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n570), .A2(KEYINPUT96), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT96), .B1(new_n570), .B2(new_n573), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n568), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G57gat), .B(G64gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n570), .A2(new_n573), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n570), .A2(KEYINPUT96), .A3(new_n573), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(G57gat), .A2(G64gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(G57gat), .A2(G64gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n569), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n570), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n565), .B1(new_n577), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n576), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n582), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n592), .A3(new_n568), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n593), .A3(KEYINPUT98), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(G231gat), .B(G233gat), .C1(new_n595), .C2(KEYINPUT21), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n590), .A2(new_n597), .A3(new_n594), .A4(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n331), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n521), .B1(new_n595), .B2(KEYINPUT21), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n596), .A2(new_n331), .A3(new_n599), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n603), .B1(new_n601), .B2(new_n604), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n215), .ZN(new_n608));
  XOR2_X1   g407(.A(G183gat), .B(G211gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OR3_X1    g410(.A1(new_n605), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n605), .B2(new_n606), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT7), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  INV_X1    g416(.A(G85gat), .ZN(new_n618));
  INV_X1    g417(.A(G92gat), .ZN(new_n619));
  AOI22_X1  g418(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G99gat), .B(G106gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n624), .A2(new_n616), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n512), .A2(new_n530), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n512), .A2(new_n530), .A3(KEYINPUT99), .A4(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n537), .B2(new_n626), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G190gat), .B(G218gat), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n639));
  XNOR2_X1  g438(.A(G134gat), .B(G162gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n637), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n631), .A2(new_n642), .A3(new_n635), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n641), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(new_n631), .B2(new_n635), .ZN(new_n646));
  AOI211_X1 g445(.A(new_n637), .B(new_n634), .C1(new_n629), .C2(new_n630), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n591), .A2(new_n593), .A3(KEYINPUT98), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT98), .B1(new_n591), .B2(new_n593), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n626), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n623), .A2(new_n591), .A3(new_n593), .A4(new_n625), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT10), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n595), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n650), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n654), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n595), .B2(new_n626), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n658), .B1(new_n650), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n658), .B(new_n665), .C1(new_n650), .C2(new_n661), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n614), .A2(new_n649), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n564), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n395), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(new_n514), .ZN(G1324gat));
  INV_X1    g474(.A(new_n673), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n421), .A2(new_n418), .A3(KEYINPUT84), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT84), .B1(new_n421), .B2(new_n418), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n519), .B1(new_n676), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n673), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  INV_X1    g484(.A(new_n426), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n673), .A2(G15gat), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n483), .ZN(new_n688));
  OAI21_X1  g487(.A(G15gat), .B1(new_n673), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n673), .A2(new_n268), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n614), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n670), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(new_n649), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n564), .A2(new_n491), .A3(new_n396), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT45), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n699));
  INV_X1    g498(.A(new_n649), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n479), .B(new_n482), .C1(new_n422), .C2(new_n268), .ZN(new_n701));
  INV_X1    g500(.A(new_n268), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n702), .B1(new_n679), .B2(new_n474), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n701), .B1(new_n703), .B2(new_n451), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n434), .B1(KEYINPUT35), .B2(new_n424), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n699), .B(new_n700), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n695), .A2(new_n562), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n649), .B1(new_n436), .B2(new_n485), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT100), .B1(new_n711), .B2(new_n699), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT100), .B(new_n700), .C1(new_n704), .C2(new_n705), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT44), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n709), .B(new_n710), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G29gat), .B1(new_n715), .B2(new_n395), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n698), .A2(KEYINPUT102), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(G1328gat));
  OAI21_X1  g520(.A(new_n696), .B1(new_n558), .B2(new_n563), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n722), .A2(G36gat), .A3(new_n681), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n715), .B2(new_n681), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1329gat));
  OAI21_X1  g528(.A(new_n497), .B1(new_n722), .B2(new_n686), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n483), .A2(G43gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n715), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g532(.A(G50gat), .B1(new_n715), .B2(new_n268), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n739), .B(new_n696), .C1(new_n558), .C2(new_n563), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n268), .A2(G50gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n742), .A2(new_n734), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n742), .B2(new_n734), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(new_n734), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(KEYINPUT106), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT48), .B1(new_n734), .B2(KEYINPUT105), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n742), .A2(new_n734), .A3(new_n743), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n746), .A2(new_n751), .ZN(G1331gat));
  NAND4_X1  g551(.A1(new_n614), .A2(new_n562), .A3(new_n649), .A4(new_n669), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n753), .B1(new_n436), .B2(new_n485), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n396), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g555(.A(new_n681), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(KEYINPUT107), .Z(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1333gat));
  NAND2_X1  g560(.A1(new_n754), .A2(new_n483), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n686), .A2(G71gat), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n762), .A2(G71gat), .B1(new_n754), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n754), .A2(new_n702), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g566(.A1(new_n614), .A2(new_n557), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n711), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n711), .A2(KEYINPUT51), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT108), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n774), .A2(new_n618), .A3(new_n396), .A4(new_n669), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n706), .A2(new_n707), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(KEYINPUT44), .A3(new_n713), .ZN(new_n777));
  INV_X1    g576(.A(new_n768), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(new_n670), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n709), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780), .B2(new_n395), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n775), .A2(new_n781), .ZN(G1336gat));
  AND4_X1   g581(.A1(new_n619), .A2(new_n773), .A3(new_n679), .A4(new_n669), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n777), .A2(new_n679), .A3(new_n709), .A4(new_n779), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(G92gat), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT109), .B1(new_n784), .B2(G92gat), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n785), .B(new_n787), .ZN(G1337gat));
  NOR3_X1   g587(.A1(new_n686), .A2(G99gat), .A3(new_n670), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT110), .Z(new_n790));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G99gat), .B1(new_n780), .B2(new_n688), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1338gat));
  OAI21_X1  g592(.A(G106gat), .B1(new_n780), .B2(new_n268), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n268), .A2(G106gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n669), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  INV_X1    g599(.A(new_n650), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n595), .A2(new_n656), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n801), .B(new_n802), .C1(new_n660), .C2(KEYINPUT10), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n658), .A2(new_n803), .A3(KEYINPUT54), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n805), .B(new_n650), .C1(new_n655), .C2(new_n657), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n666), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n668), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n806), .A2(new_n666), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n809), .B2(new_n804), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n539), .A2(new_n540), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n532), .B1(new_n531), .B2(new_n534), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n551), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n541), .B(new_n553), .C1(new_n544), .C2(new_n545), .ZN(new_n815));
  AND4_X1   g614(.A1(new_n644), .A2(new_n648), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n800), .B1(new_n811), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n658), .A2(new_n803), .A3(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n806), .A2(new_n666), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n821), .A2(new_n668), .A3(new_n807), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n644), .A2(new_n648), .A3(new_n814), .A4(new_n815), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT112), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n669), .A2(new_n814), .A3(new_n815), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(new_n562), .B2(new_n822), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n649), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n614), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n671), .A2(new_n557), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT113), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n808), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(new_n561), .A3(new_n554), .A4(new_n821), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n700), .B1(new_n833), .B2(new_n826), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n811), .A2(new_n816), .A3(new_n800), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT112), .B1(new_n822), .B2(new_n823), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n694), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n672), .A2(new_n562), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n831), .A2(new_n841), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n842), .A2(new_n268), .A3(new_n426), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n396), .A3(new_n681), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n320), .A3(new_n562), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n842), .A2(new_n396), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n365), .A3(new_n423), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT114), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n681), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n557), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n845), .B1(new_n850), .B2(new_n320), .ZN(G1340gat));
  NOR3_X1   g650(.A1(new_n844), .A2(new_n318), .A3(new_n670), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n669), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n318), .ZN(G1341gat));
  NAND3_X1  g653(.A1(new_n849), .A2(new_n331), .A3(new_n614), .ZN(new_n855));
  OAI21_X1  g654(.A(G127gat), .B1(new_n844), .B2(new_n694), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NOR2_X1   g656(.A1(new_n679), .A2(new_n649), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n848), .A2(new_n332), .A3(new_n858), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g659(.A(G134gat), .B1(new_n844), .B2(new_n649), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(G1343gat));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n702), .A3(new_n688), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n679), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n205), .A3(new_n557), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n864), .B1(new_n867), .B2(KEYINPUT118), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT115), .B1(new_n819), .B2(new_n820), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n809), .A2(new_n871), .A3(new_n804), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n818), .A3(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n870), .A2(new_n872), .A3(KEYINPUT116), .A4(new_n818), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n875), .A2(new_n557), .A3(new_n832), .A4(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n700), .B1(new_n877), .B2(new_n826), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n694), .B1(new_n878), .B2(new_n837), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n840), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n869), .B1(new_n883), .B2(new_n702), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n842), .A2(new_n869), .A3(new_n702), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n483), .A2(new_n679), .A3(new_n395), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n884), .A2(new_n887), .A3(new_n562), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n867), .B1(new_n888), .B2(new_n205), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n868), .B(new_n889), .ZN(G1344gat));
  NAND3_X1  g689(.A1(new_n866), .A2(new_n207), .A3(new_n669), .ZN(new_n891));
  XNOR2_X1  g690(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n822), .A2(new_n823), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n694), .B1(new_n878), .B2(new_n894), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n895), .A2(KEYINPUT121), .A3(new_n840), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT121), .B1(new_n895), .B2(new_n840), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n896), .A2(new_n897), .A3(new_n268), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n893), .B1(new_n898), .B2(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n840), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n268), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n895), .A2(KEYINPUT121), .A3(new_n840), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(KEYINPUT122), .A3(new_n869), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n831), .A2(KEYINPUT57), .A3(new_n702), .A4(new_n841), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT120), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n899), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n669), .A3(new_n886), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n892), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n884), .A2(new_n887), .A3(new_n670), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(KEYINPUT59), .A3(new_n207), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n891), .B1(new_n910), .B2(new_n912), .ZN(G1345gat));
  NAND3_X1  g712(.A1(new_n866), .A2(new_n215), .A3(new_n614), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n884), .A2(new_n887), .A3(new_n694), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n215), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n884), .A2(new_n887), .A3(new_n649), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n858), .A2(new_n216), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n917), .A2(new_n216), .B1(new_n865), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n681), .A2(new_n396), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n843), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(G169gat), .B1(new_n921), .B2(new_n562), .ZN(new_n922));
  XOR2_X1   g721(.A(new_n922), .B(KEYINPUT123), .Z(new_n923));
  AND2_X1   g722(.A1(new_n842), .A2(new_n395), .ZN(new_n924));
  AND4_X1   g723(.A1(new_n679), .A2(new_n924), .A3(new_n365), .A4(new_n423), .ZN(new_n925));
  INV_X1    g724(.A(G169gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n557), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n923), .A2(new_n927), .ZN(G1348gat));
  INV_X1    g727(.A(G176gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n929), .A3(new_n669), .ZN(new_n930));
  OAI21_X1  g729(.A(G176gat), .B1(new_n921), .B2(new_n670), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n925), .A2(new_n302), .A3(new_n614), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n921), .B2(new_n694), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G183gat), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n921), .A2(KEYINPUT124), .A3(new_n694), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n921), .B2(new_n649), .ZN(new_n939));
  XOR2_X1   g738(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n272), .A3(new_n700), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1351gat));
  NOR3_X1   g742(.A1(new_n681), .A2(new_n268), .A3(new_n483), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n924), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(G197gat), .B1(new_n946), .B2(new_n557), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n920), .A2(new_n688), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n908), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n557), .A2(G197gat), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(G1352gat));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n669), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G204gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n945), .A2(G204gat), .A3(new_n670), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  OR3_X1    g756(.A1(new_n945), .A2(G211gat), .A3(new_n694), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n908), .A2(KEYINPUT126), .A3(new_n614), .A4(new_n949), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(G211gat), .ZN(new_n960));
  AOI21_X1  g759(.A(KEYINPUT57), .B1(new_n902), .B2(new_n903), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n963));
  OAI22_X1  g762(.A1(new_n961), .A2(KEYINPUT122), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n898), .A2(new_n893), .A3(KEYINPUT57), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n614), .B(new_n949), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(KEYINPUT63), .B1(new_n960), .B2(new_n968), .ZN(new_n969));
  AND4_X1   g768(.A1(KEYINPUT63), .A2(new_n968), .A3(G211gat), .A4(new_n959), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n958), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  INV_X1    g770(.A(G218gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n972), .B1(new_n945), .B2(new_n649), .ZN(new_n973));
  XOR2_X1   g772(.A(new_n973), .B(KEYINPUT127), .Z(new_n974));
  NOR2_X1   g773(.A1(new_n649), .A2(new_n972), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n950), .B2(new_n975), .ZN(G1355gat));
endmodule


