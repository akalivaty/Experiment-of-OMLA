

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U545 ( .A1(n718), .A2(n710), .ZN(n711) );
  NOR2_X2 U546 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  NOR2_X2 U547 ( .A1(n546), .A2(n545), .ZN(G160) );
  XNOR2_X1 U548 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n539) );
  OR2_X1 U549 ( .A1(n712), .A2(G168), .ZN(n713) );
  AND2_X1 U550 ( .A1(n534), .A2(n533), .ZN(n863) );
  XOR2_X1 U551 ( .A(KEYINPUT28), .B(n679), .Z(n511) );
  NAND2_X1 U552 ( .A1(n793), .A2(n792), .ZN(n512) );
  NOR2_X1 U553 ( .A1(n742), .A2(n791), .ZN(n513) );
  AND2_X1 U554 ( .A1(n794), .A2(n512), .ZN(n514) );
  INV_X1 U555 ( .A(n726), .ZN(n693) );
  NAND2_X1 U556 ( .A1(n674), .A2(n757), .ZN(n726) );
  NOR2_X1 U557 ( .A1(G164), .A2(G1384), .ZN(n757) );
  NOR2_X1 U558 ( .A1(G651), .A2(n632), .ZN(n635) );
  XNOR2_X1 U559 ( .A(n540), .B(n539), .ZN(n542) );
  NOR2_X1 U560 ( .A1(n538), .A2(n537), .ZN(G164) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n640) );
  NAND2_X1 U562 ( .A1(n640), .A2(G89), .ZN(n515) );
  XNOR2_X1 U563 ( .A(KEYINPUT4), .B(n515), .ZN(n518) );
  XOR2_X1 U564 ( .A(G543), .B(KEYINPUT0), .Z(n632) );
  INV_X1 U565 ( .A(G651), .ZN(n520) );
  NOR2_X1 U566 ( .A1(n632), .A2(n520), .ZN(n637) );
  NAND2_X1 U567 ( .A1(n637), .A2(G76), .ZN(n516) );
  XOR2_X1 U568 ( .A(KEYINPUT73), .B(n516), .Z(n517) );
  NAND2_X1 U569 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U570 ( .A(n519), .B(KEYINPUT5), .ZN(n526) );
  NOR2_X1 U571 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n521), .Z(n636) );
  NAND2_X1 U573 ( .A1(G63), .A2(n636), .ZN(n523) );
  NAND2_X1 U574 ( .A1(G51), .A2(n635), .ZN(n522) );
  NAND2_X1 U575 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT6), .B(n524), .Z(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U578 ( .A(n527), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U579 ( .A(KEYINPUT64), .B(G2104), .ZN(n534) );
  INV_X1 U580 ( .A(G2105), .ZN(n533) );
  NOR2_X2 U581 ( .A1(n534), .A2(n533), .ZN(n868) );
  NAND2_X1 U582 ( .A1(G126), .A2(n868), .ZN(n528) );
  XNOR2_X1 U583 ( .A(n528), .B(KEYINPUT86), .ZN(n532) );
  XOR2_X2 U584 ( .A(KEYINPUT17), .B(n529), .Z(n864) );
  NAND2_X1 U585 ( .A1(n864), .A2(G138), .ZN(n530) );
  XOR2_X1 U586 ( .A(n530), .B(KEYINPUT87), .Z(n531) );
  NAND2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n538) );
  AND2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n867) );
  NAND2_X1 U589 ( .A1(G114), .A2(n867), .ZN(n536) );
  NAND2_X1 U590 ( .A1(G102), .A2(n863), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U592 ( .A1(G101), .A2(n863), .ZN(n540) );
  NAND2_X1 U593 ( .A1(G113), .A2(n867), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U595 ( .A1(G137), .A2(n864), .ZN(n544) );
  NAND2_X1 U596 ( .A1(G125), .A2(n868), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U598 ( .A1(G72), .A2(n637), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G85), .A2(n640), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U601 ( .A1(G60), .A2(n636), .ZN(n550) );
  NAND2_X1 U602 ( .A1(G47), .A2(n635), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U604 ( .A1(n552), .A2(n551), .ZN(G290) );
  XNOR2_X1 U605 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G77), .A2(n637), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G90), .A2(n640), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n556), .B(n555), .ZN(n561) );
  NAND2_X1 U610 ( .A1(n636), .A2(G64), .ZN(n557) );
  XNOR2_X1 U611 ( .A(n557), .B(KEYINPUT66), .ZN(n559) );
  NAND2_X1 U612 ( .A1(G52), .A2(n635), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U614 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U619 ( .A(n562), .B(KEYINPUT10), .ZN(n563) );
  XNOR2_X1 U620 ( .A(KEYINPUT70), .B(n563), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n813) );
  NAND2_X1 U622 ( .A1(n813), .A2(G567), .ZN(n564) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U624 ( .A1(n636), .A2(G56), .ZN(n565) );
  XOR2_X1 U625 ( .A(KEYINPUT14), .B(n565), .Z(n573) );
  NAND2_X1 U626 ( .A1(G68), .A2(n637), .ZN(n569) );
  XOR2_X1 U627 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n567) );
  NAND2_X1 U628 ( .A1(G81), .A2(n640), .ZN(n566) );
  XNOR2_X1 U629 ( .A(n567), .B(n566), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT72), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT13), .B(n571), .Z(n572) );
  NOR2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n635), .A2(G43), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n910) );
  INV_X1 U636 ( .A(G860), .ZN(n594) );
  OR2_X1 U637 ( .A1(n910), .A2(n594), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n584) );
  NAND2_X1 U640 ( .A1(G92), .A2(n640), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G54), .A2(n635), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G66), .A2(n636), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G79), .A2(n637), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(KEYINPUT15), .ZN(n918) );
  INV_X1 U648 ( .A(G868), .ZN(n647) );
  NAND2_X1 U649 ( .A1(n918), .A2(n647), .ZN(n583) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G78), .A2(n637), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G91), .A2(n640), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT68), .B(n587), .Z(n591) );
  NAND2_X1 U655 ( .A1(G65), .A2(n636), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G53), .A2(n635), .ZN(n588) );
  AND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(G299) );
  XOR2_X1 U659 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U661 ( .A1(G286), .A2(n647), .ZN(n592) );
  NOR2_X1 U662 ( .A1(n593), .A2(n592), .ZN(G297) );
  NAND2_X1 U663 ( .A1(n594), .A2(G559), .ZN(n595) );
  INV_X1 U664 ( .A(n918), .ZN(n884) );
  NAND2_X1 U665 ( .A1(n595), .A2(n884), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n596), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U667 ( .A1(G868), .A2(n910), .ZN(n599) );
  NAND2_X1 U668 ( .A1(n884), .A2(G868), .ZN(n597) );
  NOR2_X1 U669 ( .A1(G559), .A2(n597), .ZN(n598) );
  NOR2_X1 U670 ( .A1(n599), .A2(n598), .ZN(G282) );
  XNOR2_X1 U671 ( .A(G2100), .B(KEYINPUT75), .ZN(n609) );
  NAND2_X1 U672 ( .A1(G111), .A2(n867), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G135), .A2(n864), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G123), .A2(n868), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n602), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G99), .A2(n863), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT74), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n987) );
  XNOR2_X1 U681 ( .A(n987), .B(G2096), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U683 ( .A(KEYINPUT76), .B(n610), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G559), .A2(n884), .ZN(n611) );
  XNOR2_X1 U685 ( .A(n611), .B(n910), .ZN(n654) );
  NOR2_X1 U686 ( .A1(n654), .A2(G860), .ZN(n620) );
  NAND2_X1 U687 ( .A1(G80), .A2(n637), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G93), .A2(n640), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n614), .B(KEYINPUT77), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G67), .A2(n636), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n635), .A2(G55), .ZN(n617) );
  XOR2_X1 U694 ( .A(KEYINPUT78), .B(n617), .Z(n618) );
  NOR2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n650) );
  XNOR2_X1 U696 ( .A(n620), .B(n650), .ZN(G145) );
  NAND2_X1 U697 ( .A1(G73), .A2(n637), .ZN(n621) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT2), .ZN(n628) );
  NAND2_X1 U699 ( .A1(G61), .A2(n636), .ZN(n623) );
  NAND2_X1 U700 ( .A1(G86), .A2(n640), .ZN(n622) );
  NAND2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U702 ( .A1(G48), .A2(n635), .ZN(n624) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n624), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(G305) );
  NAND2_X1 U706 ( .A1(G49), .A2(n635), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n636), .A2(n631), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U712 ( .A1(G50), .A2(n635), .ZN(n645) );
  NAND2_X1 U713 ( .A1(G62), .A2(n636), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G75), .A2(n637), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n640), .A2(G88), .ZN(n641) );
  XOR2_X1 U717 ( .A(KEYINPUT80), .B(n641), .Z(n642) );
  NOR2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT81), .ZN(G166) );
  NAND2_X1 U721 ( .A1(n647), .A2(n650), .ZN(n658) );
  XNOR2_X1 U722 ( .A(KEYINPUT19), .B(G305), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n648), .B(G288), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n650), .B(n649), .ZN(n652) );
  XNOR2_X1 U725 ( .A(G290), .B(G166), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U727 ( .A(n653), .B(G299), .ZN(n883) );
  XNOR2_X1 U728 ( .A(n654), .B(n883), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(KEYINPUT82), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n656), .A2(G868), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT83), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U735 ( .A1(G2090), .A2(n661), .ZN(n663) );
  XNOR2_X1 U736 ( .A(KEYINPUT84), .B(KEYINPUT21), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U738 ( .A1(G2072), .A2(n664), .ZN(G158) );
  XNOR2_X1 U739 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U741 ( .A1(G220), .A2(G219), .ZN(n665) );
  XNOR2_X1 U742 ( .A(KEYINPUT22), .B(n665), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n666), .A2(G96), .ZN(n667) );
  NOR2_X1 U744 ( .A1(n667), .A2(G218), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(KEYINPUT85), .ZN(n817) );
  NAND2_X1 U746 ( .A1(n817), .A2(G2106), .ZN(n672) );
  NAND2_X1 U747 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U748 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G108), .A2(n670), .ZN(n818) );
  NAND2_X1 U750 ( .A1(n818), .A2(G567), .ZN(n671) );
  NAND2_X1 U751 ( .A1(n672), .A2(n671), .ZN(n838) );
  NAND2_X1 U752 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U753 ( .A1(n838), .A2(n673), .ZN(n816) );
  NAND2_X1 U754 ( .A1(n816), .A2(G36), .ZN(G176) );
  INV_X1 U755 ( .A(G166), .ZN(G303) );
  NAND2_X1 U756 ( .A1(G160), .A2(G40), .ZN(n758) );
  INV_X1 U757 ( .A(n758), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n726), .A2(G8), .ZN(n791) );
  NOR2_X1 U759 ( .A1(G1976), .A2(G288), .ZN(n739) );
  NAND2_X1 U760 ( .A1(n739), .A2(KEYINPUT33), .ZN(n675) );
  NOR2_X1 U761 ( .A1(n791), .A2(n675), .ZN(n746) );
  NAND2_X1 U762 ( .A1(n693), .A2(G2072), .ZN(n676) );
  XNOR2_X1 U763 ( .A(n676), .B(KEYINPUT27), .ZN(n678) );
  XNOR2_X1 U764 ( .A(KEYINPUT95), .B(G1956), .ZN(n936) );
  NOR2_X1 U765 ( .A1(n936), .A2(n693), .ZN(n677) );
  NOR2_X1 U766 ( .A1(n678), .A2(n677), .ZN(n680) );
  INV_X1 U767 ( .A(G299), .ZN(n911) );
  NOR2_X1 U768 ( .A1(n680), .A2(n911), .ZN(n679) );
  NAND2_X1 U769 ( .A1(n680), .A2(n911), .ZN(n700) );
  NAND2_X1 U770 ( .A1(G1348), .A2(n918), .ZN(n681) );
  XNOR2_X1 U771 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n690) );
  NAND2_X1 U772 ( .A1(n681), .A2(n690), .ZN(n682) );
  NOR2_X1 U773 ( .A1(G1341), .A2(n682), .ZN(n683) );
  NOR2_X1 U774 ( .A1(n693), .A2(n683), .ZN(n684) );
  NOR2_X1 U775 ( .A1(n910), .A2(n684), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n918), .A2(G2067), .ZN(n686) );
  NAND2_X1 U777 ( .A1(G1996), .A2(n690), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U779 ( .A1(n687), .A2(n693), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(n692) );
  NOR2_X1 U781 ( .A1(G1996), .A2(n690), .ZN(n691) );
  NOR2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n698) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n726), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G2067), .A2(n693), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U786 ( .A1(n696), .A2(n918), .ZN(n697) );
  NOR2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U789 ( .A1(n511), .A2(n701), .ZN(n703) );
  XNOR2_X1 U790 ( .A(KEYINPUT97), .B(KEYINPUT29), .ZN(n702) );
  XNOR2_X1 U791 ( .A(n703), .B(n702), .ZN(n707) );
  XNOR2_X1 U792 ( .A(G2078), .B(KEYINPUT25), .ZN(n962) );
  NOR2_X1 U793 ( .A1(n726), .A2(n962), .ZN(n705) );
  AND2_X1 U794 ( .A1(n726), .A2(G1961), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n708) );
  NAND2_X1 U796 ( .A1(n708), .A2(G171), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n717) );
  OR2_X1 U798 ( .A1(G171), .A2(n708), .ZN(n714) );
  NOR2_X1 U799 ( .A1(G1966), .A2(n791), .ZN(n718) );
  NOR2_X1 U800 ( .A1(G2084), .A2(n726), .ZN(n721) );
  INV_X1 U801 ( .A(n721), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n709), .A2(G8), .ZN(n710) );
  XNOR2_X1 U803 ( .A(KEYINPUT30), .B(n711), .ZN(n712) );
  AND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U805 ( .A(KEYINPUT31), .B(n715), .Z(n716) );
  NAND2_X1 U806 ( .A1(n717), .A2(n716), .ZN(n725) );
  XNOR2_X1 U807 ( .A(n725), .B(KEYINPUT98), .ZN(n720) );
  INV_X1 U808 ( .A(n718), .ZN(n719) );
  AND2_X1 U809 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U810 ( .A1(G8), .A2(n721), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U812 ( .A(KEYINPUT99), .B(n724), .ZN(n736) );
  XOR2_X1 U813 ( .A(KEYINPUT100), .B(KEYINPUT32), .Z(n734) );
  NAND2_X1 U814 ( .A1(G286), .A2(n725), .ZN(n731) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n791), .ZN(n728) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n726), .ZN(n727) );
  NOR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n729), .A2(G303), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U820 ( .A1(G8), .A2(n732), .ZN(n733) );
  XNOR2_X1 U821 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U822 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U823 ( .A(n737), .B(KEYINPUT101), .ZN(n786) );
  NOR2_X1 U824 ( .A1(G1971), .A2(G303), .ZN(n738) );
  NOR2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n922) );
  INV_X1 U826 ( .A(KEYINPUT33), .ZN(n740) );
  AND2_X1 U827 ( .A1(n922), .A2(n740), .ZN(n741) );
  NAND2_X1 U828 ( .A1(n786), .A2(n741), .ZN(n744) );
  NAND2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n913) );
  INV_X1 U830 ( .A(n913), .ZN(n742) );
  OR2_X1 U831 ( .A1(KEYINPUT33), .A2(n513), .ZN(n743) );
  NAND2_X1 U832 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n746), .A2(n745), .ZN(n783) );
  XOR2_X1 U834 ( .A(G1981), .B(G305), .Z(n906) );
  NAND2_X1 U835 ( .A1(G104), .A2(n863), .ZN(n748) );
  NAND2_X1 U836 ( .A1(G140), .A2(n864), .ZN(n747) );
  NAND2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U838 ( .A(KEYINPUT34), .B(n749), .ZN(n755) );
  NAND2_X1 U839 ( .A1(n868), .A2(G128), .ZN(n750) );
  XOR2_X1 U840 ( .A(KEYINPUT89), .B(n750), .Z(n752) );
  NAND2_X1 U841 ( .A1(n867), .A2(G116), .ZN(n751) );
  NAND2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n753) );
  XOR2_X1 U843 ( .A(KEYINPUT35), .B(n753), .Z(n754) );
  NOR2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U845 ( .A(KEYINPUT36), .B(n756), .ZN(n880) );
  XNOR2_X1 U846 ( .A(KEYINPUT37), .B(G2067), .ZN(n806) );
  NOR2_X1 U847 ( .A1(n880), .A2(n806), .ZN(n995) );
  NOR2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U849 ( .A(n759), .B(KEYINPUT88), .Z(n779) );
  INV_X1 U850 ( .A(n779), .ZN(n808) );
  NAND2_X1 U851 ( .A1(n995), .A2(n808), .ZN(n804) );
  NAND2_X1 U852 ( .A1(n863), .A2(G105), .ZN(n760) );
  XNOR2_X1 U853 ( .A(n760), .B(KEYINPUT38), .ZN(n762) );
  NAND2_X1 U854 ( .A1(G129), .A2(n868), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G117), .A2(n867), .ZN(n763) );
  XNOR2_X1 U857 ( .A(KEYINPUT91), .B(n763), .ZN(n764) );
  NOR2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U859 ( .A(n766), .B(KEYINPUT92), .ZN(n768) );
  NAND2_X1 U860 ( .A1(G141), .A2(n864), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n874) );
  NAND2_X1 U862 ( .A1(G1996), .A2(n874), .ZN(n769) );
  XNOR2_X1 U863 ( .A(n769), .B(KEYINPUT93), .ZN(n778) );
  NAND2_X1 U864 ( .A1(G107), .A2(n867), .ZN(n771) );
  NAND2_X1 U865 ( .A1(G119), .A2(n868), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U867 ( .A1(n864), .A2(G131), .ZN(n772) );
  XOR2_X1 U868 ( .A(KEYINPUT90), .B(n772), .Z(n773) );
  NOR2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U870 ( .A1(n863), .A2(G95), .ZN(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n859) );
  AND2_X1 U872 ( .A1(G1991), .A2(n859), .ZN(n777) );
  NOR2_X1 U873 ( .A1(n778), .A2(n777), .ZN(n997) );
  NOR2_X1 U874 ( .A1(n779), .A2(n997), .ZN(n801) );
  INV_X1 U875 ( .A(n801), .ZN(n780) );
  NAND2_X1 U876 ( .A1(n804), .A2(n780), .ZN(n781) );
  XOR2_X1 U877 ( .A(n781), .B(KEYINPUT94), .Z(n793) );
  AND2_X1 U878 ( .A1(n906), .A2(n793), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n795) );
  NOR2_X1 U880 ( .A1(G2090), .A2(G303), .ZN(n784) );
  NAND2_X1 U881 ( .A1(G8), .A2(n784), .ZN(n785) );
  NAND2_X1 U882 ( .A1(n786), .A2(n785), .ZN(n788) );
  AND2_X1 U883 ( .A1(n791), .A2(n793), .ZN(n787) );
  NAND2_X1 U884 ( .A1(n788), .A2(n787), .ZN(n794) );
  NOR2_X1 U885 ( .A1(G1981), .A2(G305), .ZN(n789) );
  XOR2_X1 U886 ( .A(n789), .B(KEYINPUT24), .Z(n790) );
  NOR2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n795), .A2(n514), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n796), .B(KEYINPUT102), .ZN(n798) );
  XNOR2_X1 U890 ( .A(G1986), .B(G290), .ZN(n915) );
  NAND2_X1 U891 ( .A1(n915), .A2(n808), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n811) );
  NOR2_X1 U893 ( .A1(G1996), .A2(n874), .ZN(n983) );
  NOR2_X1 U894 ( .A1(G1991), .A2(n859), .ZN(n991) );
  NOR2_X1 U895 ( .A1(G1986), .A2(G290), .ZN(n799) );
  NOR2_X1 U896 ( .A1(n991), .A2(n799), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n802) );
  NOR2_X1 U898 ( .A1(n983), .A2(n802), .ZN(n803) );
  XNOR2_X1 U899 ( .A(KEYINPUT39), .B(n803), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n880), .A2(n806), .ZN(n988) );
  NAND2_X1 U902 ( .A1(n807), .A2(n988), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U905 ( .A(n812), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n813), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n814) );
  NAND2_X1 U908 ( .A1(G661), .A2(n814), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(G188) );
  NOR2_X1 U911 ( .A1(n818), .A2(n817), .ZN(G325) );
  XNOR2_X1 U912 ( .A(KEYINPUT103), .B(G325), .ZN(G261) );
  INV_X1 U914 ( .A(G120), .ZN(G236) );
  INV_X1 U915 ( .A(G96), .ZN(G221) );
  INV_X1 U916 ( .A(G69), .ZN(G235) );
  XOR2_X1 U917 ( .A(G2100), .B(KEYINPUT43), .Z(n820) );
  XNOR2_X1 U918 ( .A(G2090), .B(G2678), .ZN(n819) );
  XNOR2_X1 U919 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U920 ( .A(n821), .B(KEYINPUT104), .Z(n823) );
  XNOR2_X1 U921 ( .A(G2067), .B(G2072), .ZN(n822) );
  XNOR2_X1 U922 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U923 ( .A(KEYINPUT42), .B(G2096), .Z(n825) );
  XNOR2_X1 U924 ( .A(G2078), .B(G2084), .ZN(n824) );
  XNOR2_X1 U925 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n827), .B(n826), .ZN(G227) );
  XOR2_X1 U927 ( .A(G1981), .B(G1961), .Z(n829) );
  XNOR2_X1 U928 ( .A(G1986), .B(G1971), .ZN(n828) );
  XNOR2_X1 U929 ( .A(n829), .B(n828), .ZN(n833) );
  XOR2_X1 U930 ( .A(G1966), .B(G1956), .Z(n831) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1991), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U933 ( .A(n833), .B(n832), .Z(n835) );
  XNOR2_X1 U934 ( .A(G2474), .B(KEYINPUT41), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n837) );
  XOR2_X1 U936 ( .A(G1976), .B(KEYINPUT105), .Z(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(G229) );
  INV_X1 U938 ( .A(n838), .ZN(G319) );
  NAND2_X1 U939 ( .A1(G100), .A2(n863), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n839), .B(KEYINPUT108), .ZN(n848) );
  NAND2_X1 U941 ( .A1(G124), .A2(n868), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n840), .B(KEYINPUT44), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n841), .B(KEYINPUT106), .ZN(n843) );
  NAND2_X1 U944 ( .A1(G136), .A2(n864), .ZN(n842) );
  NAND2_X1 U945 ( .A1(n843), .A2(n842), .ZN(n846) );
  NAND2_X1 U946 ( .A1(G112), .A2(n867), .ZN(n844) );
  XNOR2_X1 U947 ( .A(KEYINPUT107), .B(n844), .ZN(n845) );
  NOR2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n847) );
  NAND2_X1 U949 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U950 ( .A(KEYINPUT109), .B(n849), .ZN(G162) );
  NAND2_X1 U951 ( .A1(G118), .A2(n867), .ZN(n851) );
  NAND2_X1 U952 ( .A1(G130), .A2(n868), .ZN(n850) );
  NAND2_X1 U953 ( .A1(n851), .A2(n850), .ZN(n856) );
  NAND2_X1 U954 ( .A1(G106), .A2(n863), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G142), .A2(n864), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n854) );
  XOR2_X1 U957 ( .A(n854), .B(KEYINPUT45), .Z(n855) );
  NOR2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U959 ( .A(KEYINPUT48), .B(n857), .Z(n858) );
  XOR2_X1 U960 ( .A(n858), .B(KEYINPUT46), .Z(n861) );
  XOR2_X1 U961 ( .A(n859), .B(KEYINPUT110), .Z(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n987), .B(n862), .ZN(n876) );
  NAND2_X1 U964 ( .A1(G103), .A2(n863), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G139), .A2(n864), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n873) );
  NAND2_X1 U967 ( .A1(G115), .A2(n867), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G127), .A2(n868), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  NOR2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n999) );
  XNOR2_X1 U972 ( .A(n874), .B(n999), .ZN(n875) );
  XNOR2_X1 U973 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U974 ( .A(n877), .B(G162), .Z(n879) );
  XNOR2_X1 U975 ( .A(G164), .B(G160), .ZN(n878) );
  XNOR2_X1 U976 ( .A(n879), .B(n878), .ZN(n881) );
  XNOR2_X1 U977 ( .A(n881), .B(n880), .ZN(n882) );
  NOR2_X1 U978 ( .A1(G37), .A2(n882), .ZN(G395) );
  XOR2_X1 U979 ( .A(KEYINPUT111), .B(n883), .Z(n886) );
  XNOR2_X1 U980 ( .A(G286), .B(n884), .ZN(n885) );
  XNOR2_X1 U981 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U982 ( .A(G171), .B(n887), .ZN(n888) );
  XNOR2_X1 U983 ( .A(n888), .B(n910), .ZN(n889) );
  NOR2_X1 U984 ( .A1(G37), .A2(n889), .ZN(G397) );
  NOR2_X1 U985 ( .A1(G227), .A2(G229), .ZN(n891) );
  XNOR2_X1 U986 ( .A(KEYINPUT112), .B(KEYINPUT49), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n902) );
  XOR2_X1 U988 ( .A(G2451), .B(G2430), .Z(n893) );
  XNOR2_X1 U989 ( .A(G2438), .B(G2443), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n899) );
  XOR2_X1 U991 ( .A(G2435), .B(G2454), .Z(n895) );
  XNOR2_X1 U992 ( .A(G1348), .B(G1341), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U994 ( .A(G2446), .B(G2427), .Z(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U996 ( .A(n899), .B(n898), .Z(n900) );
  NAND2_X1 U997 ( .A1(G14), .A2(n900), .ZN(n905) );
  NAND2_X1 U998 ( .A1(G319), .A2(n905), .ZN(n901) );
  NOR2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  INV_X1 U1004 ( .A(n905), .ZN(G401) );
  XNOR2_X1 U1005 ( .A(G168), .B(G1966), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1007 ( .A(KEYINPUT57), .B(n908), .Z(n931) );
  XOR2_X1 U1008 ( .A(G1341), .B(KEYINPUT121), .Z(n909) );
  XNOR2_X1 U1009 ( .A(n910), .B(n909), .ZN(n928) );
  XNOR2_X1 U1010 ( .A(n911), .B(G1956), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(G1971), .A2(G303), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n925) );
  XOR2_X1 U1015 ( .A(n918), .B(G1348), .Z(n920) );
  XNOR2_X1 U1016 ( .A(G171), .B(G1961), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(KEYINPUT119), .B(n921), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1021 ( .A(KEYINPUT120), .B(n926), .Z(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1023 ( .A(KEYINPUT122), .B(n929), .Z(n930) );
  NOR2_X1 U1024 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1025 ( .A(G16), .B(KEYINPUT56), .Z(n932) );
  NOR2_X1 U1026 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1027 ( .A(KEYINPUT123), .B(n934), .ZN(n1013) );
  XOR2_X1 U1028 ( .A(G16), .B(KEYINPUT124), .Z(n959) );
  XNOR2_X1 U1029 ( .A(KEYINPUT125), .B(G1966), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(n935), .B(G21), .ZN(n948) );
  XNOR2_X1 U1031 ( .A(G20), .B(n936), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(G6), .B(G1981), .ZN(n937) );
  NOR2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1036 ( .A(KEYINPUT59), .B(G1348), .Z(n941) );
  XNOR2_X1 U1037 ( .A(G4), .B(n941), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(KEYINPUT60), .B(n944), .Z(n946) );
  XNOR2_X1 U1040 ( .A(G1961), .B(G5), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n956) );
  XOR2_X1 U1043 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n954) );
  XOR2_X1 U1044 ( .A(G1986), .B(G24), .Z(n952) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G22), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G23), .B(G1976), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1049 ( .A(n954), .B(n953), .Z(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT61), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n960), .ZN(n1011) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n961), .ZN(n977) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n975) );
  XNOR2_X1 U1057 ( .A(G27), .B(n962), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G1996), .B(G32), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(KEYINPUT116), .B(n969), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(G28), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(G25), .B(G1991), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n978), .B(KEYINPUT118), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(KEYINPUT117), .B(n979), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(G29), .A2(n980), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n981), .B(KEYINPUT55), .ZN(n1009) );
  XOR2_X1 U1075 ( .A(G2090), .B(G162), .Z(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT51), .B(n984), .Z(n993) );
  XNOR2_X1 U1078 ( .A(G2084), .B(G160), .ZN(n985) );
  XNOR2_X1 U1079 ( .A(KEYINPUT113), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT114), .B(n998), .ZN(n1005) );
  XNOR2_X1 U1087 ( .A(G2072), .B(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(G164), .B(G2078), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(KEYINPUT50), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(KEYINPUT115), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1006), .Z(n1007) );
  NAND2_X1 U1094 ( .A1(G29), .A2(n1007), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(n1014), .B(KEYINPUT62), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(KEYINPUT127), .B(n1015), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

