

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G2104), .A2(G2105), .ZN(n553) );
  NOR2_X2 U549 ( .A1(G2104), .A2(n550), .ZN(n558) );
  XOR2_X1 U550 ( .A(n742), .B(KEYINPUT99), .Z(n514) );
  AND2_X1 U551 ( .A1(n745), .A2(n699), .ZN(n515) );
  INV_X1 U552 ( .A(G8), .ZN(n698) );
  NOR2_X1 U553 ( .A1(n774), .A2(G1966), .ZN(n696) );
  NOR2_X1 U554 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U555 ( .A1(n697), .A2(G8), .ZN(n774) );
  NOR2_X1 U556 ( .A1(n778), .A2(n777), .ZN(n798) );
  NOR2_X1 U557 ( .A1(G651), .A2(G543), .ZN(n640) );
  XNOR2_X1 U558 ( .A(KEYINPUT80), .B(KEYINPUT7), .ZN(n532) );
  XOR2_X1 U559 ( .A(KEYINPUT0), .B(G543), .Z(n637) );
  INV_X1 U560 ( .A(G651), .ZN(n522) );
  NOR2_X1 U561 ( .A1(n637), .A2(n522), .ZN(n641) );
  NAND2_X1 U562 ( .A1(n641), .A2(G76), .ZN(n516) );
  XNOR2_X1 U563 ( .A(KEYINPUT78), .B(n516), .ZN(n520) );
  XOR2_X1 U564 ( .A(KEYINPUT77), .B(KEYINPUT4), .Z(n518) );
  NAND2_X1 U565 ( .A1(G89), .A2(n640), .ZN(n517) );
  XNOR2_X1 U566 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U568 ( .A(n521), .B(KEYINPUT5), .ZN(n530) );
  XNOR2_X1 U569 ( .A(KEYINPUT79), .B(KEYINPUT6), .ZN(n528) );
  NOR2_X1 U570 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U571 ( .A(KEYINPUT1), .B(n523), .Z(n644) );
  NAND2_X1 U572 ( .A1(n644), .A2(G63), .ZN(n526) );
  NOR2_X1 U573 ( .A1(G651), .A2(n637), .ZN(n524) );
  XNOR2_X1 U574 ( .A(KEYINPUT66), .B(n524), .ZN(n645) );
  NAND2_X1 U575 ( .A1(G51), .A2(n645), .ZN(n525) );
  NAND2_X1 U576 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U577 ( .A(n528), .B(n527), .ZN(n529) );
  NAND2_X1 U578 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U579 ( .A(n532), .B(n531), .ZN(G168) );
  XOR2_X1 U580 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U581 ( .A1(G60), .A2(n644), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G85), .A2(n640), .ZN(n533) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U584 ( .A1(n641), .A2(G72), .ZN(n536) );
  NAND2_X1 U585 ( .A1(G47), .A2(n645), .ZN(n535) );
  NAND2_X1 U586 ( .A1(n536), .A2(n535), .ZN(n537) );
  OR2_X1 U587 ( .A1(n538), .A2(n537), .ZN(G290) );
  NAND2_X1 U588 ( .A1(G52), .A2(n645), .ZN(n539) );
  XNOR2_X1 U589 ( .A(n539), .B(KEYINPUT68), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G64), .A2(n644), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n547) );
  NAND2_X1 U592 ( .A1(G90), .A2(n640), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G77), .A2(n641), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U595 ( .A(KEYINPUT69), .B(n544), .ZN(n545) );
  XNOR2_X1 U596 ( .A(KEYINPUT9), .B(n545), .ZN(n546) );
  NOR2_X1 U597 ( .A1(n547), .A2(n546), .ZN(G171) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G57), .ZN(G237) );
  INV_X1 U600 ( .A(G132), .ZN(G219) );
  INV_X1 U601 ( .A(G82), .ZN(G220) );
  AND2_X1 U602 ( .A1(G2105), .A2(G2104), .ZN(n867) );
  NAND2_X1 U603 ( .A1(G113), .A2(n867), .ZN(n549) );
  INV_X1 U604 ( .A(G2105), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G125), .A2(n558), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n557) );
  NAND2_X1 U607 ( .A1(n550), .A2(G2104), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n551), .B(KEYINPUT67), .ZN(n603) );
  NAND2_X1 U609 ( .A1(G101), .A2(n603), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT23), .B(n552), .Z(n555) );
  XOR2_X2 U611 ( .A(KEYINPUT17), .B(n553), .Z(n870) );
  NAND2_X1 U612 ( .A1(n870), .A2(G137), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U614 ( .A1(n557), .A2(n556), .ZN(G160) );
  AND2_X1 U615 ( .A1(G138), .A2(n870), .ZN(n563) );
  NAND2_X1 U616 ( .A1(G114), .A2(n867), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G126), .A2(n558), .ZN(n559) );
  AND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U619 ( .A1(G102), .A2(n603), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(n675) );
  NOR2_X1 U621 ( .A1(n563), .A2(n675), .ZN(G164) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U623 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U624 ( .A(G223), .B(KEYINPUT72), .Z(n815) );
  NAND2_X1 U625 ( .A1(n815), .A2(G567), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT73), .ZN(n566) );
  XNOR2_X1 U627 ( .A(KEYINPUT11), .B(n566), .ZN(G234) );
  NAND2_X1 U628 ( .A1(n644), .A2(G56), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT14), .B(n567), .ZN(n574) );
  NAND2_X1 U630 ( .A1(G81), .A2(n640), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(KEYINPUT12), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT74), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G68), .A2(n641), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(n572), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U637 ( .A(n575), .B(KEYINPUT75), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G43), .A2(n645), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n968) );
  INV_X1 U640 ( .A(G860), .ZN(n623) );
  NOR2_X1 U641 ( .A1(n968), .A2(n623), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT76), .B(n578), .Z(G153) );
  INV_X1 U643 ( .A(G171), .ZN(G301) );
  NAND2_X1 U644 ( .A1(G868), .A2(G301), .ZN(n587) );
  NAND2_X1 U645 ( .A1(G66), .A2(n644), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G92), .A2(n640), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U648 ( .A1(n641), .A2(G79), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G54), .A2(n645), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U652 ( .A(KEYINPUT15), .B(n585), .Z(n971) );
  OR2_X1 U653 ( .A1(n971), .A2(G868), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G91), .A2(n640), .ZN(n589) );
  NAND2_X1 U656 ( .A1(G78), .A2(n641), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n589), .A2(n588), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G65), .A2(n644), .ZN(n590) );
  XNOR2_X1 U659 ( .A(n590), .B(KEYINPUT70), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G53), .A2(n645), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n973) );
  XNOR2_X1 U663 ( .A(n973), .B(KEYINPUT71), .ZN(G299) );
  XNOR2_X1 U664 ( .A(KEYINPUT81), .B(G868), .ZN(n595) );
  NOR2_X1 U665 ( .A1(G286), .A2(n595), .ZN(n597) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(G297) );
  NAND2_X1 U668 ( .A1(n623), .A2(G559), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n598), .A2(n971), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U671 ( .A1(G868), .A2(n968), .ZN(n602) );
  NAND2_X1 U672 ( .A1(G868), .A2(n971), .ZN(n600) );
  NOR2_X1 U673 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U674 ( .A1(n602), .A2(n601), .ZN(G282) );
  XNOR2_X1 U675 ( .A(G2100), .B(KEYINPUT83), .ZN(n614) );
  NAND2_X1 U676 ( .A1(G111), .A2(n867), .ZN(n606) );
  INV_X1 U677 ( .A(n603), .ZN(n604) );
  INV_X1 U678 ( .A(n604), .ZN(n871) );
  NAND2_X1 U679 ( .A1(G99), .A2(n871), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U681 ( .A(KEYINPUT82), .B(n607), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n558), .A2(G123), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G135), .A2(n870), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n912) );
  XNOR2_X1 U687 ( .A(n912), .B(G2096), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U689 ( .A1(G93), .A2(n640), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G80), .A2(n641), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G67), .A2(n644), .ZN(n617) );
  XNOR2_X1 U693 ( .A(n617), .B(KEYINPUT84), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G55), .A2(n645), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  OR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n658) );
  NAND2_X1 U697 ( .A1(G559), .A2(n971), .ZN(n622) );
  XOR2_X1 U698 ( .A(n968), .B(n622), .Z(n656) );
  NAND2_X1 U699 ( .A1(n623), .A2(n656), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n624), .B(KEYINPUT85), .ZN(n625) );
  XOR2_X1 U701 ( .A(n658), .B(n625), .Z(G145) );
  XOR2_X1 U702 ( .A(KEYINPUT86), .B(KEYINPUT2), .Z(n627) );
  NAND2_X1 U703 ( .A1(G73), .A2(n641), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n627), .B(n626), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G61), .A2(n644), .ZN(n629) );
  NAND2_X1 U706 ( .A1(G86), .A2(n640), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G48), .A2(n645), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U711 ( .A1(G651), .A2(G74), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G49), .A2(n645), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U714 ( .A1(n644), .A2(n636), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G88), .A2(n640), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G75), .A2(n641), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n649) );
  NAND2_X1 U720 ( .A1(n644), .A2(G62), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G50), .A2(n645), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U723 ( .A1(n649), .A2(n648), .ZN(G166) );
  INV_X1 U724 ( .A(G166), .ZN(G303) );
  XOR2_X1 U725 ( .A(n658), .B(G305), .Z(n650) );
  XNOR2_X1 U726 ( .A(n650), .B(G299), .ZN(n651) );
  XNOR2_X1 U727 ( .A(KEYINPUT87), .B(n651), .ZN(n653) );
  XNOR2_X1 U728 ( .A(G288), .B(KEYINPUT19), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U730 ( .A(n654), .B(G303), .ZN(n655) );
  XNOR2_X1 U731 ( .A(n655), .B(G290), .ZN(n885) );
  XNOR2_X1 U732 ( .A(n656), .B(n885), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(G868), .ZN(n661) );
  INV_X1 U734 ( .A(G868), .ZN(n659) );
  NAND2_X1 U735 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U736 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n662) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U745 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U746 ( .A1(G96), .A2(n668), .ZN(n819) );
  NAND2_X1 U747 ( .A1(n819), .A2(G2106), .ZN(n672) );
  NAND2_X1 U748 ( .A1(G120), .A2(G108), .ZN(n669) );
  NOR2_X1 U749 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G69), .A2(n670), .ZN(n820) );
  NAND2_X1 U751 ( .A1(n820), .A2(G567), .ZN(n671) );
  NAND2_X1 U752 ( .A1(n672), .A2(n671), .ZN(n821) );
  NAND2_X1 U753 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U754 ( .A1(n821), .A2(n673), .ZN(n818) );
  NAND2_X1 U755 ( .A1(n818), .A2(G36), .ZN(G176) );
  INV_X1 U756 ( .A(G1384), .ZN(n676) );
  AND2_X1 U757 ( .A1(G138), .A2(n676), .ZN(n674) );
  NAND2_X1 U758 ( .A1(n870), .A2(n674), .ZN(n678) );
  NAND2_X1 U759 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U761 ( .A(KEYINPUT65), .B(n679), .Z(n691) );
  NAND2_X1 U762 ( .A1(G160), .A2(G40), .ZN(n693) );
  NOR2_X1 U763 ( .A1(n691), .A2(n693), .ZN(n810) );
  XNOR2_X1 U764 ( .A(G2067), .B(KEYINPUT37), .ZN(n807) );
  XNOR2_X1 U765 ( .A(KEYINPUT88), .B(KEYINPUT34), .ZN(n683) );
  NAND2_X1 U766 ( .A1(G140), .A2(n870), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G104), .A2(n871), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U769 ( .A(n683), .B(n682), .ZN(n689) );
  NAND2_X1 U770 ( .A1(n558), .A2(G128), .ZN(n684) );
  XOR2_X1 U771 ( .A(KEYINPUT89), .B(n684), .Z(n686) );
  NAND2_X1 U772 ( .A1(n867), .A2(G116), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U774 ( .A(KEYINPUT35), .B(n687), .Z(n688) );
  NOR2_X1 U775 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U776 ( .A(KEYINPUT36), .B(n690), .ZN(n882) );
  NOR2_X1 U777 ( .A1(n807), .A2(n882), .ZN(n914) );
  NAND2_X1 U778 ( .A1(n810), .A2(n914), .ZN(n805) );
  INV_X1 U779 ( .A(n805), .ZN(n778) );
  INV_X1 U780 ( .A(KEYINPUT64), .ZN(n695) );
  INV_X1 U781 ( .A(n691), .ZN(n692) );
  XNOR2_X1 U782 ( .A(n695), .B(n694), .ZN(n697) );
  XNOR2_X1 U783 ( .A(n696), .B(KEYINPUT93), .ZN(n745) );
  INV_X1 U784 ( .A(n697), .ZN(n718) );
  INV_X1 U785 ( .A(n718), .ZN(n736) );
  NOR2_X1 U786 ( .A1(n736), .A2(G2084), .ZN(n744) );
  NOR2_X1 U787 ( .A1(n744), .A2(n698), .ZN(n699) );
  XOR2_X1 U788 ( .A(KEYINPUT30), .B(n515), .Z(n700) );
  NOR2_X1 U789 ( .A1(G168), .A2(n700), .ZN(n701) );
  XNOR2_X1 U790 ( .A(n701), .B(KEYINPUT97), .ZN(n706) );
  XNOR2_X1 U791 ( .A(G1961), .B(KEYINPUT94), .ZN(n993) );
  NOR2_X1 U792 ( .A1(n718), .A2(n993), .ZN(n703) );
  XOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .Z(n941) );
  NOR2_X1 U794 ( .A1(n736), .A2(n941), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U796 ( .A(KEYINPUT95), .B(n704), .ZN(n731) );
  OR2_X1 U797 ( .A1(n731), .A2(G171), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U799 ( .A(n707), .B(KEYINPUT31), .ZN(n735) );
  NAND2_X1 U800 ( .A1(G2072), .A2(n718), .ZN(n708) );
  XNOR2_X1 U801 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  AND2_X1 U802 ( .A1(n736), .A2(G1956), .ZN(n709) );
  NOR2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n712) );
  NOR2_X1 U804 ( .A1(n973), .A2(n712), .ZN(n711) );
  XOR2_X1 U805 ( .A(n711), .B(KEYINPUT28), .Z(n729) );
  NAND2_X1 U806 ( .A1(n973), .A2(n712), .ZN(n727) );
  NAND2_X1 U807 ( .A1(n718), .A2(G1996), .ZN(n713) );
  XNOR2_X1 U808 ( .A(n713), .B(KEYINPUT26), .ZN(n715) );
  NAND2_X1 U809 ( .A1(n736), .A2(G1341), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U811 ( .A1(n968), .A2(n716), .ZN(n717) );
  OR2_X1 U812 ( .A1(n971), .A2(n717), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n971), .A2(n717), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n718), .A2(G2067), .ZN(n719) );
  XNOR2_X1 U815 ( .A(n719), .B(KEYINPUT96), .ZN(n721) );
  NAND2_X1 U816 ( .A1(n736), .A2(G1348), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U818 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U822 ( .A(KEYINPUT29), .B(n730), .Z(n733) );
  NAND2_X1 U823 ( .A1(G171), .A2(n731), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n746), .A2(G286), .ZN(n741) );
  NOR2_X1 U827 ( .A1(n736), .A2(G2090), .ZN(n738) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n774), .ZN(n737) );
  NOR2_X1 U829 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U830 ( .A1(n739), .A2(G303), .ZN(n740) );
  NAND2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(G8), .A2(n514), .ZN(n743) );
  XNOR2_X1 U833 ( .A(n743), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U834 ( .A1(G8), .A2(n744), .ZN(n750) );
  INV_X1 U835 ( .A(n745), .ZN(n748) );
  XOR2_X1 U836 ( .A(n746), .B(KEYINPUT98), .Z(n747) );
  NOR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n767) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n972), .A2(n753), .ZN(n755) );
  INV_X1 U843 ( .A(KEYINPUT33), .ZN(n754) );
  AND2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n767), .A2(n756), .ZN(n764) );
  NAND2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n966) );
  INV_X1 U847 ( .A(n966), .ZN(n757) );
  NOR2_X1 U848 ( .A1(n774), .A2(n757), .ZN(n758) );
  NOR2_X1 U849 ( .A1(KEYINPUT33), .A2(n758), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n972), .A2(KEYINPUT33), .ZN(n759) );
  OR2_X1 U851 ( .A1(n759), .A2(n774), .ZN(n760) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n978) );
  NAND2_X1 U853 ( .A1(n760), .A2(n978), .ZN(n761) );
  NOR2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n770) );
  NOR2_X1 U856 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U857 ( .A1(G8), .A2(n765), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n768), .A2(n774), .ZN(n769) );
  NAND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n776) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XOR2_X1 U862 ( .A(n771), .B(KEYINPUT92), .Z(n772) );
  XNOR2_X1 U863 ( .A(KEYINPUT24), .B(n772), .ZN(n773) );
  NOR2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U866 ( .A1(G131), .A2(n870), .ZN(n780) );
  NAND2_X1 U867 ( .A1(G95), .A2(n871), .ZN(n779) );
  NAND2_X1 U868 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U869 ( .A(KEYINPUT90), .B(n781), .ZN(n785) );
  NAND2_X1 U870 ( .A1(G107), .A2(n867), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G119), .A2(n558), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n851) );
  INV_X1 U874 ( .A(G1991), .ZN(n937) );
  NOR2_X1 U875 ( .A1(n851), .A2(n937), .ZN(n795) );
  NAND2_X1 U876 ( .A1(G117), .A2(n867), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G129), .A2(n558), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U879 ( .A(n788), .B(KEYINPUT91), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G141), .A2(n870), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n871), .A2(G105), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n850) );
  INV_X1 U885 ( .A(G1996), .ZN(n938) );
  NOR2_X1 U886 ( .A1(n850), .A2(n938), .ZN(n794) );
  NOR2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n910) );
  XOR2_X1 U888 ( .A(G1986), .B(G290), .Z(n961) );
  NAND2_X1 U889 ( .A1(n910), .A2(n961), .ZN(n796) );
  NAND2_X1 U890 ( .A1(n796), .A2(n810), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n813) );
  AND2_X1 U892 ( .A1(n938), .A2(n850), .ZN(n925) );
  INV_X1 U893 ( .A(n910), .ZN(n802) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n799) );
  AND2_X1 U895 ( .A1(n937), .A2(n851), .ZN(n913) );
  NOR2_X1 U896 ( .A1(n799), .A2(n913), .ZN(n800) );
  XNOR2_X1 U897 ( .A(n800), .B(KEYINPUT100), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U899 ( .A1(n925), .A2(n803), .ZN(n804) );
  XNOR2_X1 U900 ( .A(n804), .B(KEYINPUT39), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n807), .A2(n882), .ZN(n909) );
  NAND2_X1 U903 ( .A1(n808), .A2(n909), .ZN(n809) );
  XOR2_X1 U904 ( .A(KEYINPUT101), .B(n809), .Z(n811) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U907 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n815), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n816) );
  NAND2_X1 U910 ( .A1(G661), .A2(n816), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(G188) );
  XOR2_X1 U913 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U915 ( .A(G120), .ZN(G236) );
  INV_X1 U916 ( .A(G96), .ZN(G221) );
  NOR2_X1 U917 ( .A1(n820), .A2(n819), .ZN(G325) );
  INV_X1 U918 ( .A(G325), .ZN(G261) );
  INV_X1 U919 ( .A(n821), .ZN(G319) );
  XOR2_X1 U920 ( .A(G2474), .B(G1976), .Z(n823) );
  XNOR2_X1 U921 ( .A(G1966), .B(G1956), .ZN(n822) );
  XNOR2_X1 U922 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U923 ( .A(n824), .B(KEYINPUT105), .Z(n826) );
  XNOR2_X1 U924 ( .A(G1996), .B(G1991), .ZN(n825) );
  XNOR2_X1 U925 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U926 ( .A(G1986), .B(G1981), .Z(n828) );
  XNOR2_X1 U927 ( .A(G1961), .B(G1971), .ZN(n827) );
  XNOR2_X1 U928 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U929 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U930 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n831) );
  XNOR2_X1 U931 ( .A(n832), .B(n831), .ZN(G229) );
  XOR2_X1 U932 ( .A(G2100), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U933 ( .A(G2090), .B(G2678), .ZN(n833) );
  XNOR2_X1 U934 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U935 ( .A(n835), .B(KEYINPUT104), .Z(n837) );
  XNOR2_X1 U936 ( .A(G2072), .B(G2067), .ZN(n836) );
  XNOR2_X1 U937 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U938 ( .A(KEYINPUT42), .B(G2096), .Z(n839) );
  XNOR2_X1 U939 ( .A(G2084), .B(G2078), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(G227) );
  NAND2_X1 U942 ( .A1(G124), .A2(n558), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n842), .B(KEYINPUT44), .ZN(n845) );
  NAND2_X1 U944 ( .A1(G112), .A2(n867), .ZN(n843) );
  XOR2_X1 U945 ( .A(KEYINPUT107), .B(n843), .Z(n844) );
  NAND2_X1 U946 ( .A1(n845), .A2(n844), .ZN(n849) );
  NAND2_X1 U947 ( .A1(G136), .A2(n870), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G100), .A2(n871), .ZN(n846) );
  NAND2_X1 U949 ( .A1(n847), .A2(n846), .ZN(n848) );
  NOR2_X1 U950 ( .A1(n849), .A2(n848), .ZN(G162) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n852), .B(n912), .ZN(n857) );
  XOR2_X1 U953 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n854) );
  XNOR2_X1 U954 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(G164), .B(n855), .Z(n856) );
  XOR2_X1 U957 ( .A(n857), .B(n856), .Z(n881) );
  NAND2_X1 U958 ( .A1(G139), .A2(n870), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G103), .A2(n871), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n865) );
  NAND2_X1 U961 ( .A1(n558), .A2(G127), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT108), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G115), .A2(n867), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n863), .Z(n864) );
  NOR2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U967 ( .A(KEYINPUT109), .B(n866), .Z(n918) );
  XNOR2_X1 U968 ( .A(G160), .B(G162), .ZN(n878) );
  NAND2_X1 U969 ( .A1(G118), .A2(n867), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G130), .A2(n558), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G142), .A2(n870), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G106), .A2(n871), .ZN(n872) );
  NAND2_X1 U974 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n918), .B(n879), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n881), .B(n880), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n884) );
  NOR2_X1 U981 ( .A1(G37), .A2(n884), .ZN(G395) );
  XOR2_X1 U982 ( .A(KEYINPUT112), .B(n885), .Z(n887) );
  XNOR2_X1 U983 ( .A(G171), .B(n971), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  XOR2_X1 U985 ( .A(n888), .B(n968), .Z(n889) );
  XNOR2_X1 U986 ( .A(G286), .B(n889), .ZN(n890) );
  NOR2_X1 U987 ( .A1(G37), .A2(n890), .ZN(G397) );
  XNOR2_X1 U988 ( .A(G2446), .B(KEYINPUT102), .ZN(n900) );
  XOR2_X1 U989 ( .A(G2430), .B(G2427), .Z(n892) );
  XNOR2_X1 U990 ( .A(KEYINPUT103), .B(G2438), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U992 ( .A(G2435), .B(G2454), .Z(n894) );
  XNOR2_X1 U993 ( .A(G1341), .B(G1348), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U996 ( .A(G2443), .B(G2451), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n901), .A2(G14), .ZN(n908) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n908), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n902) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n902), .Z(n903) );
  XNOR2_X1 U1003 ( .A(n903), .B(KEYINPUT113), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G69), .ZN(G235) );
  INV_X1 U1009 ( .A(n908), .ZN(G401) );
  NAND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n932) );
  XOR2_X1 U1011 ( .A(G2084), .B(G160), .Z(n911) );
  NOR2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT115), .B(n917), .ZN(n930) );
  XNOR2_X1 U1016 ( .A(G2072), .B(n918), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(G164), .B(G2078), .ZN(n919) );
  XNOR2_X1 U1018 ( .A(n919), .B(KEYINPUT116), .ZN(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n922), .B(KEYINPUT50), .ZN(n923) );
  XOR2_X1 U1021 ( .A(KEYINPUT117), .B(n923), .Z(n928) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n926), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n933), .ZN(n935) );
  INV_X1 U1029 ( .A(KEYINPUT55), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n936), .A2(G29), .ZN(n1019) );
  XOR2_X1 U1032 ( .A(G2090), .B(G35), .Z(n953) );
  XNOR2_X1 U1033 ( .A(n937), .B(G25), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(n938), .B(G32), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(G27), .B(n941), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n949) );
  XOR2_X1 U1038 ( .A(G2067), .B(G26), .Z(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(G28), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(KEYINPUT118), .B(G2072), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G33), .B(n945), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1044 ( .A(KEYINPUT119), .B(n950), .Z(n951) );
  XNOR2_X1 U1045 ( .A(n951), .B(KEYINPUT53), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1047 ( .A(G34), .B(G2084), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(n954), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(n957), .Z(n958) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n958), .ZN(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT120), .B(n959), .Z(n960) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n960), .ZN(n1017) );
  XNOR2_X1 U1054 ( .A(G16), .B(KEYINPUT56), .ZN(n986) );
  XNOR2_X1 U1055 ( .A(G171), .B(G1961), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1057 ( .A(G1971), .B(G166), .Z(n963) );
  XNOR2_X1 U1058 ( .A(KEYINPUT122), .B(n963), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(G1341), .B(n968), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n984) );
  XNOR2_X1 U1063 ( .A(n971), .B(G1348), .ZN(n977) );
  XOR2_X1 U1064 ( .A(n972), .B(KEYINPUT121), .Z(n975) );
  XOR2_X1 U1065 ( .A(n973), .B(G1956), .Z(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n982) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G168), .ZN(n979) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT57), .B(n980), .Z(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n1015) );
  INV_X1 U1074 ( .A(G16), .ZN(n1013) );
  XNOR2_X1 U1075 ( .A(G1986), .B(G24), .ZN(n991) );
  XNOR2_X1 U1076 ( .A(G1971), .B(G22), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(G1976), .B(G23), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n989), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(KEYINPUT58), .B(n992), .ZN(n1006) );
  XNOR2_X1 U1082 ( .A(n993), .B(G5), .ZN(n1004) );
  XNOR2_X1 U1083 ( .A(KEYINPUT59), .B(G1348), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n994), .B(G4), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G20), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G1981), .B(G6), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT123), .B(n997), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT60), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(G1966), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(G21), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT126), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(KEYINPUT61), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1020), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

