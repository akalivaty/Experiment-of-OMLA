

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U551 ( .A1(n562), .A2(G2104), .ZN(n890) );
  NOR2_X1 U552 ( .A1(n709), .A2(n782), .ZN(n734) );
  NAND2_X1 U553 ( .A1(G8), .A2(n753), .ZN(n823) );
  AND2_X1 U554 ( .A1(n820), .A2(n819), .ZN(n827) );
  NAND2_X1 U555 ( .A1(n545), .A2(n546), .ZN(n753) );
  NOR2_X2 U556 ( .A1(n782), .A2(G1384), .ZN(n545) );
  INV_X1 U557 ( .A(G1341), .ZN(n538) );
  NAND2_X1 U558 ( .A1(n544), .A2(n545), .ZN(n543) );
  OR2_X1 U559 ( .A1(G164), .A2(G1384), .ZN(n709) );
  INV_X1 U560 ( .A(KEYINPUT104), .ZN(n524) );
  NAND2_X1 U561 ( .A1(n536), .A2(n562), .ZN(n535) );
  INV_X1 U562 ( .A(G2104), .ZN(n536) );
  AND2_X1 U563 ( .A1(n543), .A2(n541), .ZN(n540) );
  NOR2_X1 U564 ( .A1(n539), .A2(n519), .ZN(n537) );
  NOR2_X1 U565 ( .A1(n719), .A2(n718), .ZN(n720) );
  AND2_X1 U566 ( .A1(n527), .A2(n526), .ZN(n529) );
  INV_X1 U567 ( .A(G2105), .ZN(n562) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n562), .ZN(n895) );
  NOR2_X1 U569 ( .A1(n781), .A2(n780), .ZN(n814) );
  NOR2_X1 U570 ( .A1(n827), .A2(n826), .ZN(n828) );
  AND2_X1 U571 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U572 ( .A1(n707), .A2(n706), .ZN(G160) );
  AND2_X1 U573 ( .A1(n757), .A2(n524), .ZN(n515) );
  AND2_X1 U574 ( .A1(G286), .A2(KEYINPUT104), .ZN(n516) );
  AND2_X1 U575 ( .A1(n752), .A2(n751), .ZN(n517) );
  AND2_X1 U576 ( .A1(n531), .A2(n515), .ZN(n518) );
  AND2_X1 U577 ( .A1(n547), .A2(n538), .ZN(n519) );
  INV_X1 U578 ( .A(KEYINPUT98), .ZN(n547) );
  NAND2_X1 U579 ( .A1(n530), .A2(KEYINPUT104), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n520), .A2(n731), .ZN(n733) );
  XNOR2_X1 U581 ( .A(n522), .B(n521), .ZN(n520) );
  INV_X1 U582 ( .A(KEYINPUT100), .ZN(n521) );
  NAND2_X1 U583 ( .A1(n523), .A2(n727), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n726), .A2(n725), .ZN(n523) );
  NAND2_X1 U585 ( .A1(n531), .A2(n757), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n525), .A2(n518), .ZN(n528) );
  NAND2_X1 U587 ( .A1(n533), .A2(G286), .ZN(n525) );
  INV_X1 U588 ( .A(n752), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n533), .A2(n516), .ZN(n527) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n758) );
  NAND2_X1 U591 ( .A1(n532), .A2(G286), .ZN(n531) );
  INV_X1 U592 ( .A(n751), .ZN(n532) );
  XNOR2_X1 U593 ( .A(n534), .B(KEYINPUT89), .ZN(n566) );
  NAND2_X1 U594 ( .A1(n891), .A2(G138), .ZN(n534) );
  XNOR2_X2 U595 ( .A(n535), .B(KEYINPUT17), .ZN(n891) );
  INV_X1 U596 ( .A(G164), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n540), .A2(n537), .ZN(n713) );
  NOR2_X1 U598 ( .A1(n546), .A2(n542), .ZN(n539) );
  OR2_X1 U599 ( .A1(n545), .A2(n542), .ZN(n541) );
  NAND2_X1 U600 ( .A1(KEYINPUT98), .A2(G1341), .ZN(n542) );
  NOR2_X1 U601 ( .A1(G164), .A2(KEYINPUT98), .ZN(n544) );
  INV_X1 U602 ( .A(KEYINPUT107), .ZN(n776) );
  XNOR2_X1 U603 ( .A(n777), .B(n776), .ZN(n781) );
  NOR2_X1 U604 ( .A1(n657), .A2(G651), .ZN(n660) );
  INV_X1 U605 ( .A(G651), .ZN(n553) );
  NOR2_X1 U606 ( .A1(G543), .A2(n553), .ZN(n548) );
  XOR2_X1 U607 ( .A(KEYINPUT1), .B(n548), .Z(n663) );
  NAND2_X1 U608 ( .A1(G63), .A2(n663), .ZN(n550) );
  XOR2_X1 U609 ( .A(KEYINPUT0), .B(G543), .Z(n657) );
  NAND2_X1 U610 ( .A1(G51), .A2(n660), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(n551), .ZN(n558) );
  NOR2_X1 U613 ( .A1(G543), .A2(G651), .ZN(n662) );
  NAND2_X1 U614 ( .A1(n662), .A2(G89), .ZN(n552) );
  XNOR2_X1 U615 ( .A(n552), .B(KEYINPUT4), .ZN(n555) );
  NOR2_X1 U616 ( .A1(n657), .A2(n553), .ZN(n666) );
  NAND2_X1 U617 ( .A1(G76), .A2(n666), .ZN(n554) );
  NAND2_X1 U618 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U619 ( .A(n556), .B(KEYINPUT5), .Z(n557) );
  NOR2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT73), .B(n559), .Z(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT7), .B(n560), .Z(G168) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U624 ( .A1(n890), .A2(G102), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT88), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G126), .A2(n895), .ZN(n564) );
  AND2_X1 U627 ( .A1(G2104), .A2(G2105), .ZN(n894) );
  NAND2_X1 U628 ( .A1(G114), .A2(n894), .ZN(n563) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X2 U631 ( .A(KEYINPUT90), .B(n569), .ZN(G164) );
  NAND2_X1 U632 ( .A1(G85), .A2(n662), .ZN(n571) );
  NAND2_X1 U633 ( .A1(G72), .A2(n666), .ZN(n570) );
  NAND2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G60), .A2(n663), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G47), .A2(n660), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  OR2_X1 U638 ( .A1(n575), .A2(n574), .ZN(G290) );
  NAND2_X1 U639 ( .A1(G64), .A2(n663), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G52), .A2(n660), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n584) );
  XNOR2_X1 U642 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n666), .A2(G77), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n662), .A2(G90), .ZN(n578) );
  XOR2_X1 U645 ( .A(KEYINPUT65), .B(n578), .Z(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(n582), .B(n581), .Z(n583) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(G171) );
  AND2_X1 U649 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U650 ( .A1(G123), .A2(n895), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n585), .B(KEYINPUT18), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n586), .B(KEYINPUT76), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G135), .A2(n891), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(KEYINPUT77), .B(n589), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G99), .A2(n890), .ZN(n591) );
  NAND2_X1 U657 ( .A1(G111), .A2(n894), .ZN(n590) );
  AND2_X1 U658 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n970) );
  XNOR2_X1 U660 ( .A(G2096), .B(n970), .ZN(n594) );
  OR2_X1 U661 ( .A1(G2100), .A2(n594), .ZN(G156) );
  INV_X1 U662 ( .A(G57), .ZN(G237) );
  INV_X1 U663 ( .A(G132), .ZN(G219) );
  INV_X1 U664 ( .A(G82), .ZN(G220) );
  NAND2_X1 U665 ( .A1(G62), .A2(n663), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G50), .A2(n660), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n597), .B(KEYINPUT81), .ZN(n599) );
  NAND2_X1 U669 ( .A1(G75), .A2(n666), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n662), .A2(G88), .ZN(n600) );
  XOR2_X1 U672 ( .A(KEYINPUT82), .B(n600), .Z(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G166) );
  NAND2_X1 U674 ( .A1(G7), .A2(G661), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT10), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT68), .B(n604), .Z(n847) );
  NAND2_X1 U677 ( .A1(n847), .A2(G567), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT69), .ZN(n606) );
  XNOR2_X1 U679 ( .A(KEYINPUT11), .B(n606), .ZN(G234) );
  NAND2_X1 U680 ( .A1(n663), .A2(G56), .ZN(n607) );
  XOR2_X1 U681 ( .A(KEYINPUT14), .B(n607), .Z(n613) );
  NAND2_X1 U682 ( .A1(n662), .A2(G81), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U684 ( .A1(G68), .A2(n666), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT13), .B(n611), .Z(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT70), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G43), .A2(n660), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n1003) );
  INV_X1 U691 ( .A(G860), .ZN(n637) );
  OR2_X1 U692 ( .A1(n1003), .A2(n637), .ZN(G153) );
  XNOR2_X1 U693 ( .A(G171), .B(KEYINPUT71), .ZN(G301) );
  NAND2_X1 U694 ( .A1(G868), .A2(G301), .ZN(n626) );
  NAND2_X1 U695 ( .A1(G79), .A2(n666), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G54), .A2(n660), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G92), .A2(n662), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G66), .A2(n663), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U701 ( .A(KEYINPUT72), .B(n621), .ZN(n622) );
  NOR2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U703 ( .A(n624), .B(KEYINPUT15), .Z(n1000) );
  INV_X1 U704 ( .A(n1000), .ZN(n719) );
  INV_X1 U705 ( .A(G868), .ZN(n682) );
  NAND2_X1 U706 ( .A1(n719), .A2(n682), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(G284) );
  NAND2_X1 U708 ( .A1(G78), .A2(n666), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G65), .A2(n663), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G91), .A2(n662), .ZN(n629) );
  XNOR2_X1 U712 ( .A(KEYINPUT67), .B(n629), .ZN(n630) );
  NOR2_X1 U713 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n660), .A2(G53), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(G299) );
  NOR2_X1 U716 ( .A1(G286), .A2(n682), .ZN(n634) );
  XNOR2_X1 U717 ( .A(n634), .B(KEYINPUT74), .ZN(n636) );
  NOR2_X1 U718 ( .A1(G299), .A2(G868), .ZN(n635) );
  NOR2_X1 U719 ( .A1(n636), .A2(n635), .ZN(G297) );
  NAND2_X1 U720 ( .A1(n637), .A2(G559), .ZN(n638) );
  NAND2_X1 U721 ( .A1(n638), .A2(n1000), .ZN(n639) );
  XNOR2_X1 U722 ( .A(n639), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U723 ( .A1(G868), .A2(n1003), .ZN(n640) );
  XOR2_X1 U724 ( .A(KEYINPUT75), .B(n640), .Z(n643) );
  NAND2_X1 U725 ( .A1(G868), .A2(n1000), .ZN(n641) );
  NOR2_X1 U726 ( .A1(G559), .A2(n641), .ZN(n642) );
  NOR2_X1 U727 ( .A1(n643), .A2(n642), .ZN(G282) );
  NAND2_X1 U728 ( .A1(G559), .A2(n1000), .ZN(n644) );
  XNOR2_X1 U729 ( .A(n644), .B(n1003), .ZN(n679) );
  XNOR2_X1 U730 ( .A(KEYINPUT78), .B(n679), .ZN(n645) );
  NOR2_X1 U731 ( .A1(G860), .A2(n645), .ZN(n653) );
  NAND2_X1 U732 ( .A1(G93), .A2(n662), .ZN(n647) );
  NAND2_X1 U733 ( .A1(G80), .A2(n666), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U735 ( .A1(G55), .A2(n660), .ZN(n648) );
  XNOR2_X1 U736 ( .A(KEYINPUT79), .B(n648), .ZN(n649) );
  NOR2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U738 ( .A1(n663), .A2(G67), .ZN(n651) );
  NAND2_X1 U739 ( .A1(n652), .A2(n651), .ZN(n681) );
  XOR2_X1 U740 ( .A(n653), .B(n681), .Z(G145) );
  NAND2_X1 U741 ( .A1(G49), .A2(n660), .ZN(n655) );
  NAND2_X1 U742 ( .A1(G74), .A2(G651), .ZN(n654) );
  NAND2_X1 U743 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U744 ( .A1(n663), .A2(n656), .ZN(n659) );
  NAND2_X1 U745 ( .A1(n657), .A2(G87), .ZN(n658) );
  NAND2_X1 U746 ( .A1(n659), .A2(n658), .ZN(G288) );
  NAND2_X1 U747 ( .A1(G48), .A2(n660), .ZN(n661) );
  XNOR2_X1 U748 ( .A(n661), .B(KEYINPUT80), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G86), .A2(n662), .ZN(n665) );
  NAND2_X1 U750 ( .A1(G61), .A2(n663), .ZN(n664) );
  NAND2_X1 U751 ( .A1(n665), .A2(n664), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n666), .A2(G73), .ZN(n667) );
  XOR2_X1 U753 ( .A(KEYINPUT2), .B(n667), .Z(n668) );
  NOR2_X1 U754 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n671), .A2(n670), .ZN(G305) );
  XNOR2_X1 U756 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n673) );
  XNOR2_X1 U757 ( .A(G288), .B(KEYINPUT19), .ZN(n672) );
  XNOR2_X1 U758 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U759 ( .A(G166), .B(n674), .ZN(n676) );
  XOR2_X1 U760 ( .A(G290), .B(G299), .Z(n675) );
  XNOR2_X1 U761 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U762 ( .A(n677), .B(G305), .ZN(n678) );
  XNOR2_X1 U763 ( .A(n678), .B(n681), .ZN(n919) );
  XNOR2_X1 U764 ( .A(n679), .B(n919), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n680), .A2(G868), .ZN(n684) );
  NAND2_X1 U766 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U767 ( .A1(n684), .A2(n683), .ZN(G295) );
  NAND2_X1 U768 ( .A1(G2078), .A2(G2084), .ZN(n685) );
  XNOR2_X1 U769 ( .A(n685), .B(KEYINPUT85), .ZN(n686) );
  XNOR2_X1 U770 ( .A(n686), .B(KEYINPUT20), .ZN(n687) );
  NAND2_X1 U771 ( .A1(n687), .A2(G2090), .ZN(n688) );
  XNOR2_X1 U772 ( .A(KEYINPUT21), .B(n688), .ZN(n689) );
  NAND2_X1 U773 ( .A1(n689), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U774 ( .A(KEYINPUT86), .B(n690), .ZN(G158) );
  XNOR2_X1 U775 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U776 ( .A1(G220), .A2(G219), .ZN(n691) );
  XOR2_X1 U777 ( .A(KEYINPUT22), .B(n691), .Z(n692) );
  NOR2_X1 U778 ( .A1(G218), .A2(n692), .ZN(n693) );
  NAND2_X1 U779 ( .A1(G96), .A2(n693), .ZN(n937) );
  NAND2_X1 U780 ( .A1(n937), .A2(G2106), .ZN(n697) );
  NAND2_X1 U781 ( .A1(G120), .A2(G108), .ZN(n694) );
  NOR2_X1 U782 ( .A1(G237), .A2(n694), .ZN(n695) );
  NAND2_X1 U783 ( .A1(G69), .A2(n695), .ZN(n938) );
  NAND2_X1 U784 ( .A1(n938), .A2(G567), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n697), .A2(n696), .ZN(n851) );
  NAND2_X1 U786 ( .A1(G483), .A2(G661), .ZN(n698) );
  NOR2_X1 U787 ( .A1(n851), .A2(n698), .ZN(n699) );
  XOR2_X1 U788 ( .A(KEYINPUT87), .B(n699), .Z(n850) );
  NAND2_X1 U789 ( .A1(n850), .A2(G36), .ZN(G176) );
  NAND2_X1 U790 ( .A1(n890), .A2(G101), .ZN(n700) );
  XOR2_X1 U791 ( .A(KEYINPUT23), .B(n700), .Z(n702) );
  NAND2_X1 U792 ( .A1(n895), .A2(G125), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U794 ( .A(n703), .B(KEYINPUT64), .ZN(n707) );
  NAND2_X1 U795 ( .A1(G137), .A2(n891), .ZN(n705) );
  NAND2_X1 U796 ( .A1(G113), .A2(n894), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U798 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NAND2_X1 U799 ( .A1(G160), .A2(G40), .ZN(n782) );
  NAND2_X1 U800 ( .A1(n734), .A2(G2072), .ZN(n708) );
  XOR2_X1 U801 ( .A(KEYINPUT27), .B(n708), .Z(n711) );
  NAND2_X1 U802 ( .A1(G1956), .A2(n753), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n728) );
  OR2_X1 U804 ( .A1(G299), .A2(n728), .ZN(n723) );
  INV_X1 U805 ( .A(n723), .ZN(n717) );
  NAND2_X1 U806 ( .A1(G1996), .A2(n734), .ZN(n712) );
  XNOR2_X1 U807 ( .A(KEYINPUT26), .B(n712), .ZN(n715) );
  NOR2_X1 U808 ( .A1(n1003), .A2(n713), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n716) );
  OR2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n727) );
  XNOR2_X1 U812 ( .A(n720), .B(KEYINPUT99), .ZN(n726) );
  NOR2_X1 U813 ( .A1(n734), .A2(G1348), .ZN(n722) );
  NOR2_X1 U814 ( .A1(G2067), .A2(n753), .ZN(n721) );
  NOR2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n724) );
  AND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U817 ( .A(KEYINPUT97), .B(KEYINPUT28), .Z(n730) );
  NAND2_X1 U818 ( .A1(n728), .A2(G299), .ZN(n729) );
  XNOR2_X1 U819 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U820 ( .A(KEYINPUT101), .B(KEYINPUT29), .ZN(n732) );
  XNOR2_X1 U821 ( .A(n733), .B(n732), .ZN(n738) );
  XNOR2_X1 U822 ( .A(G2078), .B(KEYINPUT25), .ZN(n1024) );
  NOR2_X1 U823 ( .A1(n753), .A2(n1024), .ZN(n736) );
  INV_X1 U824 ( .A(G1961), .ZN(n986) );
  NOR2_X1 U825 ( .A1(n734), .A2(n986), .ZN(n735) );
  NOR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n745) );
  NAND2_X1 U827 ( .A1(n745), .A2(G171), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n752) );
  NOR2_X1 U829 ( .A1(n823), .A2(G1966), .ZN(n739) );
  XNOR2_X1 U830 ( .A(n739), .B(KEYINPUT96), .ZN(n761) );
  NOR2_X1 U831 ( .A1(n753), .A2(G2084), .ZN(n740) );
  XOR2_X1 U832 ( .A(n740), .B(KEYINPUT95), .Z(n760) );
  INV_X1 U833 ( .A(n760), .ZN(n741) );
  NAND2_X1 U834 ( .A1(G8), .A2(n741), .ZN(n742) );
  NOR2_X1 U835 ( .A1(n761), .A2(n742), .ZN(n743) );
  XOR2_X1 U836 ( .A(KEYINPUT30), .B(n743), .Z(n744) );
  NOR2_X1 U837 ( .A1(G168), .A2(n744), .ZN(n748) );
  NOR2_X1 U838 ( .A1(G171), .A2(n745), .ZN(n746) );
  XNOR2_X1 U839 ( .A(KEYINPUT102), .B(n746), .ZN(n747) );
  NOR2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n750) );
  XNOR2_X1 U841 ( .A(KEYINPUT103), .B(KEYINPUT31), .ZN(n749) );
  XNOR2_X1 U842 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U843 ( .A1(G1971), .A2(n823), .ZN(n755) );
  NOR2_X1 U844 ( .A1(G2090), .A2(n753), .ZN(n754) );
  NOR2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n756), .A2(G303), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n758), .A2(G8), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n759), .B(KEYINPUT32), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G8), .A2(n760), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n517), .A2(n761), .ZN(n762) );
  NAND2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n818) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n766) );
  XNOR2_X1 U854 ( .A(KEYINPUT105), .B(n766), .ZN(n990) );
  INV_X1 U855 ( .A(n990), .ZN(n778) );
  NOR2_X1 U856 ( .A1(G1971), .A2(G303), .ZN(n767) );
  NOR2_X1 U857 ( .A1(n778), .A2(n767), .ZN(n769) );
  INV_X1 U858 ( .A(KEYINPUT33), .ZN(n768) );
  AND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n818), .A2(n770), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G288), .A2(G1976), .ZN(n771) );
  XNOR2_X1 U862 ( .A(n771), .B(KEYINPUT106), .ZN(n989) );
  INV_X1 U863 ( .A(n989), .ZN(n772) );
  NOR2_X1 U864 ( .A1(n772), .A2(n823), .ZN(n773) );
  OR2_X1 U865 ( .A1(KEYINPUT33), .A2(n773), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U867 ( .A1(n778), .A2(KEYINPUT33), .ZN(n779) );
  NOR2_X1 U868 ( .A1(n823), .A2(n779), .ZN(n780) );
  XOR2_X1 U869 ( .A(G1981), .B(G305), .Z(n996) );
  NOR2_X1 U870 ( .A1(G1384), .A2(G164), .ZN(n783) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n840) );
  XNOR2_X1 U872 ( .A(KEYINPUT37), .B(G2067), .ZN(n838) );
  NAND2_X1 U873 ( .A1(G104), .A2(n890), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G140), .A2(n891), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G116), .A2(n894), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G128), .A2(n895), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U880 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U882 ( .A(KEYINPUT36), .B(n792), .ZN(n911) );
  NOR2_X1 U883 ( .A1(n838), .A2(n911), .ZN(n969) );
  NAND2_X1 U884 ( .A1(n840), .A2(n969), .ZN(n836) );
  NAND2_X1 U885 ( .A1(G119), .A2(n895), .ZN(n799) );
  NAND2_X1 U886 ( .A1(G95), .A2(n890), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G107), .A2(n894), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n891), .A2(G131), .ZN(n795) );
  XOR2_X1 U890 ( .A(KEYINPUT92), .B(n795), .Z(n796) );
  NOR2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U892 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U893 ( .A(n800), .B(KEYINPUT93), .Z(n905) );
  AND2_X1 U894 ( .A1(n905), .A2(G1991), .ZN(n810) );
  XOR2_X1 U895 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n802) );
  NAND2_X1 U896 ( .A1(G105), .A2(n890), .ZN(n801) );
  XNOR2_X1 U897 ( .A(n802), .B(n801), .ZN(n806) );
  NAND2_X1 U898 ( .A1(G117), .A2(n894), .ZN(n804) );
  NAND2_X1 U899 ( .A1(G129), .A2(n895), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n891), .A2(G141), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n906) );
  AND2_X1 U904 ( .A1(n906), .A2(G1996), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n974) );
  INV_X1 U906 ( .A(n974), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n811), .A2(n840), .ZN(n830) );
  AND2_X1 U908 ( .A1(n836), .A2(n830), .ZN(n825) );
  AND2_X1 U909 ( .A1(n996), .A2(n825), .ZN(n812) );
  XNOR2_X1 U910 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U911 ( .A1(n993), .A2(n840), .ZN(n815) );
  AND2_X1 U912 ( .A1(n812), .A2(n815), .ZN(n813) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n845) );
  INV_X1 U914 ( .A(n815), .ZN(n829) );
  NOR2_X1 U915 ( .A1(G2090), .A2(G303), .ZN(n816) );
  NAND2_X1 U916 ( .A1(G8), .A2(n816), .ZN(n817) );
  NAND2_X1 U917 ( .A1(n818), .A2(n817), .ZN(n820) );
  AND2_X1 U918 ( .A1(n823), .A2(n825), .ZN(n819) );
  NOR2_X1 U919 ( .A1(G1981), .A2(G305), .ZN(n821) );
  XOR2_X1 U920 ( .A(n821), .B(KEYINPUT24), .Z(n822) );
  NOR2_X1 U921 ( .A1(n823), .A2(n822), .ZN(n824) );
  AND2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U923 ( .A1(n829), .A2(n828), .ZN(n843) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n906), .ZN(n964) );
  INV_X1 U925 ( .A(n830), .ZN(n833) );
  NOR2_X1 U926 ( .A1(G1991), .A2(n905), .ZN(n968) );
  NOR2_X1 U927 ( .A1(G1986), .A2(G290), .ZN(n831) );
  NOR2_X1 U928 ( .A1(n968), .A2(n831), .ZN(n832) );
  NOR2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n834) );
  NOR2_X1 U930 ( .A1(n964), .A2(n834), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n835), .B(KEYINPUT39), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n839) );
  NAND2_X1 U933 ( .A1(n838), .A2(n911), .ZN(n966) );
  NAND2_X1 U934 ( .A1(n839), .A2(n966), .ZN(n841) );
  AND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  NOR2_X1 U936 ( .A1(n843), .A2(n842), .ZN(n844) );
  NAND2_X1 U937 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U938 ( .A(n846), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n847), .ZN(G217) );
  INV_X1 U940 ( .A(n847), .ZN(G223) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n848) );
  NAND2_X1 U942 ( .A1(G661), .A2(n848), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U944 ( .A1(n850), .A2(n849), .ZN(G188) );
  INV_X1 U945 ( .A(n851), .ZN(G319) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n853) );
  XNOR2_X1 U947 ( .A(G2090), .B(G2678), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U949 ( .A(n854), .B(KEYINPUT108), .Z(n856) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2100), .Z(n858) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U955 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n862) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1966), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U959 ( .A(n863), .B(G2474), .Z(n865) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1981), .Z(n867) );
  XOR2_X1 U963 ( .A(G1956), .B(n986), .Z(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G100), .A2(n890), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n870), .B(KEYINPUT110), .ZN(n873) );
  NAND2_X1 U968 ( .A1(G112), .A2(n894), .ZN(n871) );
  XOR2_X1 U969 ( .A(KEYINPUT109), .B(n871), .Z(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U971 ( .A1(G124), .A2(n895), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n874), .B(KEYINPUT44), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n891), .A2(G136), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G118), .A2(n894), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G130), .A2(n895), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n886) );
  NAND2_X1 U979 ( .A1(G106), .A2(n890), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G142), .A2(n891), .ZN(n881) );
  NAND2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(KEYINPUT111), .B(n883), .ZN(n884) );
  XNOR2_X1 U983 ( .A(KEYINPUT45), .B(n884), .ZN(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n910) );
  XOR2_X1 U985 ( .A(KEYINPUT114), .B(KEYINPUT116), .Z(n888) );
  XNOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(n889), .B(KEYINPUT46), .Z(n903) );
  NAND2_X1 U989 ( .A1(G103), .A2(n890), .ZN(n893) );
  NAND2_X1 U990 ( .A1(G139), .A2(n891), .ZN(n892) );
  NAND2_X1 U991 ( .A1(n893), .A2(n892), .ZN(n900) );
  NAND2_X1 U992 ( .A1(G115), .A2(n894), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G127), .A2(n895), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(KEYINPUT47), .B(n898), .Z(n899) );
  NOR2_X1 U996 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(n901), .Z(n976) );
  XNOR2_X1 U998 ( .A(n976), .B(KEYINPUT115), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(n908) );
  XOR2_X1 U1001 ( .A(G164), .B(n906), .Z(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1003 ( .A(n910), .B(n909), .ZN(n913) );
  XNOR2_X1 U1004 ( .A(n911), .B(G162), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(n913), .B(n912), .ZN(n915) );
  XNOR2_X1 U1006 ( .A(n970), .B(G160), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n916), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(G286), .B(KEYINPUT117), .ZN(n918) );
  XOR2_X1 U1010 ( .A(n1000), .B(G171), .Z(n917) );
  XNOR2_X1 U1011 ( .A(n918), .B(n917), .ZN(n921) );
  XOR2_X1 U1012 ( .A(n1003), .B(n919), .Z(n920) );
  XNOR2_X1 U1013 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n922), .ZN(G397) );
  XOR2_X1 U1015 ( .A(G2451), .B(G2430), .Z(n924) );
  XNOR2_X1 U1016 ( .A(G2438), .B(G2443), .ZN(n923) );
  XNOR2_X1 U1017 ( .A(n924), .B(n923), .ZN(n930) );
  XOR2_X1 U1018 ( .A(G2435), .B(G2454), .Z(n926) );
  XNOR2_X1 U1019 ( .A(G1348), .B(G1341), .ZN(n925) );
  XNOR2_X1 U1020 ( .A(n926), .B(n925), .ZN(n928) );
  XOR2_X1 U1021 ( .A(G2446), .B(G2427), .Z(n927) );
  XNOR2_X1 U1022 ( .A(n928), .B(n927), .ZN(n929) );
  XOR2_X1 U1023 ( .A(n930), .B(n929), .Z(n931) );
  NAND2_X1 U1024 ( .A1(G14), .A2(n931), .ZN(n939) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n939), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(G227), .A2(G229), .ZN(n932) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(n932), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n934), .A2(n933), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(G395), .A2(G397), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n936), .A2(n935), .ZN(G225) );
  XOR2_X1 U1031 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  XNOR2_X1 U1032 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U1034 ( .A(G120), .ZN(G236) );
  INV_X1 U1035 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(G325) );
  INV_X1 U1037 ( .A(G325), .ZN(G261) );
  INV_X1 U1038 ( .A(G69), .ZN(G235) );
  INV_X1 U1039 ( .A(n939), .ZN(G401) );
  XOR2_X1 U1040 ( .A(G5), .B(G1961), .Z(n957) );
  XOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .Z(n940) );
  XNOR2_X1 U1042 ( .A(G4), .B(n940), .ZN(n942) );
  XNOR2_X1 U1043 ( .A(G20), .B(G1956), .ZN(n941) );
  NOR2_X1 U1044 ( .A1(n942), .A2(n941), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1046 ( .A(G1981), .B(G6), .ZN(n943) );
  NOR2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1049 ( .A(n947), .B(KEYINPUT60), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G22), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(G23), .B(G1976), .ZN(n948) );
  NOR2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(G1986), .B(KEYINPUT127), .ZN(n950) );
  XNOR2_X1 U1054 ( .A(n950), .B(G24), .ZN(n951) );
  NAND2_X1 U1055 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1056 ( .A(KEYINPUT58), .B(n953), .ZN(n954) );
  NOR2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n959) );
  XNOR2_X1 U1059 ( .A(G21), .B(G1966), .ZN(n958) );
  NOR2_X1 U1060 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1061 ( .A(KEYINPUT61), .B(n960), .ZN(n961) );
  INV_X1 U1062 ( .A(G16), .ZN(n1011) );
  NAND2_X1 U1063 ( .A1(n961), .A2(n1011), .ZN(n962) );
  NAND2_X1 U1064 ( .A1(n962), .A2(G11), .ZN(n1017) );
  XOR2_X1 U1065 ( .A(G2090), .B(G162), .Z(n963) );
  NOR2_X1 U1066 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1067 ( .A(KEYINPUT51), .B(n965), .Z(n967) );
  NAND2_X1 U1068 ( .A1(n967), .A2(n966), .ZN(n973) );
  NOR2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n971) );
  NAND2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G160), .B(G2084), .ZN(n975) );
  NAND2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n981) );
  XOR2_X1 U1074 ( .A(G2072), .B(n976), .Z(n978) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1077 ( .A(KEYINPUT50), .B(n979), .Z(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(n984), .B(KEYINPUT52), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n985), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1082 ( .A(G171), .B(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(G299), .B(G1956), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1086 ( .A(KEYINPUT125), .B(n991), .Z(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n1009) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G168), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(n998), .B(KEYINPUT57), .ZN(n999) );
  XNOR2_X1 U1092 ( .A(KEYINPUT124), .B(n999), .ZN(n1007) );
  XOR2_X1 U1093 ( .A(G1971), .B(G303), .Z(n1002) );
  XNOR2_X1 U1094 ( .A(G1348), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(G1341), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1010), .Z(n1013) );
  XOR2_X1 U1101 ( .A(n1011), .B(KEYINPUT56), .Z(n1012) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1041) );
  XNOR2_X1 U1105 ( .A(G1991), .B(G25), .ZN(n1022) );
  XNOR2_X1 U1106 ( .A(G2067), .B(G26), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(G2072), .B(G33), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(KEYINPUT121), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(G28), .A2(n1023), .ZN(n1029) );
  XOR2_X1 U1112 ( .A(n1024), .B(G27), .Z(n1026) );
  XNOR2_X1 U1113 ( .A(G1996), .B(G32), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1115 ( .A(KEYINPUT122), .B(n1027), .Z(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1117 ( .A(KEYINPUT53), .B(n1030), .Z(n1034) );
  XNOR2_X1 U1118 ( .A(KEYINPUT54), .B(G34), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(n1031), .B(KEYINPUT123), .ZN(n1032) );
  XNOR2_X1 U1120 ( .A(G2084), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1037) );
  XNOR2_X1 U1122 ( .A(KEYINPUT120), .B(G2090), .ZN(n1035) );
  XNOR2_X1 U1123 ( .A(G35), .B(n1035), .ZN(n1036) );
  NOR2_X1 U1124 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1125 ( .A1(G29), .A2(n1038), .ZN(n1039) );
  XNOR2_X1 U1126 ( .A(n1039), .B(KEYINPUT55), .ZN(n1040) );
  NAND2_X1 U1127 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1128 ( .A(KEYINPUT62), .B(n1042), .ZN(G150) );
  INV_X1 U1129 ( .A(G150), .ZN(G311) );
endmodule

