//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n210), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT64), .Z(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n216), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT65), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G107), .B(G116), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  NAND3_X1  g0042(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(new_n211), .ZN(new_n244));
  INV_X1    g0044(.A(KEYINPUT69), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(KEYINPUT8), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT8), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT70), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n212), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI22_X1  g0063(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n265));
  OAI21_X1  g0065(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(new_n264), .B2(KEYINPUT71), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n249), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G20), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT72), .ZN(new_n271));
  INV_X1    g0071(.A(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n248), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G50), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n268), .B(new_n277), .C1(G50), .C2(new_n274), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  OAI21_X1  g0080(.A(KEYINPUT66), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT66), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G222), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G223), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n290), .B1(new_n291), .B2(new_n288), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT67), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n295), .A2(new_n298), .A3(G1), .A4(G13), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n294), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n303));
  INV_X1    g0103(.A(G274), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n296), .A2(new_n303), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(G226), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n302), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n302), .A2(KEYINPUT68), .A3(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n278), .B1(new_n314), .B2(G179), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(G169), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n278), .B(KEYINPUT9), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(G200), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(G190), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT10), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT10), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n318), .A2(new_n319), .A3(new_n323), .A4(new_n320), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n317), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  NOR2_X1   g0126(.A1(G226), .A2(G1698), .ZN(new_n327));
  INV_X1    g0127(.A(G232), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(G1698), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n281), .A2(new_n329), .A3(new_n287), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT74), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(G33), .B2(G97), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(KEYINPUT74), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n301), .ZN(new_n337));
  INV_X1    g0137(.A(new_n305), .ZN(new_n338));
  INV_X1    g0138(.A(G238), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n306), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n326), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n300), .B1(new_n330), .B2(new_n335), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n343), .A2(KEYINPUT13), .A3(new_n340), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G190), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n276), .A2(G68), .ZN(new_n347));
  INV_X1    g0147(.A(new_n274), .ZN(new_n348));
  INV_X1    g0148(.A(G68), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT12), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n262), .A2(G50), .B1(G20), .B2(new_n349), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n291), .B2(new_n260), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n249), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT11), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n249), .A2(new_n353), .A3(KEYINPUT11), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n351), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n346), .A2(new_n347), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n345), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n337), .A2(new_n326), .A3(new_n341), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT13), .B1(new_n343), .B2(new_n340), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n363), .A2(G179), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G169), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n363), .B2(new_n364), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI211_X1 g0169(.A(KEYINPUT14), .B(new_n366), .C1(new_n363), .C2(new_n364), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT75), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(G169), .B1(new_n342), .B2(new_n344), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT14), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n367), .A2(new_n368), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .A4(new_n365), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n358), .A2(new_n347), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n362), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n250), .A2(new_n349), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n380), .B2(new_n201), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n262), .A2(G159), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n279), .A2(new_n280), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT76), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n384), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n212), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n284), .A2(new_n286), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(G20), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n383), .B1(new_n392), .B2(G68), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n248), .B1(new_n393), .B2(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(new_n383), .ZN(new_n395));
  INV_X1    g0195(.A(new_n385), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n281), .A2(new_n287), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n212), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n396), .B1(new_n398), .B2(new_n389), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n395), .B1(new_n399), .B2(new_n349), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n293), .A2(new_n289), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(G226), .B2(new_n289), .C1(new_n279), .C2(new_n280), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n300), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n338), .B1(new_n306), .B2(new_n328), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT79), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n406), .A2(new_n404), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n301), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n408), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT79), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n414), .A3(new_n360), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT78), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n338), .B(KEYINPUT78), .C1(new_n328), .C2(new_n306), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(KEYINPUT80), .A2(G190), .ZN(new_n420));
  NOR2_X1   g0220(.A1(KEYINPUT80), .A2(G190), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT81), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n422), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n407), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n426), .A2(new_n427), .A3(new_n417), .A4(new_n418), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n415), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n259), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n275), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n259), .A2(new_n274), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT77), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT77), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n432), .C1(new_n276), .C2(new_n259), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n403), .A2(new_n429), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n403), .A2(new_n437), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT18), .ZN(new_n442));
  INV_X1    g0242(.A(G179), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n411), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n419), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n409), .A2(new_n414), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(new_n366), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n441), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n394), .A2(new_n402), .B1(new_n434), .B2(new_n436), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n446), .A2(G169), .B1(new_n419), .B2(new_n444), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT18), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(KEYINPUT17), .A3(new_n429), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n440), .A2(new_n449), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n288), .A2(G232), .A3(new_n289), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  OAI221_X1 g0257(.A(new_n456), .B1(new_n457), .B2(new_n288), .C1(new_n292), .C2(new_n339), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n301), .ZN(new_n459));
  INV_X1    g0259(.A(G244), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n338), .B1(new_n306), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n443), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n276), .A2(G77), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n348), .A2(new_n291), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT15), .B(G87), .ZN(new_n466));
  OAI22_X1  g0266(.A1(new_n466), .A2(new_n260), .B1(new_n212), .B2(new_n291), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n256), .A2(new_n263), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n249), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n464), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n461), .B1(new_n458), .B2(new_n301), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n473), .B2(new_n366), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n470), .B1(new_n473), .B2(G200), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(G190), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n463), .A2(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT73), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n325), .A2(new_n379), .A3(new_n455), .A4(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n482));
  INV_X1    g0282(.A(G45), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G1), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G270), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n485), .A2(new_n296), .A3(G274), .A4(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G257), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n289), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n289), .A2(G264), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n390), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G303), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n288), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n300), .B1(new_n495), .B2(KEYINPUT85), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT85), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n497), .B(new_n493), .C1(new_n288), .C2(new_n494), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n489), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n269), .A2(G33), .ZN(new_n500));
  AND3_X1   g0300(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT69), .B1(new_n243), .B2(new_n211), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n274), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G116), .ZN(new_n504));
  OR2_X1    g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  INV_X1    g0306(.A(G97), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n212), .C1(G33), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(G20), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n244), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT20), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n273), .A2(G20), .A3(new_n504), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n505), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G169), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n481), .B1(new_n499), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n499), .A2(G179), .A3(new_n514), .ZN(new_n517));
  INV_X1    g0317(.A(new_n493), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n494), .B1(new_n281), .B2(new_n287), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT85), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(new_n498), .A3(new_n301), .ZN(new_n521));
  INV_X1    g0321(.A(new_n489), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(new_n514), .A3(KEYINPUT21), .A4(G169), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n516), .A2(new_n517), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n499), .A2(new_n360), .ZN(new_n526));
  INV_X1    g0326(.A(new_n514), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n523), .B2(new_n422), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g0329(.A1(KEYINPUT5), .A2(G41), .ZN(new_n530));
  NOR2_X1   g0330(.A1(KEYINPUT5), .A2(G41), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n484), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(G264), .A3(new_n296), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G250), .A2(G1698), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n490), .B2(G1698), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(new_n390), .B1(G33), .B2(G294), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n533), .B(new_n488), .C1(new_n536), .C2(new_n300), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(G179), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n366), .B2(new_n537), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n212), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT22), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  OR3_X1    g0342(.A1(new_n542), .A2(KEYINPUT22), .A3(G20), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n397), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT23), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n457), .A3(G20), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(KEYINPUT87), .A2(KEYINPUT24), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n544), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n555), .B1(new_n544), .B2(new_n553), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n556), .A2(new_n557), .A3(new_n248), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n348), .A2(KEYINPUT25), .A3(new_n457), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n274), .B2(G107), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n503), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n248), .A2(KEYINPUT82), .A3(new_n274), .A4(new_n500), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n566), .B2(new_n457), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n539), .B1(new_n558), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n525), .A2(new_n529), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n571), .A2(new_n460), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n281), .A2(new_n287), .A3(new_n289), .A4(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n506), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n460), .A2(G1698), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n279), .B2(new_n280), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n574), .B1(new_n576), .B2(new_n571), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n281), .A2(new_n287), .A3(G250), .A4(G1698), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n301), .ZN(new_n580));
  INV_X1    g0380(.A(G190), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n532), .A2(G257), .A3(new_n296), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n488), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n580), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n583), .B1(new_n579), .B2(new_n301), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(G200), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n274), .A2(G97), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n457), .A2(KEYINPUT6), .A3(G97), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT6), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n592), .A2(new_n212), .B1(new_n291), .B2(new_n263), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n399), .B2(new_n457), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n588), .B1(new_n595), .B2(new_n249), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n564), .A2(new_n565), .A3(G97), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n587), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n535), .A2(new_n390), .ZN(new_n599));
  NAND2_X1  g0399(.A1(G33), .A2(G294), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n301), .B1(new_n486), .B2(G264), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(KEYINPUT88), .A3(new_n581), .A4(new_n488), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n537), .B2(new_n360), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n537), .A2(G190), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n603), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n544), .A2(new_n553), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n248), .B1(new_n608), .B2(new_n554), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n608), .B2(new_n554), .ZN(new_n610));
  INV_X1    g0410(.A(new_n567), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n588), .ZN(new_n613));
  AOI21_X1  g0413(.A(G20), .B1(new_n281), .B2(new_n287), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n385), .B1(new_n614), .B2(KEYINPUT7), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n593), .B1(new_n615), .B2(G107), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n597), .B(new_n613), .C1(new_n616), .C2(new_n248), .ZN(new_n617));
  AOI211_X1 g0417(.A(G179), .B(new_n583), .C1(new_n579), .C2(new_n301), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n580), .A2(new_n584), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n366), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n598), .A2(new_n612), .A3(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n466), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n564), .A2(new_n565), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT19), .B1(new_n332), .B2(new_n334), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n212), .B1(new_n542), .B2(new_n204), .ZN(new_n627));
  AOI21_X1  g0427(.A(G20), .B1(new_n284), .B2(new_n286), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G68), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT19), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n249), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n624), .A2(new_n274), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n625), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT84), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n333), .A2(KEYINPUT74), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n331), .A2(G33), .A3(G97), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n631), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n642), .A2(G20), .B1(G87), .B2(new_n205), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n628), .A2(G68), .B1(new_n631), .B2(new_n630), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n635), .B1(new_n645), .B2(new_n249), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(KEYINPUT84), .A3(new_n625), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n283), .A2(new_n504), .ZN(new_n648));
  NOR2_X1   g0448(.A1(G238), .A2(G1698), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n460), .B2(G1698), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(new_n390), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(new_n300), .ZN(new_n652));
  INV_X1    g0452(.A(G250), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n484), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n296), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n654), .A2(KEYINPUT83), .A3(new_n296), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n484), .A2(G274), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n652), .A2(new_n659), .A3(G179), .A4(new_n660), .ZN(new_n661));
  NOR4_X1   g0461(.A1(new_n482), .A2(new_n656), .A3(new_n484), .A4(new_n653), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT83), .B1(new_n654), .B2(new_n296), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n660), .B1(new_n651), .B2(new_n300), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n661), .B1(new_n666), .B2(new_n366), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n639), .A2(new_n647), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(G200), .B1(new_n664), .B2(new_n665), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n652), .A2(new_n659), .A3(G190), .A4(new_n660), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n564), .A2(new_n565), .A3(G87), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n634), .A3(new_n636), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n668), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n623), .A2(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n480), .A2(new_n570), .A3(new_n677), .ZN(G372));
  NAND3_X1  g0478(.A1(new_n652), .A2(new_n659), .A3(new_n660), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G169), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n680), .A2(new_n661), .B1(new_n637), .B2(new_n638), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n681), .A2(new_n647), .B1(new_n674), .B2(new_n671), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT92), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n617), .A2(new_n619), .A3(new_n621), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT26), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(KEYINPUT26), .A3(new_n675), .A4(new_n668), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(KEYINPUT92), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT89), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n646), .A2(new_n688), .A3(new_n672), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n688), .B1(new_n646), .B2(new_n672), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n671), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n667), .A2(new_n637), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND4_X1   g0493(.A1(KEYINPUT91), .A2(new_n617), .A3(new_n619), .A4(new_n621), .ZN(new_n694));
  AOI21_X1  g0494(.A(G169), .B1(new_n580), .B2(new_n584), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n618), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT91), .B1(new_n696), .B2(new_n617), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n693), .A2(new_n694), .A3(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n685), .B(new_n687), .C1(new_n698), .C2(KEYINPUT26), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n623), .A2(new_n693), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n568), .A2(new_n516), .A3(new_n517), .A4(new_n524), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT90), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND4_X1   g0502(.A1(new_n568), .A2(new_n516), .A3(new_n517), .A4(new_n524), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT90), .ZN(new_n704));
  NOR4_X1   g0504(.A1(new_n703), .A2(new_n623), .A3(new_n693), .A4(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n699), .B(new_n692), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n480), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n377), .A2(new_n378), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n463), .B(new_n470), .C1(G169), .C2(new_n472), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n362), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n440), .A3(new_n453), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n449), .A2(new_n452), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n322), .A2(new_n324), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n317), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n707), .A2(new_n715), .ZN(G369));
  INV_X1    g0516(.A(new_n273), .ZN(new_n717));
  OR3_X1    g0517(.A1(new_n717), .A2(KEYINPUT27), .A3(G20), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT27), .B1(new_n717), .B2(G20), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G213), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G343), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n527), .A2(new_n723), .ZN(new_n724));
  OR3_X1    g0524(.A1(new_n525), .A2(new_n529), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n525), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n569), .A2(new_n722), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n722), .B1(new_n558), .B2(new_n567), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n612), .A2(new_n568), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n727), .A2(G330), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n569), .A2(new_n723), .ZN(new_n733));
  INV_X1    g0533(.A(new_n525), .ZN(new_n734));
  OR3_X1    g0534(.A1(new_n734), .A2(new_n722), .A3(new_n730), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(G399));
  INV_X1    g0536(.A(new_n208), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G41), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n739), .A2(G1), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n214), .B2(new_n739), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  OR2_X1    g0543(.A1(KEYINPUT93), .A2(KEYINPUT30), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n586), .A2(new_n666), .A3(new_n602), .A4(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n521), .A2(G179), .A3(new_n522), .ZN(new_n746));
  NAND2_X1  g0546(.A1(KEYINPUT93), .A2(KEYINPUT30), .ZN(new_n747));
  OR3_X1    g0547(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n747), .B1(new_n745), .B2(new_n746), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n537), .A2(new_n443), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n523), .A2(new_n679), .A3(new_n620), .A4(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n752), .A2(KEYINPUT31), .A3(new_n722), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT31), .B1(new_n752), .B2(new_n722), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n570), .A2(new_n677), .A3(new_n723), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G330), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n680), .A2(new_n661), .B1(new_n646), .B2(new_n625), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n673), .A2(KEYINPUT89), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n646), .A2(new_n688), .A3(new_n672), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n762), .B1(new_n765), .B2(new_n671), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n766), .A2(new_n622), .A3(new_n598), .A4(new_n612), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n704), .B1(new_n767), .B2(new_n703), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n700), .A2(KEYINPUT90), .A3(new_n701), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n762), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n722), .B1(new_n770), .B2(new_n699), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n682), .A2(new_n684), .ZN(new_n775));
  MUX2_X1   g0575(.A(new_n775), .B(new_n698), .S(KEYINPUT26), .Z(new_n776));
  AOI21_X1  g0576(.A(new_n762), .B1(new_n700), .B2(new_n701), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n722), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT29), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n761), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n743), .B1(new_n780), .B2(G1), .ZN(G364));
  NOR2_X1   g0581(.A1(new_n272), .A2(G20), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n269), .B1(new_n782), .B2(G45), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n738), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(new_n727), .B2(G330), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G330), .B2(new_n727), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT95), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT95), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n211), .B1(G20), .B2(new_n366), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT97), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n737), .A2(new_n390), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G45), .B2(new_n214), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n241), .B2(G45), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n288), .A2(new_n208), .ZN(new_n799));
  INV_X1    g0599(.A(G355), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n799), .A2(new_n800), .B1(G116), .B2(new_n208), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n795), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n785), .B(KEYINPUT96), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n212), .A2(new_n443), .A3(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n425), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n581), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n807), .A2(G322), .B1(G311), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G294), .ZN(new_n811));
  NOR3_X1   g0611(.A1(new_n581), .A2(G179), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(new_n212), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n810), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n422), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT98), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n816), .A2(new_n817), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n814), .B1(G326), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n815), .A2(G190), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT102), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n360), .A2(G179), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(G20), .A3(G190), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n212), .A2(G190), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n830), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n832), .A2(G303), .B1(new_n835), .B2(G283), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n829), .A2(new_n397), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n833), .A2(new_n443), .A3(new_n360), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n838), .A2(KEYINPUT101), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(KEYINPUT101), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n837), .B1(G329), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n823), .A2(new_n843), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n813), .A2(new_n507), .B1(new_n825), .B2(new_n349), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT100), .Z(new_n846));
  XOR2_X1   g0646(.A(KEYINPUT99), .B(G159), .Z(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n838), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT32), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n806), .A2(new_n250), .B1(new_n291), .B2(new_n808), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n834), .A2(new_n457), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n397), .B(new_n854), .C1(G87), .C2(new_n832), .ZN(new_n855));
  INV_X1    g0655(.A(G50), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n853), .B(new_n855), .C1(new_n856), .C2(new_n821), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n844), .B1(new_n846), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n804), .B1(new_n858), .B2(new_n793), .ZN(new_n859));
  INV_X1    g0659(.A(new_n792), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n727), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n788), .A2(new_n789), .A3(new_n861), .ZN(G396));
  NAND2_X1  g0662(.A1(new_n470), .A2(new_n722), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT104), .B1(new_n709), .B2(new_n723), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT104), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n474), .A2(new_n865), .A3(new_n463), .A4(new_n722), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n477), .A2(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n771), .B(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n761), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n785), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n384), .B1(new_n832), .B2(G50), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n873), .B1(new_n250), .B2(new_n813), .C1(new_n349), .C2(new_n834), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n807), .A2(G143), .B1(new_n809), .B2(new_n848), .ZN(new_n875));
  INV_X1    g0675(.A(G137), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n875), .B1(new_n261), .B2(new_n825), .C1(new_n821), .C2(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(new_n877), .B(KEYINPUT34), .Z(new_n878));
  AOI211_X1 g0678(.A(new_n874), .B(new_n878), .C1(G132), .C2(new_n842), .ZN(new_n879));
  INV_X1    g0679(.A(G283), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n808), .A2(new_n504), .B1(new_n825), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n822), .B2(G303), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT103), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n842), .A2(G311), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n397), .B1(new_n542), .B2(new_n834), .C1(new_n457), .C2(new_n831), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n806), .A2(new_n811), .B1(new_n507), .B2(new_n813), .ZN(new_n886));
  NOR4_X1   g0686(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n793), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n803), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n793), .A2(new_n790), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n291), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n888), .B(new_n891), .C1(new_n868), .C2(new_n791), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n872), .A2(new_n892), .ZN(G384));
  INV_X1    g0693(.A(new_n592), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT35), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(KEYINPUT35), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n895), .A2(G116), .A3(new_n213), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT36), .Z(new_n898));
  OR3_X1    g0698(.A1(new_n214), .A2(new_n291), .A3(new_n380), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n856), .A2(G68), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n269), .B(G13), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n903));
  AOI21_X1  g0703(.A(new_n867), .B1(new_n755), .B2(new_n757), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT106), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n378), .A2(new_n722), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n371), .B2(new_n376), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(KEYINPUT105), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n905), .B(new_n907), .C1(new_n379), .C2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n362), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n708), .A2(new_n910), .A3(new_n908), .ZN(new_n911));
  INV_X1    g0711(.A(new_n907), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT106), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n904), .B1(new_n909), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n392), .A2(G68), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n915), .A2(KEYINPUT16), .A3(new_n395), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n249), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n393), .A2(KEYINPUT16), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n437), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n720), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n448), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n922), .A3(new_n438), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT37), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n441), .A2(new_n448), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n441), .A2(new_n920), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT37), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .A4(new_n438), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n921), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n454), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT38), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT38), .B1(new_n929), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n903), .B1(new_n914), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n911), .A2(new_n912), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n905), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n911), .A2(KEYINPUT106), .A3(new_n912), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT38), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n925), .A2(new_n926), .A3(new_n438), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n942));
  INV_X1    g0742(.A(new_n926), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n942), .A2(new_n928), .B1(new_n454), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n940), .B1(new_n944), .B2(KEYINPUT38), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n939), .A2(KEYINPUT40), .A3(new_n945), .A4(new_n904), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n935), .A2(new_n946), .A3(G330), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n480), .A2(new_n761), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT109), .Z(new_n950));
  NOR2_X1   g0750(.A1(new_n479), .A2(new_n759), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n935), .A3(new_n946), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n706), .A2(new_n723), .A3(new_n868), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n709), .A2(new_n722), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n954), .A2(new_n956), .B1(new_n937), .B2(new_n938), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n932), .B2(new_n933), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n377), .A2(new_n378), .A3(new_n723), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n944), .A2(KEYINPUT38), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT107), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT39), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n940), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT107), .B1(new_n945), .B2(KEYINPUT39), .ZN(new_n965));
  INV_X1    g0765(.A(new_n933), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n966), .B2(new_n940), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n960), .B(new_n964), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n712), .A2(new_n920), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n958), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n480), .A2(new_n779), .A3(new_n774), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n715), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n970), .B(new_n972), .Z(new_n973));
  NAND2_X1  g0773(.A1(new_n953), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n269), .B2(new_n782), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n953), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n902), .B1(new_n975), .B2(new_n976), .ZN(G367));
  INV_X1    g0777(.A(new_n780), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n735), .A2(new_n733), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n617), .A2(new_n722), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n598), .A2(new_n622), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n684), .A2(new_n722), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT110), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n986), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n985), .C2(KEYINPUT44), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n979), .A2(new_n983), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n989), .B(new_n993), .C1(KEYINPUT111), .C2(new_n732), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n732), .A2(KEYINPUT111), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n994), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n727), .A2(G330), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n734), .A2(new_n722), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n735), .B1(new_n731), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n998), .B(new_n1000), .Z(new_n1001));
  AOI21_X1  g0801(.A(new_n978), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n738), .B(KEYINPUT41), .Z(new_n1003));
  OAI21_X1  g0803(.A(new_n783), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n763), .A2(new_n764), .A3(new_n722), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n766), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n692), .B2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n735), .A2(new_n983), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT42), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n622), .B1(new_n981), .B2(new_n568), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(new_n723), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1008), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1007), .A2(KEYINPUT43), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n732), .A2(new_n983), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1004), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n813), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n807), .A2(G150), .B1(new_n1019), .B2(G68), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n825), .B2(new_n847), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n834), .A2(new_n291), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G137), .B2(new_n849), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n250), .B2(new_n831), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n288), .B1(new_n856), .B2(new_n808), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(G143), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n821), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n822), .A2(G311), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT112), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n831), .B2(new_n504), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1031), .A2(KEYINPUT46), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(KEYINPUT113), .B(G317), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n384), .B1(new_n834), .B2(new_n507), .C1(new_n838), .C2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(KEYINPUT46), .B2(new_n1031), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n806), .A2(new_n494), .B1(new_n811), .B2(new_n825), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n808), .A2(new_n880), .B1(new_n813), .B2(new_n457), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1029), .A2(new_n1032), .A3(new_n1035), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1028), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT47), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n793), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n234), .A2(new_n796), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n793), .B(new_n792), .C1(new_n737), .C2(new_n624), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n889), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1042), .B(new_n1045), .C1(new_n860), .C2(new_n1007), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1018), .A2(new_n1046), .ZN(G387));
  NAND2_X1  g0847(.A1(new_n822), .A2(G159), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n813), .A2(new_n466), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n808), .A2(new_n349), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G50), .C2(new_n807), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n831), .A2(new_n291), .B1(new_n838), .B2(new_n261), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n384), .B(new_n1052), .C1(G97), .C2(new_n835), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n430), .A2(new_n824), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1048), .A2(new_n1051), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n390), .B1(new_n849), .B2(G326), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n813), .A2(new_n880), .B1(new_n831), .B2(new_n811), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n806), .A2(new_n1033), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G311), .B2(new_n824), .ZN(new_n1059));
  INV_X1    g0859(.A(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(new_n494), .B2(new_n808), .C1(new_n821), .C2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT115), .Z(new_n1062));
  AOI21_X1  g0862(.A(new_n1057), .B1(new_n1062), .B2(KEYINPUT48), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1056), .B1(new_n504), .B2(new_n834), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1055), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n793), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n231), .A2(new_n483), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT114), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n254), .A2(new_n856), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT50), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n740), .B(new_n483), .C1(new_n349), .C2(new_n291), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n796), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(G107), .B2(new_n208), .C1(new_n740), .C2(new_n799), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n889), .B1(new_n1078), .B2(new_n795), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT116), .B1(new_n1069), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n731), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(new_n792), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1069), .A2(KEYINPUT116), .A3(new_n1079), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n1082), .A2(new_n1083), .B1(new_n784), .B2(new_n1001), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n780), .A2(new_n1001), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n738), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n780), .A2(new_n1001), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(G393));
  NAND2_X1  g0888(.A1(new_n238), .A2(new_n796), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(new_n794), .C1(new_n507), .C2(new_n208), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n889), .B1(new_n1090), .B2(KEYINPUT117), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(KEYINPUT117), .B2(new_n1090), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n822), .A2(G317), .B1(G311), .B2(new_n807), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT52), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n397), .B1(new_n825), .B2(new_n494), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n808), .A2(new_n811), .B1(new_n813), .B2(new_n504), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n854), .B1(G283), .B2(new_n832), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n1060), .C2(new_n838), .ZN(new_n1099));
  INV_X1    g0899(.A(G159), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n821), .A2(new_n261), .B1(new_n1100), .B2(new_n806), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT51), .Z(new_n1102));
  OAI22_X1  g0902(.A1(new_n813), .A2(new_n291), .B1(new_n825), .B2(new_n856), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(new_n254), .B2(new_n809), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n384), .B1(new_n835), .B2(G87), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G68), .A2(new_n832), .B1(new_n849), .B2(G143), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1094), .A2(new_n1099), .B1(new_n1102), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1092), .B1(new_n1108), .B2(new_n793), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n983), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1109), .B1(new_n1110), .B2(new_n860), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n994), .B(new_n995), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n783), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1085), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n739), .B1(new_n997), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1085), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(KEYINPUT121), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT119), .B1(new_n957), .B2(new_n960), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT119), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n955), .B1(new_n771), .B2(new_n868), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n909), .A2(new_n913), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1122), .B(new_n959), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1120), .A2(new_n1121), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n945), .A2(new_n959), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n955), .B1(new_n778), .B2(new_n868), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(KEYINPUT118), .C1(new_n1124), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT118), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n776), .A2(new_n777), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n723), .A3(new_n868), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1133), .A2(new_n956), .B1(new_n937), .B2(new_n938), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1131), .B1(new_n1134), .B2(new_n1127), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1126), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n904), .A2(G330), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1124), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1139), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1126), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1140), .A2(new_n784), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1121), .A2(new_n790), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n831), .A2(new_n261), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT53), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n397), .B1(G50), .B2(new_n835), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1147), .B(new_n1148), .C1(new_n1149), .C2(new_n841), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n807), .A2(G132), .B1(G137), .B2(new_n824), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT54), .B(G143), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1151), .B1(new_n1100), .B2(new_n813), .C1(new_n808), .C2(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1150), .B(new_n1153), .C1(G128), .C2(new_n822), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n821), .A2(new_n880), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n832), .A2(G87), .B1(new_n835), .B2(G68), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1156), .B(new_n397), .C1(new_n841), .C2(new_n811), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n808), .A2(new_n507), .B1(new_n813), .B2(new_n291), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n806), .A2(new_n504), .B1(new_n457), .B2(new_n825), .ZN(new_n1159));
  NOR4_X1   g0959(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n793), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n890), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1161), .B(new_n803), .C1(new_n430), .C2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1145), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT120), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1145), .A2(KEYINPUT120), .A3(new_n1163), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1119), .B1(new_n1144), .B2(new_n1168), .ZN(new_n1169));
  OR2_X1    g0969(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(KEYINPUT121), .A3(new_n1143), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n971), .A2(new_n948), .A3(new_n715), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1124), .A2(new_n1138), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1141), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1123), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1141), .A2(new_n1174), .A3(new_n1129), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n739), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1140), .A2(new_n1142), .A3(new_n1179), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1169), .A2(new_n1171), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(G378));
  INV_X1    g0984(.A(KEYINPUT124), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n947), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n935), .A2(new_n946), .A3(KEYINPUT124), .A4(G330), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n278), .A2(new_n920), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n322), .A2(new_n324), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n317), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n325), .A2(new_n1188), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1193), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n325), .A2(new_n1188), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1189), .B(new_n317), .C1(new_n322), .C2(new_n324), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1186), .A2(new_n1187), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1194), .A2(new_n1198), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1201), .A2(new_n947), .A3(new_n1185), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1200), .A2(new_n970), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n970), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n784), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n785), .B1(new_n1162), .B2(G50), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT123), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G41), .B(new_n390), .C1(new_n832), .C2(G77), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n250), .B2(new_n834), .C1(new_n880), .C2(new_n841), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT122), .Z(new_n1211));
  AOI22_X1  g1011(.A1(new_n1019), .A2(G68), .B1(new_n824), .B2(G97), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n457), .B2(new_n806), .C1(new_n466), .C2(new_n808), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(G116), .B2(new_n822), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n279), .A2(G41), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1215), .A2(KEYINPUT58), .B1(new_n856), .B2(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n809), .A2(G137), .B1(G132), .B2(new_n824), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G150), .B2(new_n1019), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n831), .A2(new_n1152), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n807), .B2(G128), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n1149), .C2(new_n821), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n848), .A2(new_n835), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n849), .C2(G124), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1217), .B(new_n1228), .C1(KEYINPUT58), .C2(new_n1215), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1208), .B1(new_n1229), .B2(new_n793), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1201), .B2(new_n791), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1206), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1173), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1182), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1205), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1205), .A3(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n738), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1237), .B2(KEYINPUT125), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT125), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1236), .A2(new_n1239), .A3(new_n738), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1232), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(G375));
  INV_X1    g1042(.A(new_n1003), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1177), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1180), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n783), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1124), .A2(new_n790), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n803), .B1(G68), .B2(new_n1162), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n390), .B1(new_n834), .B2(new_n250), .C1(new_n1100), .C2(new_n831), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n842), .B2(G128), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n806), .A2(new_n876), .B1(new_n261), .B2(new_n808), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n813), .A2(new_n856), .B1(new_n825), .B2(new_n1152), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G132), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1250), .B(new_n1253), .C1(new_n1254), .C2(new_n821), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n806), .A2(new_n880), .B1(new_n504), .B2(new_n825), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1049), .B(new_n1256), .C1(G107), .C2(new_n809), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1022), .B(new_n288), .C1(G97), .C2(new_n832), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n494), .C2(new_n841), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n821), .A2(new_n811), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1255), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1248), .B1(new_n1261), .B2(new_n793), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1246), .B1(new_n1247), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1245), .A2(new_n1263), .ZN(G381));
  AOI211_X1 g1064(.A(new_n1168), .B(new_n1144), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(G375), .A2(new_n1266), .ZN(new_n1267));
  OR2_X1    g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(G390), .A2(new_n1268), .A3(G384), .A4(G381), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1267), .A2(new_n1018), .A3(new_n1046), .A4(new_n1269), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n721), .A2(G213), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1267), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(G407), .A2(G213), .A3(new_n1273), .ZN(G409));
  NAND3_X1  g1074(.A1(new_n872), .A2(KEYINPUT126), .A3(new_n892), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1263), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1180), .A2(KEYINPUT60), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1278), .A2(new_n1244), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n738), .B1(new_n1278), .B2(new_n1244), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1277), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G384), .A2(new_n1282), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1277), .B(new_n1284), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1183), .B(new_n1232), .C1(new_n1238), .C2(new_n1240), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1232), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1234), .A2(new_n1205), .A3(new_n1243), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1290), .A2(new_n1265), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1271), .B(new_n1286), .C1(new_n1287), .C2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT62), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1272), .A2(G2897), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1286), .B(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1291), .B1(new_n1241), .B2(G378), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1272), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1237), .A2(KEYINPUT125), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1235), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1240), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(G378), .A3(new_n1288), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1290), .A2(new_n1265), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1271), .A4(new_n1286), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1293), .A2(new_n1294), .A3(new_n1298), .A4(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT127), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(G390), .A2(new_n1018), .A3(new_n1046), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1018), .B2(new_n1046), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(G396), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1310), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1312), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G387), .A2(new_n1117), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1314), .B1(new_n1315), .B2(new_n1309), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1308), .B1(new_n1313), .B2(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1312), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1315), .A2(new_n1314), .A3(new_n1309), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(KEYINPUT127), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1307), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1304), .A2(new_n1271), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1323), .B2(new_n1296), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1304), .A2(KEYINPUT63), .A3(new_n1271), .A4(new_n1286), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1292), .A2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1322), .A2(new_n1329), .ZN(G405));
  NAND2_X1  g1130(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1302), .B1(new_n1241), .B2(new_n1266), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1331), .A2(new_n1333), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1286), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1321), .A2(new_n1332), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1338), .A2(new_n1283), .A3(new_n1285), .A4(new_n1334), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(G402));
endmodule


