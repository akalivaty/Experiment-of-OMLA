//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1307, new_n1308;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI21_X1  g0005(.A(G50), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  AND2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT66), .Z(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G68), .A2(G238), .ZN(new_n214));
  AND3_X1   g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n211), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NAND2_X1  g0021(.A1(new_n204), .A2(new_n205), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n216), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT65), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n228), .B1(new_n219), .B2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G13), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n230), .A2(KEYINPUT65), .A3(G1), .A4(G20), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n232), .B(G250), .C1(G257), .C2(G264), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g0034(.A1(new_n221), .A2(new_n227), .A3(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G264), .ZN(new_n243));
  INV_X1    g0043(.A(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G87), .B(G97), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(G107), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(new_n217), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n254), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G223), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G77), .ZN(new_n273));
  INV_X1    g0073(.A(G222), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n266), .A2(new_n267), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT68), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n269), .B(new_n273), .C1(new_n274), .C2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n256), .ZN(new_n282));
  AOI211_X1 g0082(.A(new_n260), .B(new_n263), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G179), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(G20), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G150), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n225), .A2(G33), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT8), .B(G58), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n287), .B1(new_n288), .B2(new_n289), .C1(new_n206), .C2(new_n225), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n224), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n290), .A2(new_n292), .B1(new_n216), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n292), .B1(new_n257), .B2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G50), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n285), .B(new_n298), .C1(G169), .C2(new_n283), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n281), .A2(new_n282), .ZN(new_n301));
  INV_X1    g0101(.A(new_n260), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(new_n302), .A3(new_n262), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G200), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n304), .A2(KEYINPUT72), .B1(G190), .B2(new_n283), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n298), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n283), .A2(KEYINPUT72), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n290), .A2(new_n292), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n294), .A2(new_n216), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n310), .A2(KEYINPUT9), .A3(new_n311), .A4(new_n297), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT71), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n295), .A2(KEYINPUT71), .A3(KEYINPUT9), .A4(new_n297), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n305), .A2(new_n307), .A3(new_n309), .A4(new_n316), .ZN(new_n317));
  OR2_X1    g0117(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(KEYINPUT10), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n300), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n266), .A2(new_n225), .A3(new_n267), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n272), .A2(KEYINPUT73), .A3(KEYINPUT7), .A4(new_n225), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(G68), .A3(new_n327), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(G20), .B1(G159), .B2(new_n286), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT16), .ZN(new_n332));
  INV_X1    g0132(.A(new_n330), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n203), .B1(new_n323), .B2(new_n324), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n331), .A2(new_n292), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n289), .A2(new_n293), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n296), .B2(new_n289), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n256), .A2(G232), .A3(new_n258), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n262), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n268), .A2(G226), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n275), .A2(new_n279), .A3(G223), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G87), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n341), .B1(new_n345), .B2(new_n282), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT74), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n340), .A2(new_n262), .A3(KEYINPUT74), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n349), .A2(new_n350), .B1(new_n345), .B2(new_n282), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n308), .A2(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT17), .B1(new_n339), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n338), .ZN(new_n355));
  INV_X1    g0155(.A(new_n292), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n321), .A2(new_n322), .ZN(new_n357));
  AOI21_X1  g0157(.A(KEYINPUT7), .B1(new_n272), .B2(new_n225), .ZN(new_n358));
  OAI21_X1  g0158(.A(G68), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n330), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n356), .B1(new_n360), .B2(new_n332), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n355), .B1(new_n361), .B2(new_n331), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT17), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n349), .A2(new_n350), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n345), .A2(new_n282), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI22_X1  g0166(.A1(new_n366), .A2(G190), .B1(G200), .B2(new_n346), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n362), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n354), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n347), .B1(new_n351), .B2(new_n284), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n339), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n366), .A2(G179), .B1(G169), .B2(new_n346), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n362), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n276), .A2(new_n278), .B1(new_n266), .B2(new_n267), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(G232), .B1(new_n268), .B2(G238), .ZN(new_n379));
  INV_X1    g0179(.A(G107), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(new_n275), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n282), .ZN(new_n382));
  INV_X1    g0182(.A(new_n259), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G244), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n262), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n370), .ZN(new_n386));
  XNOR2_X1  g0186(.A(new_n289), .B(KEYINPUT69), .ZN(new_n387));
  INV_X1    g0187(.A(new_n286), .ZN(new_n388));
  XOR2_X1   g0188(.A(KEYINPUT15), .B(G87), .Z(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n387), .A2(new_n388), .B1(new_n390), .B2(new_n288), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n225), .A2(new_n207), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n292), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n294), .A2(new_n207), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n296), .A2(G77), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n382), .A2(new_n284), .A3(new_n262), .A4(new_n384), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n386), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n377), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n385), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G190), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT70), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n385), .A2(G200), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n393), .A2(KEYINPUT70), .A3(new_n394), .A4(new_n395), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n402), .A2(new_n404), .A3(new_n405), .A4(new_n406), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n275), .A2(new_n279), .A3(G226), .ZN(new_n408));
  OAI211_X1 g0208(.A(G232), .B(G1698), .C1(new_n270), .C2(new_n271), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n282), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n383), .A2(G238), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n262), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT13), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n412), .A2(new_n416), .A3(new_n262), .A4(new_n413), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT14), .B1(new_n418), .B2(new_n370), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(G179), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n417), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT14), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n422), .A3(G169), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n203), .A2(G20), .ZN(new_n425));
  OAI221_X1 g0225(.A(new_n425), .B1(new_n288), .B2(new_n207), .C1(new_n388), .C2(new_n216), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n426), .A2(KEYINPUT11), .A3(new_n292), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n296), .A2(G68), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n293), .A2(G68), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT12), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT11), .B1(new_n426), .B2(new_n292), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n418), .A2(G190), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n421), .B2(G200), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n424), .A2(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n320), .A2(new_n400), .A3(new_n407), .A4(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n257), .A2(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n261), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n275), .A2(new_n279), .A3(G238), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n275), .A2(G244), .A3(G1698), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G116), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n440), .B1(new_n444), .B2(new_n282), .ZN(new_n445));
  AND2_X1   g0245(.A1(G33), .A2(G41), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n439), .B(G250), .C1(new_n446), .C2(new_n224), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT78), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n256), .A2(KEYINPUT78), .A3(G250), .A4(new_n439), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(G169), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  AOI221_X4 g0252(.A(new_n440), .B1(new_n449), .B2(new_n450), .C1(new_n444), .C2(new_n282), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n452), .B1(new_n284), .B2(new_n453), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n410), .A2(KEYINPUT19), .A3(G20), .ZN(new_n455));
  INV_X1    g0255(.A(G87), .ZN(new_n456));
  INV_X1    g0256(.A(G97), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n457), .A3(new_n380), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n410), .A2(new_n225), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n455), .B1(new_n460), .B2(KEYINPUT19), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n225), .B(G68), .C1(new_n270), .C2(new_n271), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT79), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT79), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT19), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n458), .B2(new_n459), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n465), .B(new_n462), .C1(new_n467), .C2(new_n455), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n464), .A2(new_n292), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n390), .A2(new_n294), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n389), .B(KEYINPUT80), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n356), .B(new_n293), .C1(G1), .C2(new_n254), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n472), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G87), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n469), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n445), .A2(new_n352), .A3(new_n451), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n453), .B2(G200), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n454), .A2(new_n473), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT77), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(KEYINPUT5), .A2(G41), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n439), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G274), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n257), .B(G45), .C1(new_n486), .C2(new_n481), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n256), .ZN(new_n488));
  INV_X1    g0288(.A(G257), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OR2_X1    g0290(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(KEYINPUT76), .A2(KEYINPUT4), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G244), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(new_n280), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n275), .A2(new_n279), .A3(G244), .A4(new_n491), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n268), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI211_X1 g0298(.A(new_n480), .B(new_n490), .C1(new_n498), .C2(new_n282), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n275), .A2(G250), .A3(G1698), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n378), .A2(G244), .B1(new_n491), .B2(new_n492), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n282), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n490), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT77), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(G190), .B1(new_n499), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n472), .A2(new_n457), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n293), .A2(G97), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT75), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n380), .B1(new_n323), .B2(new_n324), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT6), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n457), .A2(new_n380), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G97), .A2(G107), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n380), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n225), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n388), .A2(new_n207), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n512), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n509), .B(new_n511), .C1(new_n520), .C2(new_n356), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n308), .B1(new_n504), .B2(new_n505), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n507), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n504), .A2(new_n505), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n480), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n504), .A2(KEYINPUT77), .A3(new_n505), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n370), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n357), .B2(new_n358), .ZN(new_n529));
  INV_X1    g0329(.A(new_n518), .ZN(new_n530));
  INV_X1    g0330(.A(new_n519), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n508), .B1(new_n532), .B2(new_n292), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n490), .B1(new_n498), .B2(new_n282), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n511), .B1(new_n284), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT83), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT25), .ZN(new_n538));
  AOI211_X1 g0338(.A(G107), .B(new_n293), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n537), .A2(new_n538), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n474), .A2(G107), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT24), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n225), .B(G87), .C1(new_n270), .C2(new_n271), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT22), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n275), .A2(new_n548), .A3(new_n225), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n443), .A2(G20), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n225), .A2(G107), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT23), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n545), .A2(new_n550), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n547), .B2(new_n549), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n545), .B1(new_n556), .B2(new_n554), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n292), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n487), .A2(G264), .A3(new_n256), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT84), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n487), .A2(new_n561), .A3(G264), .A4(new_n256), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n275), .A2(new_n279), .A3(G250), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n275), .A2(G257), .A3(G1698), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G294), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n560), .A2(new_n562), .B1(new_n566), .B2(new_n282), .ZN(new_n567));
  AOI21_X1  g0367(.A(G200), .B1(new_n567), .B2(new_n485), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n560), .A2(new_n562), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n282), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n352), .A2(new_n569), .A3(new_n570), .A4(new_n485), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n544), .B(new_n558), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n479), .A2(new_n524), .A3(new_n536), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(new_n284), .A3(new_n485), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n569), .A2(new_n570), .A3(new_n485), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n370), .ZN(new_n576));
  AOI21_X1  g0376(.A(G20), .B1(new_n266), .B2(new_n267), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n548), .B1(new_n577), .B2(G87), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n546), .A2(KEYINPUT22), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n552), .B(new_n554), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT24), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n556), .A2(new_n545), .A3(new_n554), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n356), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n574), .B(new_n576), .C1(new_n583), .C2(new_n543), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n268), .A2(G264), .B1(new_n272), .B2(G303), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n378), .A2(G257), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n256), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n485), .B1(new_n488), .B2(new_n244), .ZN(new_n588));
  OAI211_X1 g0388(.A(KEYINPUT21), .B(G169), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n280), .A2(new_n489), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n275), .A2(G264), .A3(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n272), .A2(G303), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n282), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n484), .A2(new_n282), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(G270), .B1(G274), .B2(new_n484), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(G179), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n294), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n472), .B2(new_n599), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(G20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n292), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n292), .A2(KEYINPUT81), .A3(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n500), .B(new_n225), .C1(G33), .C2(new_n457), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT20), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n292), .A2(KEYINPUT81), .A3(new_n603), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT81), .B1(new_n292), .B2(new_n603), .ZN(new_n612));
  OAI211_X1 g0412(.A(KEYINPUT20), .B(new_n609), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n602), .B1(new_n610), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n598), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n370), .B1(new_n594), .B2(new_n596), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XOR2_X1   g0418(.A(KEYINPUT82), .B(KEYINPUT21), .Z(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n608), .A2(new_n609), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n601), .B1(new_n623), .B2(new_n613), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n587), .A2(new_n588), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(G190), .ZN(new_n626));
  OAI21_X1  g0426(.A(G200), .B1(new_n587), .B2(new_n588), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n624), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n584), .A2(new_n616), .A3(new_n620), .A4(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n438), .A2(new_n573), .A3(new_n629), .ZN(G372));
  INV_X1    g0430(.A(KEYINPUT10), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n317), .B(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n422), .B1(new_n421), .B2(G169), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT14), .B(new_n370), .C1(new_n415), .C2(new_n417), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n433), .B1(new_n635), .B2(new_n420), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n398), .B1(new_n435), .B2(new_n436), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n369), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n632), .B1(new_n638), .B2(new_n376), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT86), .B1(new_n639), .B2(new_n300), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT86), .ZN(new_n641));
  INV_X1    g0441(.A(new_n376), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n424), .A2(new_n434), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n435), .A2(new_n436), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n399), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n642), .B1(new_n646), .B2(new_n369), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n641), .B(new_n299), .C1(new_n647), .C2(new_n632), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n438), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n528), .A2(new_n535), .A3(KEYINPUT85), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT85), .B1(new_n528), .B2(new_n535), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n651), .B(new_n479), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n445), .A2(new_n451), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n370), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n473), .B(new_n656), .C1(G179), .C2(new_n655), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n478), .A2(new_n476), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n572), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n528), .A2(new_n535), .B1(new_n507), .B2(new_n523), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n618), .A2(new_n619), .B1(new_n598), .B2(new_n615), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n584), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n658), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT26), .B1(new_n664), .B2(new_n536), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n654), .A2(new_n663), .A3(new_n657), .A4(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n650), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n649), .A2(new_n667), .ZN(G369));
  INV_X1    g0468(.A(new_n661), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n230), .A2(G20), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n257), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT27), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n672), .A2(G213), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G343), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n615), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n628), .A2(new_n677), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n661), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT87), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT87), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n676), .B1(new_n583), .B2(new_n543), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n572), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n584), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n584), .A2(new_n676), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n684), .A2(G330), .A3(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n661), .A2(new_n676), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n688), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(G399));
  INV_X1    g0495(.A(new_n232), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G41), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n257), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n458), .A2(G116), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n698), .A2(new_n699), .B1(new_n223), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT28), .Z(new_n701));
  INV_X1    g0501(.A(new_n629), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(new_n659), .A3(new_n660), .A4(new_n675), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n526), .A2(new_n527), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n597), .A2(new_n655), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n567), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n704), .A2(KEYINPUT30), .A3(new_n567), .A4(new_n705), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n525), .A2(new_n575), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n625), .A2(G179), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(new_n655), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT88), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n710), .A2(KEYINPUT88), .A3(new_n655), .A4(new_n711), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n708), .A2(new_n709), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n703), .A2(KEYINPUT31), .B1(new_n676), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n708), .A2(new_n709), .A3(new_n712), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n479), .B1(new_n652), .B2(new_n653), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT26), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n479), .A2(new_n651), .A3(new_n528), .A4(new_n535), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n725), .A2(new_n657), .A3(new_n663), .A4(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n723), .B1(new_n727), .B2(new_n675), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n666), .A2(new_n723), .A3(new_n675), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n722), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n701), .B1(new_n730), .B2(G1), .ZN(G364));
  AOI21_X1  g0531(.A(new_n257), .B1(new_n670), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n697), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n224), .B1(G20), .B2(new_n370), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G179), .A2(G200), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n225), .B1(new_n738), .B2(G190), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G294), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n225), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(new_n738), .ZN(new_n746));
  INV_X1    g0546(.A(G329), .ZN(new_n747));
  INV_X1    g0547(.A(G303), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n308), .A2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G20), .A3(G190), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n272), .B1(new_n746), .B2(new_n747), .C1(new_n748), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(G20), .A2(G179), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT92), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G190), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n308), .ZN(new_n755));
  XNOR2_X1  g0555(.A(KEYINPUT96), .B(G326), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n745), .A2(new_n749), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n754), .A2(G200), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n744), .B(new_n760), .C1(G322), .C2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n753), .A2(new_n352), .A3(new_n308), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n753), .A2(new_n352), .A3(G200), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(KEYINPUT94), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT33), .B(G317), .Z(new_n769));
  OAI221_X1 g0569(.A(new_n762), .B1(new_n763), .B2(new_n764), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n759), .A2(new_n380), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n275), .B1(new_n750), .B2(new_n456), .ZN(new_n772));
  INV_X1    g0572(.A(new_n768), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n771), .B(new_n772), .C1(new_n773), .C2(G68), .ZN(new_n774));
  INV_X1    g0574(.A(new_n764), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G50), .A2(new_n755), .B1(new_n775), .B2(G77), .ZN(new_n776));
  INV_X1    g0576(.A(new_n761), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n202), .B2(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT93), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT93), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n742), .A2(new_n457), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT32), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n746), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n746), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(KEYINPUT32), .A3(G159), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n781), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n774), .A2(new_n779), .A3(new_n780), .A4(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n737), .B1(new_n770), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT90), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n225), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT91), .Z(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n736), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n249), .A2(G45), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n696), .A2(new_n275), .ZN(new_n797));
  INV_X1    g0597(.A(new_n223), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n797), .C1(G45), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n232), .A2(G355), .A3(new_n275), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n799), .B(new_n800), .C1(G116), .C2(new_n232), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n735), .B(new_n789), .C1(new_n795), .C2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n684), .B2(new_n793), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n684), .A2(G330), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n735), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n684), .A2(G330), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT89), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n804), .B1(new_n806), .B2(new_n808), .ZN(G396));
  NAND2_X1  g0609(.A1(new_n666), .A2(new_n675), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n398), .A2(new_n676), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n396), .A2(new_n676), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n407), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(new_n813), .B2(new_n398), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n666), .A2(new_n675), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(new_n722), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n735), .ZN(new_n820));
  INV_X1    g0620(.A(new_n755), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n743), .A2(new_n777), .B1(new_n821), .B2(new_n748), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n272), .B1(new_n746), .B2(new_n763), .C1(new_n380), .C2(new_n750), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n759), .A2(new_n456), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n822), .A2(new_n781), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n825), .B1(new_n599), .B2(new_n764), .C1(new_n758), .C2(new_n768), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G137), .A2(new_n755), .B1(new_n761), .B2(G143), .ZN(new_n827));
  INV_X1    g0627(.A(G150), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n783), .B2(new_n764), .C1(new_n768), .C2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT34), .ZN(new_n830));
  INV_X1    g0630(.A(G132), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n275), .B1(new_n746), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n750), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G50), .B2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n830), .B(new_n834), .C1(new_n202), .C2(new_n742), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n759), .A2(new_n203), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n826), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n736), .A2(new_n790), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n837), .A2(new_n736), .B1(new_n207), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n815), .A2(new_n791), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n839), .A2(new_n734), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n820), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(KEYINPUT103), .ZN(new_n843));
  AND3_X1   g0643(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n717), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n716), .A2(KEYINPUT31), .A3(new_n676), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT31), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n524), .A2(new_n536), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n572), .A2(new_n657), .A3(new_n658), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n848), .A2(new_n629), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n850), .B2(new_n675), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n716), .A2(new_n676), .ZN(new_n852));
  OAI211_X1 g0652(.A(KEYINPUT103), .B(new_n846), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n332), .A2(KEYINPUT100), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n328), .A2(new_n330), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n328), .B2(new_n330), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n856), .A2(new_n857), .A3(new_n356), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n674), .B1(new_n858), .B2(new_n355), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n371), .B1(new_n858), .B2(new_n355), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n362), .A2(new_n367), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n339), .A2(new_n353), .ZN(new_n864));
  INV_X1    g0664(.A(new_n674), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n374), .A2(new_n865), .B1(new_n336), .B2(new_n338), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n863), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n859), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n377), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT102), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n339), .A2(KEYINPUT17), .A3(new_n353), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n363), .B1(new_n362), .B2(new_n367), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n354), .A2(KEYINPUT102), .A3(new_n368), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n878), .A2(new_n376), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n362), .A2(new_n865), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n868), .B1(new_n864), .B2(new_n866), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n880), .A2(new_n881), .B1(new_n870), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n874), .B1(new_n883), .B2(KEYINPUT38), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT99), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n643), .B2(new_n675), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n636), .A2(KEYINPUT99), .A3(new_n676), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n434), .A2(new_n676), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n886), .A2(new_n887), .B1(new_n437), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n854), .A2(new_n814), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n815), .B(new_n889), .C1(new_n845), .C2(new_n853), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n871), .B2(new_n873), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT40), .B1(new_n894), .B2(new_n874), .ZN(new_n895));
  AOI22_X1  g0695(.A1(KEYINPUT40), .A2(new_n891), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT104), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n854), .A2(new_n650), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n897), .B(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(G330), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n862), .A2(KEYINPUT37), .B1(new_n867), .B2(new_n869), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n859), .B1(new_n369), .B2(new_n376), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT39), .B1(new_n893), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT39), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n874), .B(new_n906), .C1(new_n883), .C2(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n643), .A2(new_n676), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n376), .A2(new_n674), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n811), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n817), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n914), .B(new_n890), .C1(new_n904), .C2(new_n893), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n650), .B1(new_n728), .B2(new_n729), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n649), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n900), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n257), .B2(new_n670), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n516), .A2(new_n517), .ZN(new_n922));
  OAI211_X1 g0722(.A(G116), .B(new_n226), .C1(new_n922), .C2(KEYINPUT35), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT98), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(KEYINPUT35), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  OAI21_X1  g0727(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n798), .A2(new_n928), .B1(G50), .B2(new_n203), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(G1), .A3(new_n230), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n921), .A2(new_n927), .A3(new_n930), .ZN(G367));
  INV_X1    g0731(.A(G317), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n272), .B1(new_n932), .B2(new_n746), .C1(new_n821), .C2(new_n763), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n759), .A2(new_n457), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n750), .A2(new_n599), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT46), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n742), .A2(new_n380), .B1(new_n758), .B2(new_n764), .ZN(new_n937));
  NOR4_X1   g0737(.A1(new_n933), .A2(new_n934), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n938), .B1(new_n743), .B2(new_n768), .C1(new_n748), .C2(new_n777), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n742), .A2(new_n203), .ZN(new_n940));
  INV_X1    g0740(.A(G137), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n750), .A2(new_n202), .B1(new_n746), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT109), .ZN(new_n943));
  INV_X1    g0743(.A(new_n759), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n272), .B(new_n943), .C1(G77), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n755), .A2(G143), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n777), .B2(new_n828), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G50), .B2(new_n775), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n945), .B(new_n948), .C1(new_n783), .C2(new_n768), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n939), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT47), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n735), .B1(new_n951), .B2(new_n736), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n476), .A2(new_n675), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n473), .A3(new_n454), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n664), .B2(new_n953), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n793), .ZN(new_n956));
  INV_X1    g0756(.A(new_n797), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n795), .B1(new_n232), .B2(new_n390), .C1(new_n245), .C2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n952), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n536), .A2(KEYINPUT105), .A3(new_n675), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n521), .A2(new_n676), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n660), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(KEYINPUT105), .B1(new_n536), .B2(new_n675), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n692), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n970));
  INV_X1    g0770(.A(new_n584), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n536), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT106), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n972), .A2(KEYINPUT106), .A3(new_n536), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n675), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n687), .A2(new_n689), .A3(new_n693), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n970), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT42), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n977), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n968), .A2(new_n969), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n968), .B1(new_n983), .B2(new_n969), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n961), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n969), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n967), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n960), .A3(new_n984), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT108), .ZN(new_n992));
  INV_X1    g0792(.A(new_n694), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n966), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT108), .B1(new_n970), .B2(new_n694), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n970), .A2(new_n694), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n692), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n690), .B1(new_n661), .B2(new_n676), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n805), .A2(new_n978), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n978), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n684), .A2(new_n1008), .A3(G330), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n998), .A2(new_n692), .A3(new_n1002), .A4(new_n999), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1005), .A2(new_n730), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n730), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n697), .B(KEYINPUT41), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n733), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n959), .B1(new_n991), .B2(new_n1015), .ZN(G387));
  NAND2_X1  g0816(.A1(new_n1010), .A2(new_n733), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT110), .Z(new_n1018));
  NOR2_X1   g0818(.A1(new_n387), .A2(G50), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n699), .B1(new_n203), .B2(new_n207), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1021), .A2(new_n1022), .A3(G45), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n957), .B1(new_n241), .B2(G45), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n696), .A2(new_n272), .A3(new_n699), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1024), .A2(new_n1027), .B1(G107), .B2(new_n232), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n690), .A2(new_n794), .B1(new_n795), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G322), .A2(new_n755), .B1(new_n775), .B2(G303), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n932), .B2(new_n777), .C1(new_n768), .C2(new_n763), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT48), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n758), .B2(new_n742), .C1(new_n743), .C2(new_n750), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT49), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n785), .A2(new_n756), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(KEYINPUT49), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n275), .B1(new_n944), .B2(G116), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n471), .A2(new_n742), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n275), .B1(new_n759), .B2(new_n457), .C1(new_n207), .C2(new_n750), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n761), .B2(G50), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n828), .B2(new_n746), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1040), .B(new_n1043), .C1(G68), .C2(new_n775), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n783), .B2(new_n821), .C1(new_n289), .C2(new_n768), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n734), .B(new_n1029), .C1(new_n1046), .C2(new_n737), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1010), .B(new_n730), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n697), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1018), .B(new_n1047), .C1(new_n1048), .C2(new_n1049), .ZN(G393));
  NAND3_X1  g0850(.A1(new_n1005), .A2(KEYINPUT111), .A3(new_n1011), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1011), .A2(KEYINPUT111), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1010), .A2(new_n730), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(KEYINPUT116), .A4(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1054), .A2(new_n1012), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1053), .A3(new_n1052), .ZN(new_n1056));
  INV_X1    g0856(.A(KEYINPUT116), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1049), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n733), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n795), .B1(new_n457), .B2(new_n232), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n252), .B2(new_n797), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT113), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n275), .B(new_n771), .C1(G322), .C2(new_n785), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n599), .B2(new_n742), .C1(new_n743), .C2(new_n764), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G303), .B2(new_n773), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G311), .A2(new_n761), .B1(new_n755), .B2(G317), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(new_n758), .C2(new_n750), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G150), .A2(new_n755), .B1(new_n761), .B2(G159), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT51), .Z(new_n1072));
  OR2_X1    g0872(.A1(new_n387), .A2(new_n764), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n773), .A2(G50), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n833), .A2(G68), .B1(new_n785), .B2(G143), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n275), .B1(new_n1075), .B2(KEYINPUT114), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n742), .A2(new_n207), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .A4(new_n824), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n737), .B1(new_n1070), .B2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1064), .A2(new_n735), .A3(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT115), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n966), .A2(new_n794), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT112), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1059), .A2(new_n1061), .A3(new_n1086), .ZN(G390));
  NAND3_X1  g0887(.A1(new_n905), .A2(new_n907), .A3(new_n791), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n838), .A2(new_n289), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n777), .A2(new_n599), .B1(new_n457), .B2(new_n764), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n272), .B1(new_n746), .B2(new_n743), .C1(new_n456), .C2(new_n750), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1090), .A2(new_n836), .A3(new_n1078), .A4(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1092), .B1(new_n380), .B2(new_n768), .C1(new_n758), .C2(new_n821), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT119), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  AOI22_X1  g0895(.A1(new_n773), .A2(G137), .B1(new_n775), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n783), .B2(new_n742), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1097), .A2(KEYINPUT117), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n785), .A2(G125), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(KEYINPUT117), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G128), .A2(new_n755), .B1(new_n761), .B2(G132), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT118), .Z(new_n1102));
  AND3_X1   g0902(.A1(new_n833), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1103));
  AOI21_X1  g0903(.A(KEYINPUT53), .B1(new_n833), .B2(G150), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n275), .B1(new_n216), .B2(new_n759), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1094), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n735), .B1(new_n1108), .B2(new_n736), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1088), .A2(new_n1089), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n909), .B1(new_n914), .B2(new_n890), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n813), .A2(new_n398), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n727), .A2(new_n675), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n889), .B1(new_n1114), .B2(new_n913), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n909), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n884), .A2(new_n1116), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1112), .A2(new_n908), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n854), .A2(G330), .A3(new_n814), .A4(new_n890), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(G330), .B(new_n814), .C1(new_n717), .C2(new_n719), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n889), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n1115), .B2(new_n1117), .C1(new_n1112), .C2(new_n908), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1111), .B1(new_n1124), .B2(new_n733), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n649), .B(new_n917), .C1(new_n898), .C2(new_n721), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1121), .A2(new_n889), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1119), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n914), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n716), .A2(new_n676), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n573), .A2(new_n629), .A3(new_n676), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n847), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT103), .B1(new_n1132), .B2(new_n846), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n717), .A2(new_n844), .A3(new_n843), .ZN(new_n1134));
  OAI211_X1 g0934(.A(G330), .B(new_n814), .C1(new_n1133), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n889), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n913), .B(new_n1114), .C1(new_n1121), .C2(new_n889), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1126), .B1(new_n1129), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n697), .B1(new_n1140), .B2(new_n1124), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n721), .B(new_n438), .C1(new_n845), .C2(new_n853), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n918), .A2(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1119), .A2(new_n1127), .B1(new_n913), .B2(new_n817), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1137), .B1(new_n1135), .B2(new_n889), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1125), .B1(new_n1141), .B2(new_n1148), .ZN(G378));
  OAI21_X1  g0949(.A(new_n916), .B1(new_n896), .B2(new_n721), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n891), .A2(KEYINPUT40), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n892), .A2(new_n895), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(G330), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n298), .A2(new_n674), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n320), .B(new_n1156), .Z(new_n1157));
  INV_X1    g0957(.A(KEYINPUT55), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1159), .A2(KEYINPUT56), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(KEYINPUT56), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1150), .A2(new_n1155), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1163), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n733), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n791), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n838), .A2(new_n216), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n821), .A2(new_n599), .B1(new_n471), .B2(new_n764), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G58), .A2(new_n944), .B1(new_n785), .B2(G283), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n207), .B2(new_n750), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n272), .A2(new_n255), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n1169), .A2(new_n1171), .A3(new_n940), .A4(new_n1172), .ZN(new_n1173));
  OAI221_X1 g0973(.A(new_n1173), .B1(new_n457), .B2(new_n768), .C1(new_n380), .C2(new_n777), .ZN(new_n1174));
  XOR2_X1   g0974(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n216), .B1(new_n270), .B2(G41), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(new_n785), .B2(G124), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1178), .B(new_n254), .C1(new_n783), .C2(new_n759), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT121), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n742), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1181), .A2(G150), .B1(new_n755), .B2(G125), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n761), .A2(G128), .B1(new_n833), .B2(new_n1095), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n831), .B2(new_n768), .C1(new_n941), .C2(new_n764), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT59), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1176), .B(new_n1177), .C1(new_n1180), .C2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n735), .B1(new_n1187), .B2(new_n736), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1167), .A2(new_n1168), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1166), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n896), .A2(new_n916), .A3(new_n721), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1154), .B1(new_n1153), .B2(G330), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1150), .A2(new_n1155), .A3(new_n1163), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1140), .A2(new_n1124), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1195), .A2(new_n1196), .B1(new_n1144), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n697), .B1(new_n1198), .B2(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1144), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1191), .B1(new_n1199), .B2(new_n1203), .ZN(G375));
  NOR3_X1   g1004(.A1(new_n1145), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(new_n1014), .A3(new_n1147), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n773), .A2(G116), .B1(G107), .B2(new_n775), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n743), .B2(new_n821), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT123), .Z(new_n1210));
  OAI221_X1 g1010(.A(new_n272), .B1(new_n746), .B2(new_n748), .C1(new_n207), .C2(new_n759), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1211), .B(new_n1040), .C1(G283), .C2(new_n761), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1210), .B(new_n1212), .C1(new_n457), .C2(new_n750), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n742), .A2(new_n216), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n275), .B1(new_n759), .B2(new_n202), .C1(new_n783), .C2(new_n750), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n777), .A2(new_n941), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G128), .C2(new_n785), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n773), .A2(new_n1095), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G132), .A2(new_n755), .B1(new_n775), .B2(G150), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1213), .B1(new_n1214), .B2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1221), .A2(new_n736), .B1(new_n203), .B2(new_n838), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n889), .A2(new_n790), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT122), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1223), .A2(KEYINPUT122), .ZN(new_n1226));
  NOR3_X1   g1026(.A1(new_n1225), .A2(new_n735), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1129), .A2(new_n1139), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n733), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1207), .A2(new_n1229), .ZN(G381));
  AOI21_X1  g1030(.A(new_n1049), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1198), .A2(KEYINPUT57), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n732), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1189), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1234), .A2(G378), .A3(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1238), .A2(G390), .A3(G384), .A4(G387), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1237), .A2(new_n1229), .A3(new_n1207), .A4(new_n1239), .ZN(G407));
  INV_X1    g1040(.A(new_n1237), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G343), .C2(new_n1241), .ZN(G409));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(G343), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1198), .A2(new_n1014), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1244), .B1(new_n1236), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1190), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1247));
  INV_X1    g1047(.A(G378), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n697), .B1(new_n1205), .B2(KEYINPUT60), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1129), .A2(new_n1139), .A3(KEYINPUT60), .A4(new_n1126), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1147), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1229), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(G384), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G384), .B(new_n1229), .C1(new_n1250), .C2(new_n1252), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT124), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(KEYINPUT124), .A3(new_n1256), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1244), .A2(G2897), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1259), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1255), .A2(KEYINPUT124), .A3(new_n1256), .A4(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1257), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT61), .B1(new_n1249), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1246), .B(new_n1266), .C1(new_n1247), .C2(new_n1248), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(KEYINPUT62), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G375), .A2(G378), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT62), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1269), .A2(new_n1270), .A3(new_n1266), .A4(new_n1246), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1264), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n959), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n991), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1015), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(G390), .A2(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1055), .A2(new_n1058), .B1(new_n1085), .B2(new_n1083), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G387), .B1(new_n1278), .B2(new_n1061), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G393), .A2(G396), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G390), .A2(new_n1276), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1280), .A2(new_n1238), .A3(new_n1281), .A4(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT125), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1238), .B(new_n1281), .C1(new_n1279), .C2(new_n1285), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G390), .B(new_n1276), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1284), .A2(new_n1288), .A3(KEYINPUT126), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1249), .B2(new_n1263), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1267), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1284), .B(new_n1288), .C1(new_n1267), .C2(new_n1295), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1272), .A2(new_n1293), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT127), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1264), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1303), .B(new_n1304), .C1(new_n1299), .C2(new_n1298), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1301), .A2(new_n1305), .ZN(G405));
  NAND2_X1  g1106(.A1(new_n1241), .A2(new_n1269), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1307), .B(new_n1265), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1289), .ZN(G402));
endmodule


