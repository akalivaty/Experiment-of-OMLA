

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741;

  XOR2_X1 U364 ( .A(n711), .B(KEYINPUT121), .Z(n712) );
  XNOR2_X1 U365 ( .A(n431), .B(n430), .ZN(n660) );
  NAND2_X1 U366 ( .A1(n563), .A2(n600), .ZN(n664) );
  NOR2_X1 U367 ( .A1(n680), .A2(n422), .ZN(n431) );
  XNOR2_X1 U368 ( .A(n383), .B(n484), .ZN(n612) );
  NOR2_X1 U369 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U370 ( .A1(n554), .A2(n459), .ZN(n383) );
  NOR2_X1 U371 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U372 ( .A(n420), .B(n439), .ZN(n717) );
  XNOR2_X1 U373 ( .A(G134), .B(n344), .ZN(n528) );
  BUF_X1 U374 ( .A(G107), .Z(n344) );
  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n518) );
  NAND2_X2 U376 ( .A1(n541), .A2(n396), .ZN(n402) );
  XNOR2_X1 U377 ( .A(n343), .B(n370), .ZN(n369) );
  NAND2_X1 U378 ( .A1(n356), .A2(n372), .ZN(n343) );
  XNOR2_X1 U379 ( .A(n365), .B(KEYINPUT85), .ZN(n381) );
  AND2_X2 U380 ( .A1(n415), .A2(n676), .ZN(n651) );
  INV_X1 U381 ( .A(G953), .ZN(n732) );
  NOR2_X1 U382 ( .A1(n740), .A2(KEYINPUT67), .ZN(n409) );
  XNOR2_X2 U383 ( .A(n451), .B(KEYINPUT39), .ZN(n541) );
  AND2_X2 U384 ( .A1(n423), .A2(n425), .ZN(n408) );
  NOR2_X2 U385 ( .A1(n675), .A2(n573), .ZN(n445) );
  XNOR2_X2 U386 ( .A(n446), .B(KEYINPUT21), .ZN(n675) );
  NAND2_X2 U387 ( .A1(n408), .A2(n608), .ZN(n440) );
  XNOR2_X2 U388 ( .A(n400), .B(n477), .ZN(n366) );
  INV_X1 U389 ( .A(G902), .ZN(n525) );
  NOR2_X1 U390 ( .A1(n616), .A2(n552), .ZN(n399) );
  INV_X1 U391 ( .A(n544), .ZN(n554) );
  XNOR2_X1 U392 ( .A(n354), .B(G146), .ZN(n447) );
  XNOR2_X1 U393 ( .A(G110), .B(G107), .ZN(n435) );
  XNOR2_X1 U394 ( .A(n561), .B(KEYINPUT19), .ZN(n591) );
  NOR2_X1 U395 ( .A1(n510), .A2(n589), .ZN(n573) );
  XNOR2_X1 U396 ( .A(n465), .B(n466), .ZN(n711) );
  XNOR2_X1 U397 ( .A(n717), .B(n418), .ZN(n704) );
  XNOR2_X1 U398 ( .A(n447), .B(n455), .ZN(n729) );
  XNOR2_X1 U399 ( .A(n428), .B(n426), .ZN(n439) );
  XNOR2_X1 U400 ( .A(n436), .B(n435), .ZN(n499) );
  XNOR2_X1 U401 ( .A(G104), .B(G101), .ZN(n436) );
  XNOR2_X1 U402 ( .A(KEYINPUT99), .B(KEYINPUT31), .ZN(n430) );
  XNOR2_X1 U403 ( .A(n543), .B(KEYINPUT69), .ZN(n552) );
  XNOR2_X1 U404 ( .A(KEYINPUT83), .B(KEYINPUT8), .ZN(n460) );
  INV_X1 U405 ( .A(G125), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n359), .B(n358), .ZN(n545) );
  INV_X1 U407 ( .A(KEYINPUT109), .ZN(n358) );
  NAND2_X2 U408 ( .A1(n376), .A2(n374), .ZN(n560) );
  OR2_X1 U409 ( .A1(n704), .A2(n375), .ZN(n374) );
  AND2_X1 U410 ( .A1(n378), .A2(n377), .ZN(n376) );
  XNOR2_X1 U411 ( .A(n538), .B(G478), .ZN(n571) );
  XNOR2_X1 U412 ( .A(G101), .B(G146), .ZN(n488) );
  INV_X1 U413 ( .A(G137), .ZN(n487) );
  XNOR2_X1 U414 ( .A(G134), .B(G131), .ZN(n477) );
  XNOR2_X1 U415 ( .A(n427), .B(G119), .ZN(n426) );
  XNOR2_X1 U416 ( .A(n429), .B(n491), .ZN(n428) );
  INV_X1 U417 ( .A(KEYINPUT3), .ZN(n427) );
  INV_X1 U418 ( .A(G900), .ZN(n454) );
  AND2_X1 U419 ( .A1(n619), .A2(n475), .ZN(n459) );
  XNOR2_X1 U420 ( .A(n472), .B(n471), .ZN(n597) );
  NOR2_X1 U421 ( .A1(n711), .A2(G902), .ZN(n472) );
  INV_X1 U422 ( .A(n581), .ZN(n401) );
  XNOR2_X1 U423 ( .A(n487), .B(G140), .ZN(n478) );
  XNOR2_X1 U424 ( .A(G128), .B(KEYINPUT24), .ZN(n462) );
  XOR2_X1 U425 ( .A(KEYINPUT23), .B(KEYINPUT73), .Z(n463) );
  XNOR2_X1 U426 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n455) );
  XNOR2_X1 U427 ( .A(n366), .B(n478), .ZN(n730) );
  XNOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT92), .ZN(n508) );
  INV_X1 U429 ( .A(KEYINPUT108), .ZN(n398) );
  INV_X1 U430 ( .A(KEYINPUT34), .ZN(n594) );
  NAND2_X1 U431 ( .A1(n386), .A2(n593), .ZN(n385) );
  INV_X1 U432 ( .A(KEYINPUT1), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n530), .B(n360), .ZN(n537) );
  XNOR2_X1 U434 ( .A(n531), .B(n361), .ZN(n360) );
  AND2_X1 U435 ( .A1(n630), .A2(G953), .ZN(n714) );
  XNOR2_X1 U436 ( .A(n411), .B(KEYINPUT20), .ZN(n473) );
  NAND2_X1 U437 ( .A1(n468), .A2(G234), .ZN(n411) );
  XNOR2_X1 U438 ( .A(n558), .B(n357), .ZN(n356) );
  AND2_X1 U439 ( .A1(n579), .A2(n578), .ZN(n372) );
  INV_X1 U440 ( .A(KEYINPUT46), .ZN(n357) );
  INV_X1 U441 ( .A(KEYINPUT48), .ZN(n370) );
  XNOR2_X1 U442 ( .A(G116), .B(G113), .ZN(n429) );
  INV_X1 U443 ( .A(KEYINPUT72), .ZN(n491) );
  XNOR2_X1 U444 ( .A(n467), .B(n525), .ZN(n625) );
  XNOR2_X1 U445 ( .A(KEYINPUT90), .B(KEYINPUT15), .ZN(n467) );
  XNOR2_X1 U446 ( .A(n560), .B(KEYINPUT38), .ZN(n687) );
  INV_X1 U447 ( .A(G237), .ZN(n495) );
  XNOR2_X1 U448 ( .A(G143), .B(G104), .ZN(n519) );
  XNOR2_X1 U449 ( .A(KEYINPUT11), .B(KEYINPUT100), .ZN(n513) );
  XOR2_X1 U450 ( .A(G140), .B(KEYINPUT12), .Z(n514) );
  XNOR2_X1 U451 ( .A(G113), .B(G131), .ZN(n516) );
  INV_X1 U452 ( .A(KEYINPUT107), .ZN(n397) );
  NOR2_X1 U453 ( .A1(n609), .A2(n410), .ZN(n585) );
  NAND2_X1 U454 ( .A1(n388), .A2(n459), .ZN(n609) );
  INV_X1 U455 ( .A(KEYINPUT70), .ZN(n444) );
  XNOR2_X1 U456 ( .A(n493), .B(n366), .ZN(n634) );
  XNOR2_X1 U457 ( .A(G116), .B(G122), .ZN(n531) );
  INV_X1 U458 ( .A(KEYINPUT103), .ZN(n361) );
  XOR2_X1 U459 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n529) );
  XNOR2_X1 U460 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n476) );
  XNOR2_X1 U461 ( .A(n421), .B(n499), .ZN(n420) );
  NAND2_X1 U462 ( .A1(n624), .A2(n434), .ZN(n665) );
  XNOR2_X1 U463 ( .A(n449), .B(n448), .ZN(n668) );
  INV_X1 U464 ( .A(KEYINPUT41), .ZN(n448) );
  XNOR2_X1 U465 ( .A(n610), .B(n432), .ZN(n680) );
  INV_X1 U466 ( .A(KEYINPUT98), .ZN(n432) );
  NOR2_X1 U467 ( .A1(n611), .A2(n609), .ZN(n610) );
  XNOR2_X1 U468 ( .A(n452), .B(KEYINPUT106), .ZN(n510) );
  NOR2_X1 U469 ( .A1(n587), .A2(n453), .ZN(n452) );
  NAND2_X1 U470 ( .A1(n454), .A2(G953), .ZN(n453) );
  XNOR2_X1 U471 ( .A(n527), .B(n526), .ZN(n570) );
  BUF_X1 U472 ( .A(n616), .Z(n410) );
  XNOR2_X1 U473 ( .A(n729), .B(n382), .ZN(n466) );
  XNOR2_X1 U474 ( .A(n478), .B(n348), .ZN(n382) );
  XNOR2_X1 U475 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U476 ( .A(n730), .B(n481), .ZN(n641) );
  AND2_X1 U477 ( .A1(n368), .A2(n560), .ZN(n580) );
  XNOR2_X1 U478 ( .A(n557), .B(n556), .ZN(n639) );
  INV_X1 U479 ( .A(KEYINPUT42), .ZN(n556) );
  NOR2_X1 U480 ( .A1(n668), .A2(n564), .ZN(n557) );
  XNOR2_X1 U481 ( .A(n364), .B(n363), .ZN(n563) );
  INV_X1 U482 ( .A(KEYINPUT36), .ZN(n363) );
  XNOR2_X1 U483 ( .A(KEYINPUT35), .B(KEYINPUT78), .ZN(n442) );
  XNOR2_X1 U484 ( .A(n413), .B(n412), .ZN(n741) );
  INV_X1 U485 ( .A(KEYINPUT32), .ZN(n412) );
  AND2_X1 U486 ( .A1(n457), .A2(n676), .ZN(n414) );
  NOR2_X1 U487 ( .A1(n599), .A2(n388), .ZN(n417) );
  XNOR2_X1 U488 ( .A(n708), .B(n405), .ZN(n710) );
  XNOR2_X1 U489 ( .A(n709), .B(KEYINPUT120), .ZN(n405) );
  AND2_X1 U490 ( .A1(n593), .A2(n349), .ZN(n345) );
  XOR2_X1 U491 ( .A(n665), .B(KEYINPUT81), .Z(n346) );
  AND2_X1 U492 ( .A1(n665), .A2(n404), .ZN(n347) );
  XNOR2_X1 U493 ( .A(n394), .B(n398), .ZN(n562) );
  XOR2_X1 U494 ( .A(G119), .B(G110), .Z(n348) );
  INV_X1 U495 ( .A(n565), .ZN(n396) );
  AND2_X1 U496 ( .A1(n612), .A2(n611), .ZN(n349) );
  NOR2_X1 U497 ( .A1(n688), .A2(n598), .ZN(n350) );
  XOR2_X1 U498 ( .A(KEYINPUT22), .B(KEYINPUT74), .Z(n351) );
  BUF_X1 U499 ( .A(n597), .Z(n619) );
  AND2_X1 U500 ( .A1(n567), .A2(n438), .ZN(n352) );
  XOR2_X1 U501 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n353) );
  INV_X1 U502 ( .A(KEYINPUT2), .ZN(n434) );
  XNOR2_X1 U503 ( .A(n400), .B(n419), .ZN(n418) );
  INV_X1 U504 ( .A(n646), .ZN(n424) );
  XNOR2_X2 U505 ( .A(n355), .B(n351), .ZN(n617) );
  NAND2_X1 U506 ( .A1(n593), .A2(n350), .ZN(n355) );
  NAND2_X1 U507 ( .A1(n562), .A2(n686), .ZN(n359) );
  NOR2_X1 U508 ( .A1(n597), .A2(n542), .ZN(n543) );
  NAND2_X1 U509 ( .A1(n395), .A2(n396), .ZN(n394) );
  XNOR2_X1 U510 ( .A(n417), .B(n416), .ZN(n415) );
  INV_X1 U511 ( .A(n388), .ZN(n620) );
  XNOR2_X2 U512 ( .A(n544), .B(n362), .ZN(n388) );
  NAND2_X1 U513 ( .A1(n369), .A2(n367), .ZN(n365) );
  NAND2_X1 U514 ( .A1(n562), .A2(n561), .ZN(n364) );
  NAND2_X1 U515 ( .A1(n381), .A2(n433), .ZN(n583) );
  INV_X1 U516 ( .A(n580), .ZN(n367) );
  XNOR2_X1 U517 ( .A(n546), .B(n353), .ZN(n368) );
  XNOR2_X1 U518 ( .A(n502), .B(n373), .ZN(n419) );
  XNOR2_X1 U519 ( .A(n447), .B(n501), .ZN(n373) );
  NAND2_X1 U520 ( .A1(n704), .A2(n506), .ZN(n378) );
  OR2_X1 U521 ( .A1(n404), .A2(n506), .ZN(n375) );
  NAND2_X1 U522 ( .A1(n506), .A2(n404), .ZN(n377) );
  XNOR2_X2 U523 ( .A(n548), .B(KEYINPUT111), .ZN(n438) );
  AND2_X1 U524 ( .A1(n379), .A2(G210), .ZN(n391) );
  AND2_X1 U525 ( .A1(n379), .A2(G472), .ZN(n392) );
  AND2_X1 U526 ( .A1(n379), .A2(G475), .ZN(n389) );
  AND2_X1 U527 ( .A1(n379), .A2(G217), .ZN(n390) );
  AND2_X1 U528 ( .A1(n379), .A2(n347), .ZN(n393) );
  NAND2_X1 U529 ( .A1(n346), .A2(n379), .ZN(n671) );
  XNOR2_X2 U530 ( .A(n403), .B(KEYINPUT76), .ZN(n379) );
  NAND2_X1 U531 ( .A1(n380), .A2(n639), .ZN(n558) );
  XNOR2_X1 U532 ( .A(n380), .B(G131), .ZN(G33) );
  XNOR2_X2 U533 ( .A(n402), .B(KEYINPUT40), .ZN(n380) );
  AND2_X1 U534 ( .A1(n381), .A2(n401), .ZN(n731) );
  NAND2_X1 U535 ( .A1(n450), .A2(n612), .ZN(n451) );
  NAND2_X1 U536 ( .A1(n384), .A2(n596), .ZN(n443) );
  XNOR2_X1 U537 ( .A(n385), .B(n594), .ZN(n384) );
  INV_X1 U538 ( .A(n666), .ZN(n386) );
  AND2_X1 U539 ( .A1(n620), .A2(n387), .ZN(n672) );
  INV_X1 U540 ( .A(n459), .ZN(n387) );
  NOR2_X1 U541 ( .A1(n545), .A2(n388), .ZN(n546) );
  NAND2_X1 U542 ( .A1(n389), .A2(n347), .ZN(n629) );
  NAND2_X1 U543 ( .A1(n390), .A2(n347), .ZN(n713) );
  NAND2_X1 U544 ( .A1(n391), .A2(n347), .ZN(n706) );
  NAND2_X1 U545 ( .A1(n392), .A2(n347), .ZN(n636) );
  NAND2_X1 U546 ( .A1(n393), .A2(G478), .ZN(n708) );
  NAND2_X1 U547 ( .A1(n393), .A2(G469), .ZN(n644) );
  XNOR2_X1 U548 ( .A(n399), .B(n397), .ZN(n395) );
  XNOR2_X2 U549 ( .A(n533), .B(n476), .ZN(n400) );
  XNOR2_X1 U550 ( .A(n674), .B(KEYINPUT6), .ZN(n616) );
  NAND2_X1 U551 ( .A1(n623), .A2(n724), .ZN(n403) );
  XNOR2_X1 U552 ( .A(n664), .B(KEYINPUT86), .ZN(n579) );
  XNOR2_X1 U553 ( .A(n445), .B(n444), .ZN(n542) );
  BUF_X1 U554 ( .A(n625), .Z(n404) );
  NOR2_X2 U555 ( .A1(n631), .A2(n714), .ZN(n633) );
  NOR2_X2 U556 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U557 ( .A1(n615), .A2(n424), .ZN(n425) );
  XNOR2_X1 U558 ( .A(n406), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U559 ( .A1(n707), .A2(n714), .ZN(n406) );
  XNOR2_X1 U560 ( .A(n407), .B(n638), .ZN(G57) );
  NOR2_X2 U561 ( .A1(n637), .A2(n714), .ZN(n407) );
  NAND2_X1 U562 ( .A1(n509), .A2(G902), .ZN(n587) );
  NAND2_X1 U563 ( .A1(n606), .A2(n409), .ZN(n607) );
  XNOR2_X2 U564 ( .A(n494), .B(G472), .ZN(n674) );
  NOR2_X1 U565 ( .A1(n651), .A2(n741), .ZN(n606) );
  NAND2_X1 U566 ( .A1(n617), .A2(n414), .ZN(n413) );
  INV_X1 U567 ( .A(KEYINPUT65), .ZN(n416) );
  XNOR2_X2 U568 ( .A(n441), .B(G143), .ZN(n533) );
  XNOR2_X1 U569 ( .A(n498), .B(KEYINPUT16), .ZN(n421) );
  INV_X1 U570 ( .A(n593), .ZN(n422) );
  XNOR2_X2 U571 ( .A(n592), .B(KEYINPUT0), .ZN(n593) );
  NAND2_X1 U572 ( .A1(n607), .A2(KEYINPUT44), .ZN(n423) );
  NOR2_X1 U573 ( .A1(n581), .A2(n434), .ZN(n433) );
  NAND2_X1 U574 ( .A1(n438), .A2(n437), .ZN(n449) );
  INV_X1 U575 ( .A(n688), .ZN(n437) );
  XNOR2_X1 U576 ( .A(n492), .B(n439), .ZN(n493) );
  XNOR2_X2 U577 ( .A(n440), .B(KEYINPUT45), .ZN(n724) );
  XNOR2_X2 U578 ( .A(G128), .B(KEYINPUT80), .ZN(n441) );
  XNOR2_X2 U579 ( .A(n443), .B(n442), .ZN(n740) );
  NAND2_X1 U580 ( .A1(n473), .A2(G221), .ZN(n446) );
  INV_X1 U581 ( .A(n560), .ZN(n574) );
  NAND2_X1 U582 ( .A1(n612), .A2(n497), .ZN(n569) );
  AND2_X1 U583 ( .A1(n512), .A2(n497), .ZN(n450) );
  XNOR2_X1 U584 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U585 ( .A(n522), .B(n521), .Z(n456) );
  NOR2_X1 U586 ( .A1(n602), .A2(n601), .ZN(n457) );
  XOR2_X1 U587 ( .A(n463), .B(n462), .Z(n458) );
  AND2_X1 U588 ( .A1(n606), .A2(n603), .ZN(n604) );
  XNOR2_X1 U589 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U590 ( .A(n490), .B(n489), .ZN(n492) );
  INV_X1 U591 ( .A(n595), .ZN(n596) );
  XNOR2_X1 U592 ( .A(G134), .B(KEYINPUT114), .ZN(n540) );
  NAND2_X1 U593 ( .A1(n732), .A2(G234), .ZN(n461) );
  XNOR2_X1 U594 ( .A(n461), .B(n460), .ZN(n532) );
  NAND2_X1 U595 ( .A1(G221), .A2(n532), .ZN(n464) );
  XNOR2_X1 U596 ( .A(n464), .B(n458), .ZN(n465) );
  XOR2_X1 U597 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n470) );
  INV_X1 U598 ( .A(n625), .ZN(n468) );
  NAND2_X1 U599 ( .A1(G217), .A2(n473), .ZN(n469) );
  XOR2_X1 U600 ( .A(n470), .B(n469), .Z(n471) );
  INV_X1 U601 ( .A(KEYINPUT95), .ZN(n474) );
  XNOR2_X1 U602 ( .A(n675), .B(n474), .ZN(n598) );
  INV_X1 U603 ( .A(n598), .ZN(n475) );
  NAND2_X1 U604 ( .A1(n732), .A2(G227), .ZN(n479) );
  XNOR2_X1 U605 ( .A(n479), .B(G146), .ZN(n480) );
  XNOR2_X1 U606 ( .A(n499), .B(n480), .ZN(n481) );
  OR2_X2 U607 ( .A1(n641), .A2(G902), .ZN(n483) );
  XNOR2_X1 U608 ( .A(KEYINPUT71), .B(G469), .ZN(n482) );
  XNOR2_X2 U609 ( .A(n483), .B(n482), .ZN(n544) );
  INV_X1 U610 ( .A(KEYINPUT96), .ZN(n484) );
  XOR2_X1 U611 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n486) );
  NAND2_X1 U612 ( .A1(n518), .A2(G210), .ZN(n485) );
  XNOR2_X1 U613 ( .A(n486), .B(n485), .ZN(n490) );
  NAND2_X1 U614 ( .A1(n634), .A2(n525), .ZN(n494) );
  NAND2_X1 U615 ( .A1(n525), .A2(n495), .ZN(n503) );
  NAND2_X1 U616 ( .A1(n503), .A2(G214), .ZN(n686) );
  AND2_X1 U617 ( .A1(n674), .A2(n686), .ZN(n496) );
  XNOR2_X1 U618 ( .A(n496), .B(KEYINPUT30), .ZN(n497) );
  XOR2_X1 U619 ( .A(KEYINPUT75), .B(G122), .Z(n498) );
  NAND2_X1 U620 ( .A1(n732), .A2(G224), .ZN(n500) );
  XNOR2_X1 U621 ( .A(n500), .B(KEYINPUT77), .ZN(n502) );
  XNOR2_X1 U622 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n501) );
  NAND2_X1 U623 ( .A1(n503), .A2(G210), .ZN(n505) );
  INV_X1 U624 ( .A(KEYINPUT91), .ZN(n504) );
  XNOR2_X1 U625 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U626 ( .A(KEYINPUT38), .B(n574), .ZN(n511) );
  NAND2_X1 U627 ( .A1(G234), .A2(G237), .ZN(n507) );
  NAND2_X1 U628 ( .A1(G952), .A2(n509), .ZN(n697) );
  NOR2_X1 U629 ( .A1(n697), .A2(G953), .ZN(n589) );
  NOR2_X1 U630 ( .A1(n511), .A2(n573), .ZN(n512) );
  INV_X1 U631 ( .A(n541), .ZN(n539) );
  XNOR2_X1 U632 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U633 ( .A(n515), .B(G122), .Z(n517) );
  XNOR2_X1 U634 ( .A(n517), .B(n516), .ZN(n524) );
  NAND2_X1 U635 ( .A1(G214), .A2(n518), .ZN(n520) );
  XNOR2_X1 U636 ( .A(n520), .B(n519), .ZN(n522) );
  XOR2_X1 U637 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n521) );
  XNOR2_X1 U638 ( .A(n729), .B(n456), .ZN(n523) );
  XNOR2_X1 U639 ( .A(n524), .B(n523), .ZN(n627) );
  NAND2_X1 U640 ( .A1(n627), .A2(n525), .ZN(n527) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(G475), .ZN(n526) );
  XNOR2_X1 U642 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U643 ( .A1(G217), .A2(n532), .ZN(n535) );
  INV_X1 U644 ( .A(n533), .ZN(n534) );
  XNOR2_X1 U645 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U646 ( .A(n537), .B(n536), .ZN(n709) );
  OR2_X1 U647 ( .A1(n709), .A2(G902), .ZN(n538) );
  AND2_X1 U648 ( .A1(n570), .A2(n571), .ZN(n659) );
  INV_X1 U649 ( .A(n659), .ZN(n566) );
  NOR2_X1 U650 ( .A1(n539), .A2(n566), .ZN(n581) );
  XOR2_X1 U651 ( .A(n540), .B(n581), .Z(G36) );
  OR2_X1 U652 ( .A1(n570), .A2(n571), .ZN(n565) );
  XOR2_X1 U653 ( .A(G140), .B(KEYINPUT115), .Z(n547) );
  XOR2_X1 U654 ( .A(n547), .B(n580), .Z(G42) );
  NAND2_X1 U655 ( .A1(n687), .A2(n686), .ZN(n548) );
  INV_X1 U656 ( .A(n571), .ZN(n549) );
  NAND2_X1 U657 ( .A1(n570), .A2(n549), .ZN(n551) );
  INV_X1 U658 ( .A(KEYINPUT105), .ZN(n550) );
  XNOR2_X1 U659 ( .A(n551), .B(n550), .ZN(n688) );
  INV_X1 U660 ( .A(n674), .ZN(n611) );
  NOR2_X1 U661 ( .A1(n552), .A2(n611), .ZN(n553) );
  XNOR2_X1 U662 ( .A(n553), .B(KEYINPUT28), .ZN(n555) );
  NAND2_X1 U663 ( .A1(n555), .A2(n554), .ZN(n564) );
  INV_X1 U664 ( .A(n686), .ZN(n559) );
  XNOR2_X1 U665 ( .A(n620), .B(KEYINPUT89), .ZN(n600) );
  NOR2_X1 U666 ( .A1(n564), .A2(n591), .ZN(n655) );
  AND2_X1 U667 ( .A1(n566), .A2(n565), .ZN(n685) );
  INV_X1 U668 ( .A(n685), .ZN(n567) );
  NAND2_X1 U669 ( .A1(n655), .A2(n567), .ZN(n568) );
  XNOR2_X1 U670 ( .A(n568), .B(KEYINPUT47), .ZN(n577) );
  INV_X1 U671 ( .A(n570), .ZN(n572) );
  NAND2_X1 U672 ( .A1(n572), .A2(n571), .ZN(n595) );
  NOR2_X1 U673 ( .A1(n595), .A2(n573), .ZN(n575) );
  NAND2_X1 U674 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U675 ( .A1(n569), .A2(n576), .ZN(n654) );
  NOR2_X1 U676 ( .A1(n577), .A2(n654), .ZN(n578) );
  INV_X1 U677 ( .A(KEYINPUT84), .ZN(n582) );
  XNOR2_X1 U678 ( .A(n583), .B(n582), .ZN(n623) );
  XNOR2_X1 U679 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n584) );
  XNOR2_X1 U680 ( .A(n585), .B(n584), .ZN(n666) );
  NOR2_X1 U681 ( .A1(G898), .A2(n732), .ZN(n586) );
  XNOR2_X1 U682 ( .A(KEYINPUT93), .B(n586), .ZN(n718) );
  NOR2_X1 U683 ( .A1(n718), .A2(n587), .ZN(n588) );
  NOR2_X1 U684 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U685 ( .A(n740), .B(KEYINPUT67), .ZN(n605) );
  NAND2_X1 U686 ( .A1(n617), .A2(n611), .ZN(n599) );
  INV_X1 U687 ( .A(n619), .ZN(n676) );
  XNOR2_X1 U688 ( .A(KEYINPUT79), .B(n410), .ZN(n602) );
  INV_X1 U689 ( .A(n600), .ZN(n601) );
  INV_X1 U690 ( .A(KEYINPUT44), .ZN(n603) );
  NAND2_X1 U691 ( .A1(n605), .A2(n604), .ZN(n608) );
  NOR2_X1 U692 ( .A1(n660), .A2(n345), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n685), .A2(n613), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n614), .B(KEYINPUT104), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n617), .A2(n410), .ZN(n618) );
  XOR2_X1 U696 ( .A(KEYINPUT87), .B(n618), .Z(n622) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n646) );
  NAND2_X1 U699 ( .A1(n724), .A2(n731), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT119), .B(KEYINPUT59), .Z(n626) );
  XNOR2_X1 U701 ( .A(n629), .B(n628), .ZN(n631) );
  INV_X1 U702 ( .A(G952), .ZN(n630) );
  XNOR2_X1 U703 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n632) );
  XNOR2_X1 U704 ( .A(n633), .B(n632), .ZN(G60) );
  INV_X1 U705 ( .A(KEYINPUT63), .ZN(n638) );
  XOR2_X1 U706 ( .A(KEYINPUT62), .B(n634), .Z(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(G137), .B(KEYINPUT127), .ZN(n640) );
  XOR2_X1 U709 ( .A(n640), .B(n639), .Z(G39) );
  XOR2_X1 U710 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n642) );
  XNOR2_X1 U711 ( .A(n641), .B(n642), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U713 ( .A1(n645), .A2(n714), .ZN(G54) );
  XNOR2_X1 U714 ( .A(G101), .B(n646), .ZN(G3) );
  NAND2_X1 U715 ( .A1(n345), .A2(n396), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n647), .B(G104), .ZN(G6) );
  XOR2_X1 U717 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n649) );
  NAND2_X1 U718 ( .A1(n345), .A2(n659), .ZN(n648) );
  XNOR2_X1 U719 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n344), .B(n650), .ZN(G9) );
  XOR2_X1 U721 ( .A(n651), .B(G110), .Z(G12) );
  XOR2_X1 U722 ( .A(G128), .B(KEYINPUT29), .Z(n653) );
  NAND2_X1 U723 ( .A1(n655), .A2(n659), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(G30) );
  XOR2_X1 U725 ( .A(G143), .B(n654), .Z(G45) );
  NAND2_X1 U726 ( .A1(n655), .A2(n396), .ZN(n656) );
  XNOR2_X1 U727 ( .A(n656), .B(G146), .ZN(G48) );
  XNOR2_X1 U728 ( .A(G113), .B(KEYINPUT112), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n396), .A2(n660), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(G15) );
  XOR2_X1 U731 ( .A(G116), .B(KEYINPUT113), .Z(n662) );
  NAND2_X1 U732 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n662), .B(n661), .ZN(G18) );
  XOR2_X1 U734 ( .A(G125), .B(KEYINPUT37), .Z(n663) );
  XNOR2_X1 U735 ( .A(n664), .B(n663), .ZN(G27) );
  BUF_X1 U736 ( .A(n666), .Z(n667) );
  NOR2_X1 U737 ( .A1(n667), .A2(n668), .ZN(n669) );
  NOR2_X1 U738 ( .A1(n669), .A2(G953), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n700) );
  XOR2_X1 U740 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n696) );
  XNOR2_X1 U741 ( .A(n672), .B(KEYINPUT50), .ZN(n673) );
  NOR2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n679) );
  AND2_X1 U743 ( .A1(n675), .A2(n676), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(KEYINPUT49), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U747 ( .A(n682), .B(KEYINPUT116), .ZN(n683) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT51), .ZN(n684) );
  NOR2_X1 U749 ( .A1(n684), .A2(n668), .ZN(n693) );
  NOR2_X1 U750 ( .A1(n687), .A2(n686), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n352), .A2(n690), .ZN(n691) );
  NOR2_X1 U753 ( .A1(n667), .A2(n691), .ZN(n692) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U755 ( .A(n694), .B(KEYINPUT52), .ZN(n695) );
  XNOR2_X1 U756 ( .A(n696), .B(n695), .ZN(n698) );
  NOR2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U759 ( .A(KEYINPUT53), .B(n701), .ZN(G75) );
  XNOR2_X1 U760 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n702) );
  XOR2_X1 U761 ( .A(n702), .B(KEYINPUT82), .Z(n703) );
  XNOR2_X1 U762 ( .A(n704), .B(n703), .ZN(n705) );
  XNOR2_X1 U763 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U764 ( .A1(n714), .A2(n710), .ZN(G63) );
  XNOR2_X1 U765 ( .A(n713), .B(n712), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n716), .B(KEYINPUT122), .ZN(G66) );
  XNOR2_X1 U767 ( .A(n717), .B(KEYINPUT125), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U769 ( .A(n720), .B(KEYINPUT124), .ZN(n728) );
  XOR2_X1 U770 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n722) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U773 ( .A1(n723), .A2(G898), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n724), .A2(n732), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U776 ( .A(n728), .B(n727), .Z(G69) );
  XNOR2_X1 U777 ( .A(n730), .B(n729), .ZN(n735) );
  XNOR2_X1 U778 ( .A(n731), .B(n735), .ZN(n733) );
  NAND2_X1 U779 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U780 ( .A(n734), .B(KEYINPUT126), .ZN(n739) );
  XOR2_X1 U781 ( .A(G227), .B(n735), .Z(n736) );
  NAND2_X1 U782 ( .A1(n736), .A2(G900), .ZN(n737) );
  NAND2_X1 U783 ( .A1(G953), .A2(n737), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n739), .A2(n738), .ZN(G72) );
  XOR2_X1 U785 ( .A(n740), .B(G122), .Z(G24) );
  XOR2_X1 U786 ( .A(G119), .B(n741), .Z(G21) );
endmodule

