//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n616, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(new_n457), .B(KEYINPUT67), .Z(G261));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n454), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT69), .B1(new_n466), .B2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G137), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT70), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n468), .ZN(new_n482));
  INV_X1    g057(.A(G125), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n479), .A2(new_n486), .ZN(G160));
  NAND3_X1  g062(.A1(new_n469), .A2(G2105), .A3(new_n471), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n473), .A2(G136), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  NAND4_X1  g070(.A1(new_n469), .A2(G138), .A3(new_n470), .A4(new_n471), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n482), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n469), .A2(G126), .A3(G2105), .A4(new_n471), .ZN(new_n503));
  OR3_X1    g078(.A1(new_n470), .A2(KEYINPUT71), .A3(G114), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT71), .B1(new_n470), .B2(G114), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n504), .A2(G2104), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n503), .A2(KEYINPUT72), .A3(new_n507), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n502), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n515), .A2(new_n517), .A3(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n515), .A2(new_n517), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(G62), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  XOR2_X1   g106(.A(new_n531), .B(KEYINPUT74), .Z(new_n532));
  AOI21_X1  g107(.A(new_n514), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n529), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  INV_X1    g110(.A(new_n527), .ZN(new_n536));
  AND2_X1   g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n518), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n537), .A2(new_n542), .ZN(G168));
  AOI22_X1  g118(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n514), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n518), .A2(G52), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT75), .B(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n527), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT76), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n551), .A2(G651), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n536), .A2(G81), .B1(G43), .B2(new_n518), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT77), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n518), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n536), .A2(G91), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n525), .A2(G65), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT78), .Z(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  NAND2_X1  g151(.A1(new_n536), .A2(G87), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n518), .A2(G49), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n525), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n514), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n518), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n527), .B2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n518), .A2(G47), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n527), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n590), .A2(KEYINPUT80), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(KEYINPUT80), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n591), .A2(new_n592), .B1(new_n514), .B2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n527), .A2(KEYINPUT81), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT81), .B1(new_n527), .B2(new_n595), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n525), .A2(G66), .ZN(new_n601));
  INV_X1    g176(.A(G79), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n522), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n596), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G301), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n607), .ZN(G284));
  OAI21_X1  g185(.A(new_n608), .B1(new_n609), .B2(new_n607), .ZN(G321));
  NAND2_X1  g186(.A1(G299), .A2(new_n607), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g189(.A(new_n606), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g196(.A1(new_n477), .A2(new_n481), .A3(new_n468), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n629), .B(new_n630), .C1(G111), .C2(new_n470), .ZN(new_n631));
  INV_X1    g206(.A(G135), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI221_X1 g208(.A(new_n631), .B1(new_n472), .B2(new_n632), .C1(new_n633), .C2(new_n488), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT84), .B(G2096), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n626), .A2(new_n636), .ZN(G156));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT85), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  INV_X1    g226(.A(G14), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n648), .B2(new_n649), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT87), .ZN(G401));
  XNOR2_X1  g230(.A(G2084), .B(G2090), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT88), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n657), .A2(new_n659), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n662), .B2(KEYINPUT17), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n657), .B2(new_n659), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(KEYINPUT17), .A3(new_n658), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2096), .B(G2100), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n670), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(new_n674), .A3(new_n676), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n679), .B(new_n680), .C1(new_n678), .C2(new_n677), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT21), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n684), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  NOR2_X1   g265(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n691));
  INV_X1    g266(.A(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(KEYINPUT93), .B1(new_n692), .B2(G16), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n692), .A2(KEYINPUT93), .A3(G16), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n693), .B(new_n694), .C1(G166), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(G1971), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G16), .B2(G23), .ZN(new_n699));
  OR3_X1    g274(.A1(new_n698), .A2(G16), .A3(G23), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n699), .B(new_n700), .C1(G288), .C2(new_n695), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT33), .B(G1976), .Z(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(G6), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n586), .B2(new_n695), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT32), .B(G1981), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT91), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n705), .B(new_n707), .Z(new_n708));
  NOR3_X1   g283(.A1(new_n697), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT34), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n489), .A2(G119), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n473), .A2(G131), .ZN(new_n714));
  OR2_X1    g289(.A1(G95), .A2(G2105), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n715), .B(G2104), .C1(G107), .C2(new_n470), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n713), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n712), .B1(new_n718), .B2(new_n711), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT35), .B(G1991), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G1986), .ZN(new_n722));
  OR2_X1    g297(.A1(G16), .A2(G24), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G290), .B2(new_n695), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n721), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n722), .B2(new_n724), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n691), .B1(new_n710), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n727), .B(new_n728), .Z(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G35), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G162), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT29), .B(G2090), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT23), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n695), .A2(G20), .ZN(new_n735));
  AOI22_X1  g310(.A1(G299), .A2(G16), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n734), .B2(new_n735), .ZN(new_n737));
  INV_X1    g312(.A(G1956), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT30), .B(G28), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n489), .A2(G129), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n473), .A2(G141), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n477), .A2(G105), .ZN(new_n743));
  NAND3_X1  g318(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT26), .Z(new_n745));
  NAND4_X1  g320(.A1(new_n741), .A2(new_n742), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  MUX2_X1   g321(.A(G32), .B(new_n746), .S(G29), .Z(new_n747));
  XOR2_X1   g322(.A(KEYINPUT27), .B(G1996), .Z(new_n748));
  OAI221_X1 g323(.A(new_n739), .B1(G29), .B2(new_n740), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G5), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G171), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1961), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n747), .A2(new_n748), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n711), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n711), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n695), .A2(G4), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n615), .B2(new_n695), .ZN(new_n760));
  INV_X1    g335(.A(G1348), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n753), .A2(new_n754), .A3(new_n758), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n695), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n695), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT99), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT100), .B(G1966), .Z(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n766), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n476), .A2(G103), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT25), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n481), .A2(new_n468), .A3(G127), .ZN(new_n772));
  NAND2_X1  g347(.A1(G115), .A2(G2104), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n470), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n473), .A2(KEYINPUT96), .A3(G139), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n776));
  INV_X1    g351(.A(G139), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n472), .B2(new_n777), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n771), .B(new_n774), .C1(new_n775), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n711), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n711), .B2(G33), .ZN(new_n781));
  INV_X1    g356(.A(G2072), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G11), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(KEYINPUT31), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n711), .B1(new_n786), .B2(G34), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(G34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G160), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n711), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G2084), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n785), .B(new_n794), .C1(KEYINPUT31), .C2(new_n784), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n711), .A2(G26), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n489), .A2(G128), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n473), .A2(G140), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n797), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n796), .B1(new_n802), .B2(new_n711), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n796), .B(new_n803), .S(KEYINPUT28), .Z(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(G2067), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(G2067), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n805), .B(new_n806), .C1(new_n711), .C2(new_n634), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n763), .A2(new_n769), .A3(new_n795), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n729), .A2(new_n733), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n781), .A2(new_n782), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT97), .ZN(new_n811));
  NOR2_X1   g386(.A1(G16), .A2(G19), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n556), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT95), .B(G1341), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n809), .A2(new_n811), .A3(new_n816), .ZN(G311));
  INV_X1    g392(.A(G311), .ZN(G150));
  AOI22_X1  g393(.A1(new_n536), .A2(G93), .B1(G55), .B2(new_n518), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n514), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G860), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT37), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n615), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT39), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n555), .B(new_n821), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n825), .B(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n823), .B1(new_n829), .B2(G860), .ZN(G145));
  XOR2_X1   g405(.A(G160), .B(KEYINPUT102), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n489), .A2(G130), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n473), .A2(G142), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n470), .A2(G118), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT104), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n623), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n717), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT105), .ZN(new_n840));
  INV_X1    g415(.A(new_n508), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n502), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n779), .A2(KEYINPUT103), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n801), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(new_n746), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n746), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n845), .A2(new_n842), .A3(new_n846), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT105), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n839), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n848), .A2(new_n852), .A3(new_n849), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n831), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n831), .ZN(new_n856));
  INV_X1    g431(.A(new_n849), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(new_n847), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n853), .B(new_n856), .C1(new_n858), .C2(new_n840), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n494), .B(new_n634), .Z(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(G37), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n855), .A2(new_n861), .A3(new_n859), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(new_n867), .ZN(G395));
  NAND2_X1  g443(.A1(new_n821), .A2(new_n607), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n606), .B(G299), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n870), .A2(KEYINPUT41), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(KEYINPUT41), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n618), .B(new_n826), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT107), .Z(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n870), .B2(new_n874), .ZN(new_n877));
  XNOR2_X1  g452(.A(G290), .B(G288), .ZN(new_n878));
  XNOR2_X1  g453(.A(G303), .B(new_n586), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT108), .ZN(new_n881));
  MUX2_X1   g456(.A(new_n880), .B(new_n881), .S(KEYINPUT42), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n877), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n869), .B1(new_n883), .B2(new_n607), .ZN(G295));
  OAI21_X1  g459(.A(new_n869), .B1(new_n883), .B2(new_n607), .ZN(G331));
  INV_X1    g460(.A(new_n881), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n887));
  INV_X1    g462(.A(new_n826), .ZN(new_n888));
  AOI21_X1  g463(.A(G286), .B1(new_n573), .B2(new_n574), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n572), .A2(G168), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n826), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n887), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n891), .A2(new_n887), .ZN(new_n895));
  NOR3_X1   g470(.A1(new_n894), .A2(new_n895), .A3(new_n870), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n873), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n886), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n894), .A2(new_n895), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n881), .B(new_n898), .C1(new_n901), .C2(new_n870), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n902), .A3(new_n864), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT110), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n864), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n873), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n897), .A2(new_n870), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n881), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n903), .A2(new_n913), .A3(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n905), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  MUX2_X1   g490(.A(new_n903), .B(new_n910), .S(KEYINPUT43), .Z(new_n916));
  MUX2_X1   g491(.A(new_n915), .B(new_n916), .S(KEYINPUT44), .Z(G397));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n842), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n474), .A2(G40), .A3(new_n485), .A4(new_n478), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n801), .B(G2067), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n746), .B(G1996), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT112), .ZN(new_n929));
  XOR2_X1   g504(.A(new_n717), .B(new_n720), .Z(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n932), .A2(G1986), .A3(G290), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n933), .B(KEYINPUT48), .Z(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n718), .A2(new_n720), .ZN(new_n936));
  OAI22_X1  g511(.A1(new_n929), .A2(new_n936), .B1(G2067), .B2(new_n801), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n925), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n932), .B2(G1996), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n925), .B1(new_n746), .B2(new_n926), .ZN(new_n941));
  INV_X1    g516(.A(G1996), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n925), .A2(KEYINPUT46), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT47), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n935), .A2(new_n938), .A3(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT127), .Z(new_n947));
  AOI21_X1  g522(.A(new_n924), .B1(new_n919), .B2(new_n922), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n512), .A2(new_n918), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(new_n922), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n768), .ZN(new_n951));
  INV_X1    g526(.A(new_n924), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n842), .A2(new_n953), .A3(new_n918), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n503), .A2(KEYINPUT72), .A3(new_n507), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT72), .B1(new_n503), .B2(new_n507), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(G1384), .B1(new_n957), .B2(new_n502), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n952), .B(new_n954), .C1(new_n958), .C2(new_n953), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n951), .B1(G2084), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(G8), .B1(new_n960), .B2(G286), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT51), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT62), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n960), .B2(G286), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n962), .B(new_n963), .C1(new_n961), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n842), .A2(new_n967), .A3(KEYINPUT45), .A4(new_n918), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n496), .A2(KEYINPUT4), .B1(new_n500), .B2(new_n498), .ZN(new_n969));
  OAI211_X1 g544(.A(KEYINPUT45), .B(new_n918), .C1(new_n969), .C2(new_n508), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT113), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n924), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n949), .A2(new_n922), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT53), .B1(new_n974), .B2(new_n757), .ZN(new_n975));
  INV_X1    g550(.A(G1961), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(new_n959), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n757), .A2(KEYINPUT53), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n948), .B(new_n978), .C1(new_n922), .C2(new_n949), .ZN(new_n979));
  AOI21_X1  g554(.A(G301), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n966), .A2(new_n980), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n974), .A2(G1971), .B1(G2090), .B2(new_n959), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  NAND2_X1  g560(.A1(G303), .A2(G8), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT55), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n987), .B(KEYINPUT115), .Z(new_n988));
  NAND4_X1  g563(.A1(new_n984), .A2(G8), .A3(new_n985), .A4(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n586), .B(G1981), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT49), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n919), .A2(new_n924), .ZN(new_n992));
  INV_X1    g567(.A(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G1976), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n996), .B2(G288), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n997), .A2(KEYINPUT52), .ZN(new_n998));
  INV_X1    g573(.A(G288), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G1976), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n997), .A2(KEYINPUT52), .A3(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n995), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n974), .A2(G1971), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n512), .A2(new_n953), .A3(new_n918), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n924), .B1(new_n919), .B2(KEYINPUT50), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n512), .A2(KEYINPUT117), .A3(new_n953), .A4(new_n918), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1009), .A2(G2090), .ZN(new_n1010));
  OAI21_X1  g585(.A(G8), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n987), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n989), .A2(new_n1002), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT126), .B1(new_n981), .B2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n989), .A2(new_n1002), .A3(new_n1012), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT126), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(new_n966), .A4(new_n980), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n962), .B1(new_n961), .B2(new_n965), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(KEYINPUT62), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1014), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n960), .A2(G8), .A3(G168), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(KEYINPUT63), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1012), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n989), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1002), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n999), .A2(new_n996), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT116), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n991), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G305), .A2(G1981), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n994), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT63), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n984), .A2(G8), .A3(new_n985), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1021), .B1(new_n1033), .B2(new_n987), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1034), .B2(new_n1002), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1020), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n1038));
  XNOR2_X1  g613(.A(G299), .B(KEYINPUT57), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1009), .A2(new_n738), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n972), .A2(new_n973), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1040), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1041), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n606), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n924), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1348), .B1(new_n1047), .B2(new_n954), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n919), .A2(G2067), .A3(new_n924), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT118), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n959), .A2(new_n761), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1049), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1044), .B1(new_n1046), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT61), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1045), .A2(new_n1044), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n606), .B1(new_n1055), .B2(KEYINPUT60), .ZN(new_n1063));
  AOI211_X1 g638(.A(new_n1061), .B(new_n615), .C1(new_n1050), .C2(new_n1054), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1039), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1041), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT61), .B1(new_n1044), .B2(KEYINPUT121), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1060), .B(new_n1065), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n968), .A2(new_n971), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1076), .A2(new_n973), .A3(new_n942), .A4(new_n952), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT119), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n972), .A2(new_n1079), .A3(new_n942), .A4(new_n973), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g656(.A(KEYINPUT58), .B(G1341), .Z(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n919), .B2(new_n924), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT120), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1081), .A2(new_n1086), .A3(new_n1083), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n556), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1085), .A2(KEYINPUT59), .A3(new_n556), .A4(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1038), .B(new_n1057), .C1(new_n1075), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1045), .A2(new_n1044), .A3(KEYINPUT121), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1066), .A2(KEYINPUT121), .A3(new_n1039), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1058), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT122), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1070), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1052), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1101));
  AOI211_X1 g676(.A(KEYINPUT118), .B(new_n1049), .C1(new_n959), .C2(new_n761), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n615), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1059), .B1(new_n1106), .B2(new_n1062), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1100), .A2(new_n1107), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1038), .B1(new_n1108), .B2(new_n1057), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1094), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n923), .A2(new_n478), .A3(new_n474), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n1112));
  OAI21_X1  g687(.A(G2105), .B1(new_n484), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1112), .B2(new_n484), .ZN(new_n1114));
  INV_X1    g689(.A(G40), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1076), .A2(new_n978), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n977), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G171), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n977), .A2(G301), .A3(new_n979), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(KEYINPUT54), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1121), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1122));
  INV_X1    g697(.A(new_n980), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n609), .B2(new_n1118), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(KEYINPUT125), .A3(new_n1125), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1122), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1037), .B1(new_n1110), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(G290), .B(new_n722), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n931), .B1(new_n932), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n947), .B1(new_n1131), .B2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g709(.A(new_n464), .ZN(new_n1136));
  NOR3_X1   g710(.A1(G401), .A2(new_n1136), .A3(G227), .ZN(new_n1137));
  NAND4_X1  g711(.A1(new_n915), .A2(new_n1137), .A3(new_n689), .A4(new_n866), .ZN(G225));
  INV_X1    g712(.A(G225), .ZN(G308));
endmodule


