//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n613, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n468), .B2(G125), .ZN(new_n469));
  OAI211_X1 g044(.A(KEYINPUT68), .B(G125), .C1(new_n462), .C2(new_n463), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n467), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n466), .B1(new_n472), .B2(G2105), .ZN(G160));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n475));
  INV_X1    g050(.A(G136), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G124), .ZN(new_n478));
  OAI221_X1 g053(.A(new_n475), .B1(new_n464), .B2(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g058(.A(G138), .B1(new_n481), .B2(KEYINPUT69), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n464), .B2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n486), .B1(new_n487), .B2(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n468), .A2(new_n488), .A3(new_n459), .A4(new_n482), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n459), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n485), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  XNOR2_X1  g069(.A(KEYINPUT5), .B(G543), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n495), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OAI21_X1  g080(.A(G543), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n498), .A2(new_n507), .ZN(G303));
  INV_X1    g083(.A(G303), .ZN(G166));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n499), .A2(G89), .ZN(new_n513));
  NAND2_X1  g088(.A1(G63), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT7), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT7), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n518), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n506), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT70), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  OR2_X1    g099(.A1(KEYINPUT6), .A2(G651), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(new_n503), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n526), .A2(G51), .B1(new_n517), .B2(new_n519), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n499), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n527), .B(new_n528), .C1(new_n512), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(new_n530), .ZN(G168));
  INV_X1    g106(.A(KEYINPUT72), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n526), .A2(G52), .ZN(new_n533));
  XNOR2_X1  g108(.A(KEYINPUT71), .B(G90), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n495), .A2(new_n499), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g111(.A(G64), .B1(new_n510), .B2(new_n511), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n497), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n532), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n537), .A2(new_n538), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G651), .ZN(new_n542));
  NAND4_X1  g117(.A1(new_n542), .A2(KEYINPUT72), .A3(new_n533), .A4(new_n535), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n500), .A2(new_n545), .B1(new_n546), .B2(new_n506), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n495), .A2(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n497), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND2_X1  g131(.A1(new_n526), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n495), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT73), .Z(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n495), .A2(new_n499), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G91), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n558), .A2(new_n562), .A3(new_n564), .ZN(G299));
  AND3_X1   g140(.A1(new_n540), .A2(KEYINPUT74), .A3(new_n543), .ZN(new_n566));
  AOI21_X1  g141(.A(KEYINPUT74), .B1(new_n540), .B2(new_n543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  OAI21_X1  g144(.A(G651), .B1(new_n495), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n495), .A2(new_n499), .A3(G87), .ZN(new_n571));
  OAI211_X1 g146(.A(G49), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  OAI21_X1  g148(.A(G61), .B1(new_n510), .B2(new_n511), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(G48), .B2(new_n526), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n495), .A2(new_n499), .A3(G86), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n495), .A2(new_n499), .A3(KEYINPUT75), .A4(G86), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n495), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n497), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT76), .B(G85), .ZN(new_n585));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n500), .A2(new_n585), .B1(new_n586), .B2(new_n506), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n563), .A2(new_n590), .A3(G92), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT77), .B1(new_n500), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n526), .A2(G54), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT78), .B(G66), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n495), .A2(new_n598), .B1(G79), .B2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n599), .B2(new_n497), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n591), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n596), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT74), .ZN(new_n605));
  NAND2_X1  g180(.A1(G171), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n540), .A2(KEYINPUT74), .A3(new_n543), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(G868), .B2(new_n608), .ZN(G284));
  AOI21_X1  g184(.A(new_n604), .B1(G868), .B2(new_n608), .ZN(G321));
  MUX2_X1   g185(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g186(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g187(.A(G860), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n603), .B1(G559), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(KEYINPUT79), .Z(G148));
  OR2_X1    g190(.A1(new_n603), .A2(G559), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n468), .A2(new_n460), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n628));
  INV_X1    g203(.A(G135), .ZN(new_n629));
  INV_X1    g204(.A(G123), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n628), .B1(new_n464), .B2(new_n629), .C1(new_n477), .C2(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G2096), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n625), .A2(new_n626), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2427), .B(G2430), .Z(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT82), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(G401));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT83), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n632), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AOI211_X1 g250(.A(new_n672), .B(new_n675), .C1(new_n667), .C2(new_n671), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT86), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1981), .B(G1986), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT85), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(G229));
  INV_X1    g259(.A(G29), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G32), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n460), .A2(G105), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(KEYINPUT96), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(KEYINPUT96), .ZN(new_n689));
  INV_X1    g264(.A(new_n477), .ZN(new_n690));
  AOI22_X1  g265(.A1(new_n688), .A2(new_n689), .B1(G129), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT26), .Z(new_n693));
  AND2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n464), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G141), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT95), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n686), .B1(new_n699), .B2(new_n685), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT27), .B(G1996), .Z(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT97), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT24), .ZN(new_n704));
  INV_X1    g279(.A(G34), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G160), .B2(new_n685), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n703), .B1(G2084), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n685), .A2(G35), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G162), .B2(new_n685), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT29), .Z(new_n712));
  INV_X1    g287(.A(G2090), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G2072), .ZN(new_n715));
  OR2_X1    g290(.A1(G29), .A2(G33), .ZN(new_n716));
  NAND2_X1  g291(.A1(G115), .A2(G2104), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n462), .A2(new_n463), .ZN(new_n718));
  INV_X1    g293(.A(G127), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n459), .B1(new_n720), .B2(KEYINPUT94), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT94), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n695), .A2(G139), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT25), .Z(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n716), .B1(new_n726), .B2(new_n685), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n709), .B(new_n714), .C1(new_n715), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G5), .A2(G16), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(G171), .B2(G16), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G27), .A2(G29), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G164), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT100), .ZN(new_n735));
  INV_X1    g310(.A(new_n603), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G4), .B2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT93), .B(G1348), .Z(new_n740));
  OAI221_X1 g315(.A(new_n732), .B1(new_n735), .B2(G2078), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n737), .A2(G20), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G299), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n737), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n746), .A2(G1956), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(G1956), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n685), .A2(G26), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n690), .A2(G128), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n695), .A2(G140), .ZN(new_n752));
  OR2_X1    g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(new_n685), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n747), .A2(new_n748), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(G28), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n685), .B1(new_n760), .B2(G28), .ZN(new_n762));
  AND2_X1   g337(.A1(KEYINPUT31), .A2(G11), .ZN(new_n763));
  NOR2_X1   g338(.A1(KEYINPUT31), .A2(G11), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n631), .A2(new_n685), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT99), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n551), .B2(G16), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1341), .ZN(new_n772));
  NAND2_X1  g347(.A1(G286), .A2(G16), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n737), .A2(G21), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT98), .B(G1966), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AOI211_X1 g352(.A(new_n769), .B(new_n772), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n739), .A2(new_n740), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n735), .A2(G2078), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n759), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n775), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n782), .A2(new_n776), .B1(new_n715), .B2(new_n727), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n783), .B1(G2084), .B2(new_n708), .C1(new_n713), .C2(new_n712), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n728), .A2(new_n741), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(G95), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n788));
  INV_X1    g363(.A(G131), .ZN(new_n789));
  INV_X1    g364(.A(G119), .ZN(new_n790));
  OAI221_X1 g365(.A(new_n788), .B1(new_n464), .B2(new_n789), .C1(new_n477), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT87), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT88), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  MUX2_X1   g369(.A(G25), .B(new_n794), .S(G29), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT35), .B(G1991), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G24), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n588), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT90), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1986), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n799), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n737), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n737), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1971), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT32), .B(G1981), .ZN(new_n809));
  MUX2_X1   g384(.A(G6), .B(G305), .S(G16), .Z(new_n810));
  AOI21_X1  g385(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n809), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G23), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT91), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n510), .A2(new_n511), .A3(G74), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n572), .B1(new_n815), .B2(new_n497), .ZN(new_n816));
  AND3_X1   g391(.A1(new_n495), .A2(new_n499), .A3(G87), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT91), .A4(new_n572), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n813), .B1(new_n820), .B2(G16), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT33), .B(G1976), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n812), .A2(KEYINPUT92), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT92), .B1(new_n812), .B2(new_n823), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(KEYINPUT34), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT34), .ZN(new_n828));
  INV_X1    g403(.A(new_n826), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n824), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n805), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n805), .A2(new_n833), .A3(new_n827), .A4(new_n830), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n786), .B1(new_n832), .B2(new_n834), .ZN(G311));
  INV_X1    g410(.A(G311), .ZN(G150));
  NAND2_X1  g411(.A1(new_n736), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n495), .A2(new_n499), .A3(G93), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT102), .B(G55), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n506), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n495), .A2(G67), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n497), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT103), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G67), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n843), .B1(new_n512), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G651), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n506), .A2(new_n840), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .A4(new_n839), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n526), .A2(G43), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n495), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n853));
  OAI221_X1 g428(.A(new_n852), .B1(new_n500), .B2(new_n545), .C1(new_n853), .C2(new_n497), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n845), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n848), .A2(new_n839), .A3(new_n849), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n551), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n845), .A2(new_n851), .A3(new_n854), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n838), .B(new_n861), .Z(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n613), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n845), .A2(new_n851), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G860), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT37), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n865), .A2(new_n868), .ZN(G145));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n726), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n698), .B(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n695), .A2(G142), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT106), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n690), .A2(G130), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n459), .A2(G118), .ZN(new_n876));
  OAI21_X1  g451(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n872), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G164), .B(new_n755), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n882), .A3(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n792), .B(new_n622), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n884), .A2(new_n887), .A3(new_n885), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G160), .B(new_n631), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G162), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n890), .A3(new_n896), .A4(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g475(.A(G868), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n866), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n616), .B(new_n861), .Z(new_n903));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n600), .B1(new_n594), .B2(new_n595), .ZN(new_n905));
  NAND3_X1  g480(.A1(G299), .A2(new_n905), .A3(new_n602), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G299), .B1(new_n905), .B2(new_n602), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n903), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n745), .A2(new_n603), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n906), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n911), .B2(KEYINPUT41), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n913), .B1(new_n903), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT42), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(KEYINPUT109), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n919), .B(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n820), .B(G305), .ZN(new_n923));
  XNOR2_X1  g498(.A(G303), .B(new_n588), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(KEYINPUT109), .B2(new_n920), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n922), .B(new_n927), .Z(new_n928));
  OAI21_X1  g503(.A(new_n902), .B1(new_n928), .B2(new_n901), .ZN(G295));
  OAI21_X1  g504(.A(new_n902), .B1(new_n928), .B2(new_n901), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  AOI21_X1  g506(.A(G168), .B1(new_n543), .B2(new_n540), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n932), .B1(G301), .B2(G168), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n861), .A2(KEYINPUT110), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n859), .A2(new_n935), .A3(new_n860), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(G286), .A2(G171), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n608), .B2(G286), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n859), .A2(new_n935), .A3(new_n860), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n935), .B1(new_n859), .B2(new_n860), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n912), .B1(new_n943), .B2(new_n915), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n937), .A2(new_n942), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n945), .B(KEYINPUT41), .C1(new_n907), .C2(new_n908), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n926), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n911), .A2(new_n937), .A3(new_n942), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT108), .B1(new_n914), .B2(new_n906), .ZN(new_n949));
  INV_X1    g524(.A(new_n910), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT41), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n916), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n925), .B(new_n948), .C1(new_n943), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n898), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n931), .B1(new_n954), .B2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n898), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n918), .A2(new_n945), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n925), .B1(new_n957), .B2(new_n948), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(KEYINPUT43), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT43), .B1(new_n956), .B2(new_n958), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n956), .C2(new_n958), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n947), .A2(new_n965), .A3(new_n898), .A4(new_n953), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n967), .A2(KEYINPUT112), .A3(new_n931), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT112), .B1(new_n967), .B2(new_n931), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n960), .B1(new_n968), .B2(new_n969), .ZN(G397));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n493), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n466), .ZN(new_n975));
  INV_X1    g550(.A(new_n467), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT68), .ZN(new_n977));
  INV_X1    g552(.A(G125), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n977), .B1(new_n718), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n979), .B2(new_n470), .ZN(new_n980));
  OAI211_X1 g555(.A(G40), .B(new_n975), .C1(new_n980), .C2(new_n459), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n755), .B(G2067), .Z(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n699), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n985), .B2(new_n699), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n792), .B(new_n796), .Z(new_n988));
  AOI21_X1  g563(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(KEYINPUT127), .ZN(new_n992));
  NOR2_X1   g567(.A1(G290), .A2(G1986), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n982), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT48), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n699), .B1(new_n997), .B2(G1996), .ZN(new_n998));
  INV_X1    g573(.A(new_n984), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n982), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n982), .A2(new_n985), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT126), .B1(new_n1001), .B2(new_n997), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n1001), .A2(KEYINPUT126), .A3(new_n997), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n987), .A2(new_n983), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n1006), .A2(new_n796), .A3(new_n794), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n755), .A2(G2067), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n982), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n996), .A2(new_n1005), .A3(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(G160), .A2(G40), .A3(new_n971), .A4(new_n493), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT115), .B(G1981), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n577), .A2(new_n580), .A3(new_n581), .A4(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n526), .A2(G48), .ZN(new_n1014));
  INV_X1    g589(.A(new_n575), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n495), .B2(G61), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1014), .B(new_n578), .C1(new_n1016), .C2(new_n497), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G1981), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1013), .A2(new_n1018), .A3(KEYINPUT49), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1021), .A2(G8), .A3(new_n1011), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G288), .A2(G1976), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1013), .ZN(new_n1026));
  OAI211_X1 g601(.A(G8), .B(new_n1011), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n981), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n972), .A2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n493), .A2(new_n1034), .A3(new_n971), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n713), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n973), .A2(G1384), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n972), .A2(new_n973), .B1(new_n493), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1971), .B1(new_n1038), .B2(new_n1032), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1036), .B1(new_n1039), .B2(KEYINPUT113), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n493), .A2(new_n1037), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT45), .B1(new_n493), .B2(new_n971), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1042), .A2(new_n1043), .A3(new_n981), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1044), .A2(new_n1045), .A3(G1971), .ZN(new_n1046));
  OAI211_X1 g621(.A(G8), .B(new_n1031), .C1(new_n1040), .C2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n818), .A2(G1976), .A3(new_n819), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(G8), .C1(new_n981), .C2(new_n972), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT52), .ZN(new_n1050));
  INV_X1    g625(.A(G1976), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT52), .B1(G288), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1011), .A2(G8), .A3(new_n1048), .A4(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1023), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1027), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G2084), .ZN(new_n1056));
  AND4_X1   g631(.A1(new_n1056), .A2(new_n1032), .A3(new_n1033), .A4(new_n1035), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1966), .B1(new_n1038), .B2(new_n1032), .ZN(new_n1058));
  OAI211_X1 g633(.A(G8), .B(G168), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1023), .A2(KEYINPUT63), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1047), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1045), .B1(new_n1044), .B2(G1971), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1039), .A2(KEYINPUT113), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n1036), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1031), .B1(new_n1065), .B2(G8), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT117), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(G8), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1030), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1047), .A4(new_n1061), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1054), .A2(KEYINPUT116), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1023), .A2(new_n1075), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1036), .B1(new_n1044), .B2(G1971), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(G8), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n1030), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1047), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1073), .B1(new_n1081), .B2(new_n1059), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1055), .B1(new_n1072), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1032), .A2(new_n974), .A3(new_n1041), .ZN(new_n1086));
  INV_X1    g661(.A(G1966), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1032), .A2(new_n1033), .A3(new_n1056), .A4(new_n1035), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1085), .B(G8), .C1(new_n1090), .C2(G286), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1092));
  NAND2_X1  g667(.A1(G286), .A2(G8), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(KEYINPUT51), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1093), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1090), .B2(new_n1096), .ZN(new_n1097));
  AOI211_X1 g672(.A(KEYINPUT122), .B(new_n1093), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1091), .B(new_n1094), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(G2078), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1044), .A2(new_n1102), .B1(new_n1103), .B2(new_n731), .ZN(new_n1104));
  INV_X1    g679(.A(G2078), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1032), .A2(new_n974), .A3(new_n1105), .A4(new_n1041), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1101), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n731), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n980), .A2(KEYINPUT123), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n980), .A2(KEYINPUT123), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(G2105), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n975), .A2(G40), .A3(new_n1102), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n974), .A3(new_n1041), .A4(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1107), .A2(new_n1109), .A3(G301), .A4(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1100), .B1(new_n1108), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1107), .A2(new_n1109), .A3(new_n1114), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1100), .B1(new_n1118), .B2(G171), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1104), .A2(G301), .A3(new_n1107), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1099), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT124), .B1(new_n1122), .B2(new_n1081), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1038), .A2(new_n1032), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1956), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1103), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1038), .A2(KEYINPUT118), .A3(new_n1032), .A4(new_n1125), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G299), .B(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1128), .A2(new_n1134), .A3(new_n1130), .A4(new_n1131), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1124), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n981), .A2(new_n972), .A3(G2067), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1103), .A2(new_n740), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT119), .B1(new_n1011), .B2(G2067), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n603), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n736), .A2(KEYINPUT60), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1142), .A2(KEYINPUT60), .A3(new_n736), .A4(new_n1143), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1150), .A2(KEYINPUT121), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT58), .B(G1341), .Z(new_n1152));
  AOI22_X1  g727(.A1(new_n1044), .A2(new_n985), .B1(new_n1011), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1153), .B2(new_n854), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1011), .A2(new_n1152), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1086), .B2(G1996), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(new_n551), .C1(KEYINPUT121), .C2(new_n1150), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1148), .A2(new_n1149), .B1(new_n1154), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1134), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n745), .A2(new_n1133), .ZN(new_n1161));
  NOR2_X1   g736(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1162));
  OAI21_X1  g737(.A(KEYINPUT120), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1132), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1139), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n603), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1132), .A2(new_n1164), .B1(new_n1168), .B2(new_n1137), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1102), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1109), .B1(new_n1086), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1107), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n608), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1115), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1175), .A2(new_n1100), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1077), .A2(new_n1047), .A3(new_n1080), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1099), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1123), .A2(new_n1170), .A3(new_n1179), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1083), .A2(new_n1084), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1084), .B1(new_n1083), .B2(new_n1180), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1108), .B1(new_n1099), .B2(KEYINPUT62), .ZN(new_n1183));
  AOI211_X1 g758(.A(new_n1081), .B(new_n1183), .C1(KEYINPUT62), .C2(new_n1099), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  AND2_X1   g760(.A1(G290), .A2(G1986), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n982), .B1(new_n1186), .B2(new_n993), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n990), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1010), .B1(new_n1185), .B2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g764(.A(G319), .ZN(new_n1191));
  NOR3_X1   g765(.A1(G229), .A2(new_n1191), .A3(G227), .ZN(new_n1192));
  NAND4_X1  g766(.A1(new_n899), .A2(new_n967), .A3(new_n651), .A4(new_n1192), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


