//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT87), .Z(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  XOR2_X1   g011(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(G101), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT79), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n197), .A2(new_n198), .A3(new_n201), .A4(G101), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n204));
  XNOR2_X1  g018(.A(G116), .B(G119), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT2), .B(G113), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n205), .B(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G101), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n192), .A2(new_n195), .A3(new_n209), .A4(new_n196), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n210), .A2(KEYINPUT4), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n197), .A2(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n203), .A2(new_n204), .A3(new_n208), .A4(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n215), .A2(G116), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n215), .A2(G116), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n206), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n205), .A2(KEYINPUT5), .ZN(new_n219));
  INV_X1    g033(.A(G113), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT5), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n218), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n191), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n194), .A2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n210), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n214), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n200), .A2(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n204), .B1(new_n231), .B2(new_n208), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n190), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n203), .A2(new_n208), .A3(new_n213), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT80), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n235), .A2(new_n189), .A3(new_n214), .A4(new_n229), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(KEYINPUT6), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G224), .ZN(new_n238));
  OR3_X1    g052(.A1(new_n238), .A2(KEYINPUT82), .A3(G953), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT82), .B1(new_n238), .B2(G953), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT81), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT83), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  OAI21_X1  g060(.A(G128), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n244), .A2(KEYINPUT65), .A3(G146), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT65), .B1(new_n244), .B2(G146), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n249), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n248), .B2(G143), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n244), .A2(KEYINPUT65), .A3(G146), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n245), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n254), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n252), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G125), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT0), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(new_n253), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n249), .A2(new_n250), .B1(KEYINPUT0), .B2(G128), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n253), .A3(KEYINPUT64), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(KEYINPUT0), .B2(G128), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n263), .A2(new_n269), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n275), .A2(new_n266), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n243), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n190), .C1(new_n230), .C2(new_n232), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n237), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n241), .ZN(new_n282));
  AND4_X1   g096(.A1(KEYINPUT7), .A2(new_n267), .A3(new_n276), .A4(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT85), .B(KEYINPUT7), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n267), .A2(new_n276), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n227), .A2(KEYINPUT84), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n286), .A2(new_n223), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n189), .B(KEYINPUT8), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(new_n286), .B2(new_n223), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n283), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n291), .B2(new_n236), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n281), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n188), .B1(new_n293), .B2(KEYINPUT86), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT86), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n281), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n281), .A2(new_n292), .A3(new_n187), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G214), .B1(G237), .B2(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G113), .B(G122), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(new_n191), .ZN(new_n303));
  INV_X1    g117(.A(G237), .ZN(new_n304));
  INV_X1    g118(.A(G953), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G214), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n244), .ZN(new_n307));
  INV_X1    g121(.A(G131), .ZN(new_n308));
  NOR2_X1   g122(.A1(G237), .A2(G953), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT89), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n307), .A2(new_n313), .A3(new_n308), .A4(new_n310), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n309), .A2(G143), .A3(G214), .ZN(new_n315));
  AOI21_X1  g129(.A(G143), .B1(new_n309), .B2(G214), .ZN(new_n316));
  OAI21_X1  g130(.A(G131), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n266), .A2(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n266), .A2(G140), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT16), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n325), .A3(G146), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT19), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n319), .A2(G125), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n320), .A2(new_n321), .A3(KEYINPUT19), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n248), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n318), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n320), .A2(new_n321), .A3(new_n248), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n248), .B1(new_n320), .B2(new_n321), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G146), .B1(new_n323), .B2(new_n328), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n320), .A2(new_n321), .A3(new_n248), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(KEYINPUT88), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(KEYINPUT18), .A2(G131), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n315), .B2(new_n316), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n307), .A2(KEYINPUT18), .A3(G131), .A4(new_n310), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n337), .A2(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n303), .B1(new_n333), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n322), .A2(new_n325), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n248), .ZN(new_n348));
  OAI211_X1 g162(.A(KEYINPUT17), .B(G131), .C1(new_n315), .C2(new_n316), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n348), .A2(new_n349), .A3(new_n326), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT17), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n312), .A2(new_n351), .A3(new_n314), .A4(new_n317), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(new_n303), .A3(new_n345), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n344), .B1(new_n350), .B2(new_n352), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT90), .A3(new_n303), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n346), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(G475), .A2(G902), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT92), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n346), .ZN(new_n364));
  AND4_X1   g178(.A1(KEYINPUT90), .A2(new_n353), .A3(new_n303), .A4(new_n345), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT90), .B1(new_n357), .B2(new_n303), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n368));
  INV_X1    g182(.A(new_n362), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n356), .A2(new_n358), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT91), .A3(new_n364), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n360), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(KEYINPUT20), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G475), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n374), .B1(new_n303), .B2(new_n357), .ZN(new_n379));
  INV_X1    g193(.A(G902), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT93), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n383));
  INV_X1    g197(.A(new_n381), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT91), .B1(new_n374), .B2(new_n364), .ZN(new_n385));
  AOI211_X1 g199(.A(new_n372), .B(new_n346), .C1(new_n356), .C2(new_n358), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n361), .B1(new_n387), .B2(new_n360), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n383), .B(new_n384), .C1(new_n388), .C2(new_n371), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT9), .B(G234), .ZN(new_n391));
  OAI21_X1  g205(.A(G221), .B1(new_n391), .B2(G902), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT77), .ZN(new_n393));
  INV_X1    g207(.A(G469), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n380), .ZN(new_n395));
  INV_X1    g209(.A(new_n265), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT10), .A3(new_n228), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n231), .A2(new_n275), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT10), .ZN(new_n399));
  INV_X1    g213(.A(new_n263), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n259), .A2(new_n264), .B1(new_n400), .B2(new_n247), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n399), .B1(new_n401), .B2(new_n227), .ZN(new_n402));
  INV_X1    g216(.A(G137), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n403), .A2(KEYINPUT11), .A3(G134), .ZN(new_n404));
  INV_X1    g218(.A(G134), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G137), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(G137), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n404), .B(new_n406), .C1(new_n407), .C2(KEYINPUT11), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT66), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(G131), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT11), .B1(new_n403), .B2(G134), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n403), .A2(G134), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n409), .A2(G131), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n404), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n397), .A2(new_n398), .A3(new_n402), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n265), .A2(new_n227), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n227), .B2(new_n401), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n420), .A2(KEYINPUT12), .A3(new_n416), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT12), .B1(new_n420), .B2(new_n416), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n305), .A2(G227), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n397), .A2(new_n398), .A3(new_n402), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n416), .ZN(new_n428));
  INV_X1    g242(.A(new_n426), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n423), .A2(new_n426), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n395), .B1(new_n431), .B2(G469), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n421), .A2(new_n422), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n418), .A2(new_n429), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n429), .B1(new_n428), .B2(new_n418), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n394), .B(new_n380), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n393), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n244), .A2(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n253), .A2(G143), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G134), .ZN(new_n443));
  XNOR2_X1  g257(.A(G128), .B(G143), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n405), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT94), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT94), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G116), .B(G122), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT14), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G122), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G116), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n194), .B1(new_n454), .B2(KEYINPUT14), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n452), .A2(new_n455), .B1(new_n194), .B2(new_n450), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n447), .A2(new_n449), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(G134), .C1(KEYINPUT13), .C2(new_n440), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n450), .B(new_n194), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n445), .ZN(new_n461));
  INV_X1    g275(.A(G217), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n391), .A2(new_n462), .A3(G953), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n457), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n463), .B1(new_n457), .B2(new_n461), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n380), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G478), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(KEYINPUT15), .ZN(new_n470));
  OAI211_X1 g284(.A(KEYINPUT95), .B(new_n380), .C1(new_n464), .C2(new_n465), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n466), .A2(new_n470), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G952), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n476), .A2(KEYINPUT96), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(KEYINPUT96), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n305), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(G234), .B2(G237), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT21), .B(G898), .ZN(new_n482));
  NAND2_X1  g296(.A1(G234), .A2(G237), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(G902), .A3(G953), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  NOR4_X1   g300(.A1(new_n301), .A2(new_n390), .A3(new_n439), .A4(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n416), .A2(new_n275), .ZN(new_n489));
  AOI21_X1  g303(.A(G131), .B1(new_n413), .B2(new_n404), .ZN(new_n490));
  NOR3_X1   g304(.A1(new_n407), .A2(new_n412), .A3(new_n308), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n489), .B1(new_n265), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n208), .ZN(new_n494));
  OAI21_X1  g308(.A(KEYINPUT68), .B1(new_n490), .B2(new_n491), .ZN(new_n495));
  INV_X1    g309(.A(new_n491), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n408), .A2(new_n308), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT68), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n207), .B(new_n489), .C1(new_n500), .C2(new_n265), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT70), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n503), .B1(new_n494), .B2(new_n501), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n501), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n309), .A2(G210), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n513), .B(KEYINPUT27), .Z(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n493), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT30), .B(new_n489), .C1(new_n500), .C2(new_n265), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n208), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n501), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n517), .B1(new_n522), .B2(new_n516), .ZN(new_n523));
  INV_X1    g337(.A(new_n516), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n521), .A2(KEYINPUT31), .A3(new_n524), .A4(new_n501), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n512), .A2(new_n516), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(G472), .A2(G902), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n488), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n511), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n489), .B1(new_n500), .B2(new_n265), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n208), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n501), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n530), .B1(new_n533), .B2(KEYINPUT28), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n516), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n511), .B1(new_n508), .B2(KEYINPUT70), .ZN(new_n538));
  AOI211_X1 g352(.A(new_n506), .B(new_n503), .C1(new_n494), .C2(new_n501), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n538), .A2(new_n516), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n522), .A2(new_n516), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n535), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n537), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G472), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n523), .A2(new_n525), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n516), .B1(new_n538), .B2(new_n539), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n527), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n529), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n529), .A2(new_n544), .A3(new_n548), .A4(KEYINPUT71), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT22), .B(G137), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n305), .A2(G221), .A3(G234), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT24), .B(G110), .Z(new_n557));
  XNOR2_X1  g371(.A(G119), .B(G128), .ZN(new_n558));
  OR3_X1    g372(.A1(new_n557), .A2(KEYINPUT73), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT73), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n253), .A2(KEYINPUT23), .A3(G119), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n215), .A2(G128), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n215), .A2(G128), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n561), .B(new_n562), .C1(new_n563), .C2(KEYINPUT23), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n559), .B(new_n560), .C1(G110), .C2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n326), .A3(new_n339), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n348), .A2(new_n326), .B1(new_n558), .B2(new_n557), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT72), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G110), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n567), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT74), .B1(new_n566), .B2(new_n572), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n556), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n556), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n573), .B2(new_n574), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT75), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n580), .A2(new_n581), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n577), .A2(new_n586), .A3(new_n579), .A4(new_n582), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n462), .B1(G234), .B2(new_n380), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n577), .A2(new_n579), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n588), .A2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(KEYINPUT76), .B1(new_n553), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT76), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n596), .B(new_n593), .C1(new_n551), .C2(new_n552), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n487), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  NOR2_X1   g413(.A1(new_n464), .A2(new_n465), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT33), .Z(new_n601));
  NOR2_X1   g415(.A1(new_n469), .A2(G902), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n468), .A2(new_n471), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n601), .A2(new_n602), .B1(new_n603), .B2(new_n469), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n281), .A2(new_n292), .A3(new_n187), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n187), .B1(new_n281), .B2(new_n292), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n300), .B(new_n485), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  AOI211_X1 g421(.A(new_n604), .B(new_n607), .C1(new_n382), .C2(new_n389), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n547), .A2(new_n380), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G472), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n547), .A2(new_n527), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n594), .A2(new_n438), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n376), .A2(KEYINPUT20), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n373), .A2(new_n375), .A3(new_n369), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n381), .B(new_n475), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n300), .ZN(new_n620));
  INV_X1    g434(.A(new_n606), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n298), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n485), .B(KEYINPUT97), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n619), .A2(KEYINPUT98), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n625));
  INV_X1    g439(.A(new_n618), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n384), .B(new_n474), .C1(new_n388), .C2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n300), .B(new_n623), .C1(new_n605), .C2(new_n606), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n613), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT99), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n578), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n573), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n591), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n589), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n610), .A2(new_n438), .A3(new_n611), .A4(new_n638), .ZN(new_n639));
  NOR4_X1   g453(.A1(new_n301), .A2(new_n639), .A3(new_n390), .A4(new_n486), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT100), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n640), .B(new_n642), .ZN(G12));
  NAND3_X1  g457(.A1(new_n483), .A2(G902), .A3(G953), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT101), .B1(new_n644), .B2(G900), .ZN(new_n645));
  OR3_X1    g459(.A1(new_n644), .A2(KEYINPUT101), .A3(G900), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n481), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n627), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n622), .A2(new_n638), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n553), .A2(new_n438), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XNOR2_X1  g467(.A(new_n647), .B(KEYINPUT39), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n438), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT40), .Z(new_n656));
  AOI211_X1 g470(.A(new_n620), .B(new_n475), .C1(new_n382), .C2(new_n389), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n299), .A2(KEYINPUT38), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT38), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n297), .A2(new_n659), .A3(new_n298), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n522), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n516), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n380), .B1(new_n533), .B2(new_n524), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n529), .A2(new_n548), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n638), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n656), .A2(new_n657), .A3(new_n661), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  AOI211_X1 g484(.A(new_n604), .B(new_n648), .C1(new_n382), .C2(new_n389), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n553), .A2(new_n671), .A3(new_n438), .A4(new_n651), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  OAI21_X1  g487(.A(new_n380), .B1(new_n435), .B2(new_n436), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G469), .ZN(new_n675));
  INV_X1    g489(.A(new_n393), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n675), .A2(new_n676), .A3(new_n437), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n553), .A2(new_n608), .A3(new_n594), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT41), .B(G113), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G15));
  NAND4_X1  g494(.A1(new_n553), .A2(new_n630), .A3(new_n594), .A4(new_n677), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G116), .ZN(G18));
  NOR2_X1   g496(.A1(new_n390), .A2(new_n486), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n553), .A2(new_n683), .A3(new_n651), .A4(new_n677), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  OR2_X1    g499(.A1(new_n534), .A2(new_n524), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n528), .B1(new_n686), .B2(new_n545), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n609), .B2(G472), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n688), .A2(new_n594), .A3(new_n623), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n677), .A2(new_n622), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n390), .A4(new_n474), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  INV_X1    g506(.A(new_n604), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n390), .A2(new_n693), .A3(new_n647), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n677), .A2(new_n688), .A3(new_n622), .A4(new_n638), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n266), .ZN(G27));
  AND4_X1   g511(.A1(new_n438), .A2(new_n297), .A3(new_n300), .A4(new_n298), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n604), .B1(new_n382), .B2(new_n389), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n698), .A2(new_n699), .A3(new_n647), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n548), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n547), .A2(KEYINPUT103), .A3(KEYINPUT32), .A4(new_n527), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n529), .A3(new_n544), .A4(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n594), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n700), .A2(KEYINPUT104), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT104), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n698), .A2(new_n699), .A3(new_n647), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n594), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n553), .A2(new_n671), .A3(new_n594), .A4(new_n698), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n712));
  AOI22_X1  g526(.A1(new_n706), .A2(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT105), .B(G131), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G33));
  NAND4_X1  g529(.A1(new_n553), .A2(new_n594), .A3(new_n649), .A4(new_n698), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G134), .ZN(G36));
  AND2_X1   g531(.A1(new_n382), .A2(new_n389), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n693), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT43), .ZN(new_n720));
  OR3_X1    g534(.A1(new_n390), .A2(KEYINPUT43), .A3(new_n604), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n638), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n611), .B2(new_n610), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(KEYINPUT44), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT106), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT44), .B1(new_n722), .B2(new_n724), .ZN(new_n727));
  INV_X1    g541(.A(new_n437), .ZN(new_n728));
  INV_X1    g542(.A(new_n395), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n431), .A2(KEYINPUT45), .ZN(new_n730));
  OAI21_X1  g544(.A(G469), .B1(new_n431), .B2(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n728), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n733), .B2(new_n732), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(new_n676), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n297), .A2(new_n300), .A3(new_n298), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n736), .A2(new_n654), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n727), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n726), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G137), .ZN(G39));
  NAND2_X1  g556(.A1(new_n735), .A2(new_n676), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(KEYINPUT107), .B2(KEYINPUT47), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n745));
  OAI21_X1  g559(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n551), .A2(new_n738), .A3(new_n552), .A4(new_n593), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n746), .A2(new_n694), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n319), .ZN(G42));
  INV_X1    g563(.A(KEYINPUT118), .ZN(new_n750));
  NOR2_X1   g564(.A1(G952), .A2(G953), .ZN(new_n751));
  INV_X1    g565(.A(new_n699), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n299), .A2(new_n300), .A3(new_n623), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n752), .A2(new_n753), .A3(new_n612), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n640), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n382), .A2(new_n389), .A3(new_n474), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT109), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n382), .A2(new_n389), .A3(new_n758), .A4(new_n474), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n761));
  INV_X1    g575(.A(new_n753), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n613), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n598), .B(new_n755), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n688), .A2(new_n638), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n671), .A2(new_n767), .A3(new_n698), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n381), .B1(new_n617), .B2(new_n618), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n638), .A2(new_n769), .A3(new_n475), .A4(new_n647), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n737), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n553), .A2(new_n438), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n716), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT111), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n716), .A2(new_n772), .A3(new_n768), .A4(KEYINPUT111), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n766), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n711), .A2(new_n712), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT104), .B1(new_n700), .B2(new_n705), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n708), .A2(new_n709), .A3(new_n707), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n678), .A2(new_n681), .A3(new_n684), .A4(new_n691), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n778), .B1(new_n784), .B2(KEYINPUT112), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n439), .B(new_n650), .C1(new_n551), .C2(new_n552), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n696), .B1(new_n786), .B2(new_n649), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n393), .B(new_n648), .C1(new_n432), .C2(new_n437), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n666), .A2(new_n788), .A3(new_n723), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n621), .A2(new_n298), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n657), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(KEYINPUT52), .A3(new_n672), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n671), .A2(new_n690), .A3(new_n767), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n672), .A2(new_n652), .A3(new_n793), .A4(new_n791), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n681), .A2(new_n678), .A3(new_n684), .A4(new_n691), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n713), .A2(KEYINPUT112), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n777), .A2(new_n785), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  AOI211_X1 g614(.A(KEYINPUT110), .B(new_n753), .C1(new_n757), .C2(new_n759), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n765), .A2(new_n801), .A3(new_n612), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n598), .A2(new_n755), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n713), .A2(new_n798), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n775), .A2(new_n776), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n797), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n778), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n800), .A2(new_n808), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n800), .A2(new_n808), .A3(new_n810), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n805), .A4(new_n797), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n810), .B1(new_n814), .B2(new_n808), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n811), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n738), .A2(new_n677), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n722), .A2(new_n480), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n704), .A2(new_n594), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n594), .A2(new_n817), .A3(new_n480), .A4(new_n667), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n479), .B1(new_n824), .B2(new_n699), .ZN(new_n825));
  INV_X1    g639(.A(new_n690), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n688), .A2(new_n594), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n720), .A2(new_n480), .A3(new_n827), .A4(new_n721), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n822), .A2(new_n823), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n658), .A2(new_n620), .A3(new_n660), .A4(new_n677), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT115), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n833), .B2(new_n828), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT50), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n836));
  OAI211_X1 g650(.A(KEYINPUT116), .B(new_n836), .C1(new_n833), .C2(new_n828), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n818), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(new_n767), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n824), .A2(new_n718), .A3(new_n604), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(KEYINPUT114), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n767), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n841), .B1(new_n818), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n835), .B2(new_n837), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n675), .A2(new_n437), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT108), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n746), .B1(new_n676), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n828), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n738), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n847), .A2(new_n853), .A3(new_n856), .A4(new_n843), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n831), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n751), .B1(new_n816), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n849), .B(KEYINPUT49), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n593), .A2(new_n393), .A3(new_n620), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n667), .A3(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(new_n661), .A3(new_n719), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n750), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n863), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n842), .A2(new_n843), .B1(new_n847), .B2(new_n853), .ZN(new_n866));
  INV_X1    g680(.A(new_n857), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n830), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n814), .A2(new_n808), .ZN(new_n869));
  OAI211_X1 g683(.A(KEYINPUT113), .B(new_n812), .C1(new_n869), .C2(new_n810), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n870), .B2(new_n811), .ZN(new_n871));
  OAI211_X1 g685(.A(KEYINPUT118), .B(new_n865), .C1(new_n871), .C2(new_n751), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n864), .A2(new_n872), .ZN(G75));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n237), .A2(new_n280), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(new_n278), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n800), .A2(new_n808), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(G902), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n874), .B(new_n877), .C1(new_n879), .C2(new_n188), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT119), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n305), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n879), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(G210), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(new_n877), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n881), .A2(new_n886), .ZN(G51));
  NAND2_X1  g701(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(new_n812), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n395), .B(KEYINPUT120), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT57), .ZN(new_n891));
  OAI22_X1  g705(.A1(new_n889), .A2(new_n891), .B1(new_n436), .B2(new_n435), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n730), .A2(new_n731), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT121), .Z(new_n894));
  NAND2_X1  g708(.A1(new_n884), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n882), .B1(new_n892), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n373), .A2(new_n375), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n883), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(G60));
  INV_X1    g714(.A(new_n601), .ZN(new_n901));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT59), .Z(new_n903));
  AOI211_X1 g717(.A(new_n901), .B(new_n903), .C1(new_n888), .C2(new_n812), .ZN(new_n904));
  INV_X1    g718(.A(new_n903), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n870), .A2(new_n811), .A3(new_n905), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n882), .B(new_n904), .C1(new_n901), .C2(new_n906), .ZN(G63));
  XNOR2_X1  g721(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n908));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n800), .B2(new_n808), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(new_n590), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n636), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n883), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n914), .B(new_n915), .ZN(G66));
  NAND2_X1  g730(.A1(new_n804), .A2(new_n783), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n305), .ZN(new_n918));
  OAI21_X1  g732(.A(G953), .B1(new_n482), .B2(new_n238), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT123), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n875), .B1(G898), .B2(new_n305), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(G69));
  AND2_X1   g737(.A1(new_n787), .A2(new_n672), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n669), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT62), .Z(new_n926));
  INV_X1    g740(.A(new_n748), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n737), .A2(new_n655), .ZN(new_n928));
  OAI221_X1 g742(.A(new_n928), .B1(new_n699), .B2(new_n760), .C1(new_n595), .C2(new_n597), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n926), .A2(new_n741), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n305), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n519), .A2(new_n520), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n331), .B(KEYINPUT124), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n657), .A2(new_n790), .ZN(new_n936));
  INV_X1    g750(.A(new_n819), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n736), .A2(new_n654), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n924), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n939), .B(new_n748), .C1(new_n726), .C2(new_n740), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n782), .A2(new_n716), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT126), .Z(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n305), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n934), .B1(G900), .B2(G953), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n935), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n305), .B1(G227), .B2(G900), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n935), .B(new_n945), .C1(new_n948), .C2(new_n947), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(G72));
  OR3_X1    g766(.A1(new_n930), .A2(new_n516), .A3(new_n662), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n940), .A2(new_n516), .A3(new_n662), .A4(new_n942), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n917), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n522), .B(new_n516), .ZN(new_n956));
  XOR2_X1   g770(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n957));
  NAND2_X1  g771(.A1(G472), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n869), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n883), .B1(new_n956), .B2(new_n959), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n955), .A2(new_n961), .A3(new_n962), .ZN(G57));
endmodule


