//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT27), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT64), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n196), .A3(G143), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n197), .A2(new_n198), .A3(G128), .A4(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n202), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n194), .A2(new_n196), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(new_n204), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n201), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT11), .A3(G134), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(G137), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n215), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G137), .ZN(new_n218));
  OAI21_X1  g032(.A(G131), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n208), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n205), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G146), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G143), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n197), .A2(new_n200), .A3(new_n224), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n211), .A2(new_n213), .A3(new_n215), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n229), .A2(G131), .ZN(new_n230));
  INV_X1    g044(.A(new_n216), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n227), .B(new_n228), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  XOR2_X1   g046(.A(KEYINPUT2), .B(G113), .Z(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n233), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  OR2_X1    g053(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n234), .B1(new_n233), .B2(new_n239), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n237), .A2(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n220), .A2(new_n232), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n242), .B1(new_n220), .B2(new_n232), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT28), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT28), .ZN(new_n247));
  INV_X1    g061(.A(new_n242), .ZN(new_n248));
  INV_X1    g062(.A(new_n232), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n219), .A2(new_n216), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n198), .B1(new_n222), .B2(G143), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n223), .B1(new_n251), .B2(new_n202), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n252), .B2(new_n201), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n248), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n220), .A2(new_n242), .A3(new_n232), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n247), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n246), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n247), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n192), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n220), .A2(new_n262), .A3(new_n232), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n220), .B2(new_n232), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n248), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT67), .B(KEYINPUT31), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n266), .A2(new_n255), .A3(new_n192), .A4(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT30), .B1(new_n249), .B2(new_n253), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n242), .B1(new_n270), .B2(new_n263), .ZN(new_n271));
  INV_X1    g085(.A(new_n192), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n271), .A2(new_n243), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n269), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n187), .B1(new_n261), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n187), .C1(new_n261), .C2(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n272), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n245), .A2(new_n260), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n245), .A2(KEYINPUT70), .A3(new_n260), .A4(new_n283), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n256), .A2(new_n257), .ZN(new_n291));
  AOI211_X1 g105(.A(KEYINPUT68), .B(new_n247), .C1(new_n254), .C2(new_n255), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n260), .B(new_n192), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n294), .B(new_n272), .C1(new_n271), .C2(new_n243), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n270), .A2(new_n263), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n243), .B1(new_n296), .B2(new_n248), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT69), .B1(new_n297), .B2(new_n192), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n293), .A2(new_n282), .A3(new_n295), .A4(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n286), .A2(new_n300), .A3(new_n287), .A4(new_n288), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n290), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G472), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n281), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT73), .ZN(new_n309));
  OR3_X1    g123(.A1(new_n307), .A2(KEYINPUT73), .A3(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT16), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT16), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G146), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n306), .A2(new_n308), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n222), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n202), .A2(KEYINPUT23), .A3(G119), .ZN(new_n318));
  INV_X1    g132(.A(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G128), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n202), .A2(G119), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n318), .B(new_n320), .C1(new_n322), .C2(KEYINPUT23), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n320), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT24), .B(G110), .Z(new_n325));
  OAI22_X1  g139(.A1(new_n323), .A2(G110), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n315), .A2(new_n317), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(G110), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n325), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n311), .A2(new_n193), .A3(new_n313), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n315), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G953), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(G221), .A3(G234), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n334), .B(KEYINPUT74), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT22), .B(G137), .ZN(new_n336));
  XOR2_X1   g150(.A(new_n335), .B(new_n336), .Z(new_n337));
  NOR3_X1   g151(.A1(new_n327), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n335), .B(new_n336), .ZN(new_n339));
  INV_X1    g153(.A(new_n331), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n193), .B1(new_n311), .B2(new_n313), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n328), .B(new_n329), .C1(new_n340), .C2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n315), .A2(new_n317), .A3(new_n326), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n287), .B1(new_n338), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT75), .A3(KEYINPUT25), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT25), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n337), .B1(new_n327), .B2(new_n332), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n343), .A3(new_n339), .ZN(new_n349));
  AOI21_X1  g163(.A(G902), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n347), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT72), .B(G217), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(G234), .B2(new_n287), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n346), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n348), .A2(new_n349), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(G902), .ZN(new_n358));
  XOR2_X1   g172(.A(KEYINPUT76), .B(KEYINPUT77), .Z(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT78), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n356), .A2(new_n364), .A3(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT79), .B1(new_n304), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n369), .B(new_n366), .C1(new_n281), .C2(new_n303), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n333), .A2(G227), .ZN(new_n374));
  XOR2_X1   g188(.A(new_n373), .B(new_n374), .Z(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(KEYINPUT3), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT81), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT81), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n378), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(KEYINPUT81), .B(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT82), .A3(new_n378), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT80), .B(G104), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT3), .B1(new_n388), .B2(G107), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n377), .A2(KEYINPUT80), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G104), .ZN(new_n392));
  AOI21_X1  g206(.A(G107), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n385), .B(new_n387), .C1(new_n389), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G101), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n392), .A3(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n390), .A2(new_n392), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n379), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n401), .A2(new_n402), .A3(new_n385), .A4(new_n387), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n395), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n227), .A2(new_n228), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT82), .B1(new_n386), .B2(new_n378), .ZN(new_n407));
  AND4_X1   g221(.A1(KEYINPUT82), .A2(new_n378), .A3(new_n380), .A4(new_n382), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n402), .B1(new_n409), .B2(new_n401), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT83), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n394), .A2(KEYINPUT83), .A3(new_n411), .A4(G101), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n404), .B(new_n406), .C1(new_n412), .C2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n230), .A2(new_n231), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n386), .A2(G104), .ZN(new_n417));
  OAI21_X1  g231(.A(G101), .B1(new_n417), .B2(new_n393), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n403), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n421), .B1(new_n252), .B2(new_n201), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n199), .B1(new_n222), .B2(G143), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n202), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n201), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n418), .B(new_n425), .C1(new_n394), .C2(G101), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n420), .A2(new_n422), .B1(new_n426), .B2(new_n421), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n415), .A2(new_n416), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(KEYINPUT84), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n415), .A2(new_n430), .A3(new_n427), .A4(new_n416), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n426), .A2(new_n421), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n422), .A2(new_n418), .A3(new_n403), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n394), .A2(new_n411), .A3(G101), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n385), .A2(new_n387), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n393), .B1(new_n397), .B2(new_n396), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n411), .B1(new_n441), .B2(new_n402), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n438), .A2(new_n413), .B1(new_n442), .B2(new_n395), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n435), .B1(new_n443), .B2(new_n406), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n444), .A2(new_n416), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n376), .B1(new_n432), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n416), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n403), .A2(new_n418), .A3(new_n425), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n208), .B1(new_n403), .B2(new_n418), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT12), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT12), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n452), .B(new_n447), .C1(new_n448), .C2(new_n449), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n375), .B(new_n454), .C1(new_n429), .C2(new_n431), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n372), .B(new_n287), .C1(new_n446), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(G469), .A2(G902), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n432), .A2(new_n445), .A3(new_n376), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n454), .B1(new_n429), .B2(new_n431), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n458), .B(G469), .C1(new_n376), .C2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(new_n457), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G221), .ZN(new_n462));
  XOR2_X1   g276(.A(KEYINPUT9), .B(G234), .Z(new_n463));
  AOI21_X1  g277(.A(new_n462), .B1(new_n463), .B2(new_n287), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(G214), .B1(G237), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n248), .B(new_n404), .C1(new_n412), .C2(new_n414), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n237), .A2(new_n238), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n319), .A2(G116), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n472), .B(G113), .C1(KEYINPUT5), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n419), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G110), .B(G122), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(new_n478), .A3(new_n476), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT6), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n477), .A2(new_n483), .A3(new_n479), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n208), .A2(new_n307), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n307), .B2(new_n405), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n333), .A2(G224), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n487), .A2(KEYINPUT7), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n486), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n419), .B(new_n475), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n478), .B(KEYINPUT8), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(G902), .B1(new_n494), .B2(new_n481), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G210), .B1(G237), .B2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n497), .A3(new_n495), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n469), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g320(.A1(KEYINPUT18), .A2(G131), .ZN(new_n507));
  INV_X1    g321(.A(G237), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n333), .A3(G214), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n204), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT85), .A3(new_n503), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n309), .A2(G146), .A3(new_n310), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n317), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n504), .A2(new_n505), .ZN(new_n515));
  INV_X1    g329(.A(new_n507), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT86), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n510), .A2(new_n503), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n518), .A2(new_n519), .A3(new_n507), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n512), .B(new_n514), .C1(new_n517), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT19), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n309), .B2(new_n310), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n316), .A2(KEYINPUT19), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n222), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(G131), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n510), .A2(new_n214), .A3(new_n503), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n315), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n531));
  XNOR2_X1  g345(.A(G113), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(new_n377), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n526), .A2(new_n536), .A3(new_n527), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n518), .A2(KEYINPUT17), .A3(G131), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n315), .A2(new_n537), .A3(new_n331), .A4(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n521), .A3(new_n533), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n531), .B1(new_n530), .B2(new_n534), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(KEYINPUT20), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT20), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n544), .C1(new_n541), .C2(new_n542), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n539), .A2(new_n521), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n534), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n540), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n287), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G475), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G952), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  NAND2_X1  g371(.A1(G234), .A2(G237), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n559), .B(KEYINPUT90), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT21), .B(G898), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(KEYINPUT91), .Z(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n558), .A2(G902), .A3(G953), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n561), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(G116), .B(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n386), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n570));
  XNOR2_X1  g384(.A(G128), .B(G143), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n204), .A2(G128), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(G134), .C1(new_n570), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n210), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n571), .B(new_n210), .ZN(new_n577));
  INV_X1    g391(.A(G116), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(KEYINPUT14), .A3(G122), .ZN(new_n579));
  INV_X1    g393(.A(new_n568), .ZN(new_n580));
  OAI211_X1 g394(.A(G107), .B(new_n579), .C1(new_n580), .C2(KEYINPUT14), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n386), .A2(new_n568), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n463), .A2(new_n333), .A3(new_n353), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n576), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n576), .A2(new_n583), .A3(KEYINPUT89), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n583), .ZN(new_n589));
  INV_X1    g403(.A(new_n584), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n287), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT15), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(G478), .ZN(new_n595));
  INV_X1    g409(.A(G478), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n592), .B(new_n287), .C1(KEYINPUT15), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n555), .A2(new_n567), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n467), .A2(new_n501), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n371), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n402), .ZN(G3));
  AND3_X1   g416(.A1(new_n489), .A2(new_n497), .A3(new_n495), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n497), .B1(new_n489), .B2(new_n495), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n585), .A2(KEYINPUT33), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n592), .A2(new_n606), .B1(new_n591), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n596), .A2(G902), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n593), .A2(new_n596), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n555), .A2(new_n613), .ZN(new_n614));
  NOR4_X1   g428(.A1(new_n605), .A2(new_n469), .A3(new_n567), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n266), .A2(new_n255), .A3(new_n192), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n274), .B2(KEYINPUT31), .ZN(new_n617));
  AOI22_X1  g431(.A1(new_n246), .A2(new_n258), .B1(new_n247), .B2(new_n255), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n617), .B(new_n269), .C1(new_n618), .C2(new_n192), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n287), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G472), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n367), .A2(new_n277), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n615), .A2(new_n467), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n377), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  NAND3_X1  g440(.A1(new_n546), .A2(KEYINPUT93), .A3(new_n548), .ZN(new_n627));
  INV_X1    g441(.A(new_n567), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT93), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(KEYINPUT20), .C1(new_n543), .C2(new_n545), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n595), .A2(new_n597), .B1(new_n553), .B2(G475), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n627), .A2(new_n628), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT94), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n467), .A2(new_n501), .A3(new_n622), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT95), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT35), .B(G107), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G9));
  AND2_X1   g454(.A1(new_n621), .A2(new_n277), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n342), .A2(new_n343), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n339), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n360), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n356), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n600), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT37), .B(G110), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT96), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n651), .A2(KEYINPUT96), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n566), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n560), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n627), .A2(new_n630), .A3(new_n631), .A4(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n304), .A2(new_n646), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n501), .A2(new_n461), .A3(new_n465), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n202), .ZN(G30));
  XNOR2_X1  g475(.A(new_n605), .B(KEYINPUT38), .ZN(new_n662));
  INV_X1    g476(.A(G472), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n254), .A2(new_n255), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n663), .B1(new_n664), .B2(new_n272), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n616), .A2(new_n665), .B1(G472), .B2(G902), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT97), .ZN(new_n667));
  INV_X1    g481(.A(new_n280), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n279), .B1(new_n619), .B2(new_n187), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n646), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n554), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n546), .B2(new_n548), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n598), .A2(new_n468), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OR3_X1    g491(.A1(new_n662), .A2(new_n672), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT98), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n655), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n467), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT99), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(KEYINPUT40), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  INV_X1    g501(.A(new_n655), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n674), .A2(new_n612), .A3(new_n688), .ZN(new_n689));
  OAI211_X1 g503(.A(new_n689), .B(new_n468), .C1(new_n603), .C2(new_n604), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n304), .A2(new_n646), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n693), .A2(new_n466), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  AOI21_X1  g510(.A(new_n366), .B1(new_n281), .B2(new_n303), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n287), .B1(new_n446), .B2(new_n455), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(G469), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(new_n465), .A3(new_n456), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n615), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(KEYINPUT41), .B(G113), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G15));
  NOR3_X1   g517(.A1(new_n634), .A2(new_n635), .A3(new_n366), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n704), .A2(new_n700), .A3(new_n501), .A4(new_n304), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G116), .ZN(G18));
  AND2_X1   g520(.A1(new_n599), .A2(new_n646), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n700), .A2(new_n707), .A3(new_n501), .A4(new_n304), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G119), .ZN(G21));
  INV_X1    g523(.A(new_n362), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n192), .B1(new_n245), .B2(new_n260), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n187), .B1(new_n276), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n276), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n260), .B1(new_n291), .B2(new_n292), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n272), .ZN(new_n715));
  AOI21_X1  g529(.A(G902), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n710), .B(new_n712), .C1(new_n716), .C2(new_n663), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT101), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n621), .A2(new_n719), .A3(new_n710), .A4(new_n712), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n676), .B(new_n628), .C1(new_n603), .C2(new_n604), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(new_n700), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NAND3_X1  g539(.A1(new_n699), .A2(new_n465), .A3(new_n456), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n499), .A2(new_n500), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n468), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT102), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n689), .A2(new_n621), .A3(new_n646), .A4(new_n712), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n501), .A2(new_n465), .A3(new_n456), .A4(new_n699), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT102), .B1(new_n734), .B2(new_n731), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  NOR3_X1   g551(.A1(new_n603), .A2(new_n604), .A3(new_n469), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n456), .A2(new_n457), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n458), .B(KEYINPUT103), .C1(new_n376), .C2(new_n459), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n432), .A2(new_n445), .A3(new_n741), .A4(new_n376), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n372), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n738), .B(new_n465), .C1(new_n739), .C2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n741), .A2(new_n432), .A3(new_n445), .A4(new_n376), .ZN(new_n747));
  INV_X1    g561(.A(new_n454), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n430), .B1(new_n444), .B2(new_n416), .ZN(new_n749));
  INV_X1    g563(.A(new_n431), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n741), .B1(new_n751), .B2(new_n375), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n747), .B1(new_n752), .B2(new_n458), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n456), .B(new_n457), .C1(new_n753), .C2(new_n372), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT104), .A3(new_n465), .A4(new_n738), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n746), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n304), .ZN(new_n757));
  INV_X1    g571(.A(new_n689), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n362), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n697), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n761), .B1(new_n746), .B2(new_n755), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n760), .A2(KEYINPUT42), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(KEYINPUT105), .B(G131), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G33));
  AOI211_X1 g580(.A(new_n761), .B(new_n656), .C1(new_n746), .C2(new_n755), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n210), .ZN(G36));
  NAND2_X1  g582(.A1(KEYINPUT45), .A2(G469), .ZN(new_n769));
  OAI21_X1  g583(.A(G469), .B1(new_n459), .B2(new_n376), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n432), .A2(new_n445), .A3(new_n376), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT106), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT103), .B1(new_n459), .B2(new_n376), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n742), .B1(new_n775), .B2(new_n771), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT45), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n460), .A2(KEYINPUT106), .A3(new_n769), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n457), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n457), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n456), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n465), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n674), .A2(new_n613), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT43), .B1(new_n787), .B2(KEYINPUT107), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n674), .A2(KEYINPUT108), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n674), .A2(KEYINPUT108), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n613), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n788), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n641), .A2(new_n671), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(KEYINPUT44), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT44), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n605), .A2(new_n468), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n786), .A2(new_n680), .A3(new_n797), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  NOR4_X1   g616(.A1(new_n799), .A2(new_n304), .A3(new_n367), .A4(new_n758), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT109), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n465), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT47), .B1(new_n784), .B2(new_n465), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  XOR2_X1   g622(.A(new_n655), .B(KEYINPUT112), .Z(new_n809));
  NAND3_X1  g623(.A1(new_n670), .A2(new_n671), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n727), .A2(new_n676), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n754), .A2(new_n465), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n692), .A2(new_n694), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n660), .B1(new_n733), .B2(new_n735), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n764), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n705), .A2(new_n701), .A3(new_n724), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n727), .A2(new_n468), .A3(new_n628), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n549), .A2(new_n631), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n614), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n467), .A2(new_n821), .A3(new_n622), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n708), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n762), .A2(new_n657), .ZN(new_n827));
  INV_X1    g641(.A(new_n600), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n368), .A2(new_n370), .ZN(new_n829));
  INV_X1    g643(.A(new_n647), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n673), .A2(new_n598), .A3(new_n688), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n738), .A2(new_n630), .A3(new_n627), .A4(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n693), .A3(new_n466), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n756), .B2(new_n732), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n826), .A2(new_n827), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n818), .A2(new_n836), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n658), .A2(new_n659), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n730), .B1(new_n729), .B2(new_n732), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n734), .A2(KEYINPUT102), .A3(new_n731), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n812), .A2(new_n813), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n736), .A2(KEYINPUT111), .A3(new_n838), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n695), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n837), .A2(new_n847), .A3(KEYINPUT53), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n731), .B1(new_n746), .B2(new_n755), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n767), .A2(new_n850), .A3(new_n834), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n600), .B1(new_n371), .B2(new_n647), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n852), .A2(new_n819), .A3(new_n825), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n851), .A2(new_n764), .A3(new_n853), .A4(new_n817), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n849), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n848), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT114), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n848), .A2(new_n856), .A3(new_n860), .A4(new_n857), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT53), .B1(new_n837), .B2(new_n847), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n854), .A2(new_n849), .A3(new_n855), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT54), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n726), .A2(new_n799), .A3(new_n560), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n757), .A2(new_n362), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n795), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT48), .Z(new_n868));
  NAND3_X1  g682(.A1(new_n795), .A2(new_n721), .A3(new_n561), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n670), .A2(new_n366), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  OAI221_X1 g685(.A(new_n557), .B1(new_n869), .B2(new_n734), .C1(new_n871), .C2(new_n614), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n869), .A2(new_n799), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n805), .A2(new_n806), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n699), .A2(new_n456), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n465), .B1(new_n877), .B2(KEYINPUT115), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(KEYINPUT115), .B2(new_n877), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n876), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n662), .B1(new_n881), .B2(KEYINPUT50), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n869), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n726), .A2(new_n468), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT117), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n871), .A2(new_n555), .A3(new_n613), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n621), .A2(new_n712), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n646), .A2(new_n865), .A3(new_n891), .A4(new_n795), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n883), .B(new_n885), .C1(KEYINPUT118), .C2(new_n887), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n889), .A2(new_n893), .A3(new_n894), .A4(KEYINPUT51), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n873), .B1(new_n880), .B2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT47), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n785), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n465), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n879), .B(KEYINPUT116), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n874), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n889), .A2(new_n894), .A3(new_n893), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT51), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n859), .A2(new_n861), .A3(new_n864), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n556), .A2(new_n333), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n877), .B(KEYINPUT49), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n710), .A2(new_n468), .A3(new_n465), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT110), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n911), .A2(new_n791), .A3(new_n670), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(new_n662), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n908), .A2(KEYINPUT119), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n333), .A2(G952), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT120), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n287), .B1(new_n848), .B2(new_n856), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n922), .B2(G210), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n482), .A2(new_n484), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(new_n488), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT55), .Z(new_n926));
  OR2_X1    g740(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n926), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n921), .B1(new_n927), .B2(new_n928), .ZN(G51));
  XOR2_X1   g743(.A(new_n457), .B(KEYINPUT57), .Z(new_n930));
  INV_X1    g744(.A(new_n858), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n857), .B1(new_n848), .B2(new_n856), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n446), .B2(new_n455), .ZN(new_n934));
  INV_X1    g748(.A(new_n779), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n922), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n919), .B1(new_n934), .B2(new_n936), .ZN(G54));
  NAND3_X1  g751(.A1(new_n922), .A2(KEYINPUT58), .A3(G475), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n938), .A2(new_n543), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n543), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n919), .ZN(G60));
  NAND3_X1  g755(.A1(new_n859), .A2(new_n861), .A3(new_n864), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT59), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n608), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n608), .B(new_n944), .C1(new_n931), .C2(new_n932), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n920), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(G63));
  NAND2_X1  g762(.A1(new_n848), .A2(new_n856), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT60), .Z(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n644), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n949), .A2(new_n951), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n920), .B(new_n952), .C1(new_n953), .C2(new_n357), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT61), .Z(G66));
  AOI21_X1  g769(.A(new_n333), .B1(new_n563), .B2(G224), .ZN(new_n956));
  INV_X1    g770(.A(new_n853), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(KEYINPUT121), .A3(new_n333), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT121), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n853), .B2(G953), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n956), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n924), .B1(G898), .B2(new_n333), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT122), .Z(new_n963));
  XOR2_X1   g777(.A(new_n961), .B(new_n963), .Z(G69));
  INV_X1    g778(.A(new_n811), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n786), .A2(new_n680), .A3(new_n965), .A4(new_n866), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n843), .A2(new_n695), .A3(new_n845), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n801), .A2(new_n764), .A3(new_n827), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n807), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n333), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n296), .B(KEYINPUT123), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n523), .A2(new_n524), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n972), .B(new_n976), .C1(G227), .C2(new_n333), .ZN(new_n977));
  OAI21_X1  g791(.A(G900), .B1(new_n976), .B2(G227), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(G953), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n683), .A2(new_n829), .A3(new_n738), .A4(new_n823), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n807), .A2(new_n801), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT124), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n686), .A2(new_n969), .A3(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n975), .A2(new_n333), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n977), .B(new_n979), .C1(new_n988), .C2(new_n989), .ZN(G72));
  NAND2_X1  g804(.A1(G472), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT63), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT126), .Z(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(new_n971), .B2(new_n957), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n272), .A3(new_n297), .ZN(new_n995));
  INV_X1    g809(.A(new_n919), .ZN(new_n996));
  INV_X1    g810(.A(new_n992), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n298), .A2(new_n295), .A3(new_n616), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n997), .B(new_n998), .C1(new_n862), .C2(new_n863), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n995), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n297), .A2(new_n272), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n988), .A2(new_n853), .ZN(new_n1002));
  INV_X1    g816(.A(new_n993), .ZN(new_n1003));
  OAI211_X1 g817(.A(KEYINPUT127), .B(new_n1001), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1003), .B1(new_n988), .B2(new_n853), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1001), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1000), .B1(new_n1004), .B2(new_n1008), .ZN(G57));
endmodule


