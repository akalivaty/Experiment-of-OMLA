

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U545 ( .A1(n721), .A2(G8), .ZN(n759) );
  NOR2_X1 U546 ( .A1(n635), .A2(G651), .ZN(n629) );
  NOR2_X2 U547 ( .A1(n950), .A2(n688), .ZN(n687) );
  NAND2_X1 U548 ( .A1(n764), .A2(n674), .ZN(n676) );
  XNOR2_X1 U549 ( .A(n744), .B(n743), .ZN(n762) );
  INV_X1 U550 ( .A(KEYINPUT102), .ZN(n743) );
  NOR2_X2 U551 ( .A1(G2105), .A2(G2104), .ZN(n511) );
  NOR2_X1 U552 ( .A1(G2104), .A2(n515), .ZN(n881) );
  NOR2_X2 U553 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X2 U554 ( .A1(n519), .A2(n518), .ZN(G164) );
  INV_X2 U555 ( .A(n693), .ZN(n721) );
  NOR2_X2 U556 ( .A1(G164), .A2(G1384), .ZN(n764) );
  OR2_X1 U557 ( .A1(n759), .A2(n758), .ZN(n510) );
  NAND2_X1 U558 ( .A1(n693), .A2(G2072), .ZN(n681) );
  INV_X1 U559 ( .A(KEYINPUT28), .ZN(n686) );
  AND2_X1 U560 ( .A1(n726), .A2(n729), .ZN(n728) );
  XNOR2_X1 U561 ( .A(n734), .B(KEYINPUT32), .ZN(n735) );
  INV_X1 U562 ( .A(KEYINPUT64), .ZN(n675) );
  OR2_X1 U563 ( .A1(n673), .A2(n672), .ZN(n763) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n511), .Z(n877) );
  NAND2_X1 U565 ( .A1(G138), .A2(n877), .ZN(n513) );
  INV_X1 U566 ( .A(G2105), .ZN(n515) );
  AND2_X1 U567 ( .A1(n515), .A2(G2104), .ZN(n876) );
  NAND2_X1 U568 ( .A1(G102), .A2(n876), .ZN(n512) );
  NAND2_X1 U569 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U570 ( .A(n514), .B(KEYINPUT90), .ZN(n519) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n880) );
  NAND2_X1 U572 ( .A1(G114), .A2(n880), .ZN(n517) );
  NAND2_X1 U573 ( .A1(G126), .A2(n881), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n618) );
  NAND2_X1 U576 ( .A1(G85), .A2(n618), .ZN(n521) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  INV_X1 U578 ( .A(G651), .ZN(n522) );
  NOR2_X1 U579 ( .A1(n635), .A2(n522), .ZN(n622) );
  NAND2_X1 U580 ( .A1(G72), .A2(n622), .ZN(n520) );
  NAND2_X1 U581 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U582 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n523), .Z(n633) );
  NAND2_X1 U584 ( .A1(G60), .A2(n633), .ZN(n525) );
  NAND2_X1 U585 ( .A1(G47), .A2(n629), .ZN(n524) );
  NAND2_X1 U586 ( .A1(n525), .A2(n524), .ZN(n526) );
  OR2_X1 U587 ( .A1(n527), .A2(n526), .ZN(G290) );
  NAND2_X1 U588 ( .A1(G64), .A2(n633), .ZN(n529) );
  NAND2_X1 U589 ( .A1(G52), .A2(n629), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n535) );
  NAND2_X1 U591 ( .A1(n622), .A2(G77), .ZN(n530) );
  XOR2_X1 U592 ( .A(KEYINPUT65), .B(n530), .Z(n532) );
  NAND2_X1 U593 ( .A1(n618), .A2(G90), .ZN(n531) );
  NAND2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(n533), .Z(n534) );
  NOR2_X1 U596 ( .A1(n535), .A2(n534), .ZN(G171) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U598 ( .A1(n876), .A2(G99), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(KEYINPUT78), .ZN(n538) );
  NAND2_X1 U600 ( .A1(G111), .A2(n880), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U602 ( .A(KEYINPUT79), .B(n539), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT18), .B(KEYINPUT76), .Z(n541) );
  NAND2_X1 U604 ( .A1(G123), .A2(n881), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G135), .A2(n877), .ZN(n542) );
  XNOR2_X1 U607 ( .A(KEYINPUT77), .B(n542), .ZN(n543) );
  NOR2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U610 ( .A(KEYINPUT80), .B(n547), .ZN(n990) );
  XNOR2_X1 U611 ( .A(n990), .B(G2096), .ZN(n548) );
  OR2_X1 U612 ( .A1(G2100), .A2(n548), .ZN(G156) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G120), .ZN(G236) );
  INV_X1 U616 ( .A(G108), .ZN(G238) );
  NAND2_X1 U617 ( .A1(n633), .A2(G63), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n549), .B(KEYINPUT74), .ZN(n551) );
  NAND2_X1 U619 ( .A1(G51), .A2(n629), .ZN(n550) );
  NAND2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U621 ( .A(KEYINPUT6), .B(n552), .ZN(n560) );
  XOR2_X1 U622 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n554) );
  NAND2_X1 U623 ( .A1(G89), .A2(n618), .ZN(n553) );
  XNOR2_X1 U624 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U625 ( .A(KEYINPUT72), .B(n555), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n622), .A2(G76), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U628 ( .A(n558), .B(KEYINPUT5), .Z(n559) );
  NOR2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT7), .B(n561), .Z(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT75), .B(n562), .Z(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n563) );
  XOR2_X1 U634 ( .A(n563), .B(KEYINPUT10), .Z(n814) );
  NAND2_X1 U635 ( .A1(n814), .A2(G567), .ZN(n564) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(KEYINPUT68), .Z(n566) );
  NAND2_X1 U638 ( .A1(G56), .A2(n633), .ZN(n565) );
  XNOR2_X1 U639 ( .A(n566), .B(n565), .ZN(n573) );
  XNOR2_X1 U640 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n618), .A2(G81), .ZN(n567) );
  XNOR2_X1 U642 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U643 ( .A1(G68), .A2(n622), .ZN(n568) );
  NAND2_X1 U644 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U645 ( .A(n571), .B(n570), .ZN(n572) );
  NOR2_X1 U646 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n629), .A2(G43), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n575), .A2(n574), .ZN(n949) );
  INV_X1 U649 ( .A(G860), .ZN(n597) );
  NOR2_X1 U650 ( .A1(n949), .A2(n597), .ZN(n576) );
  XOR2_X1 U651 ( .A(KEYINPUT70), .B(n576), .Z(G153) );
  INV_X1 U652 ( .A(G171), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n622), .A2(G79), .ZN(n583) );
  NAND2_X1 U655 ( .A1(G66), .A2(n633), .ZN(n578) );
  NAND2_X1 U656 ( .A1(G92), .A2(n618), .ZN(n577) );
  NAND2_X1 U657 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U658 ( .A1(G54), .A2(n629), .ZN(n579) );
  XNOR2_X1 U659 ( .A(KEYINPUT71), .B(n579), .ZN(n580) );
  NOR2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U661 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U662 ( .A(KEYINPUT15), .B(n584), .ZN(n963) );
  INV_X1 U663 ( .A(n963), .ZN(n699) );
  INV_X1 U664 ( .A(G868), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n699), .A2(n594), .ZN(n585) );
  NAND2_X1 U666 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G65), .A2(n633), .ZN(n588) );
  NAND2_X1 U668 ( .A1(G78), .A2(n622), .ZN(n587) );
  NAND2_X1 U669 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n618), .A2(G91), .ZN(n589) );
  XOR2_X1 U671 ( .A(KEYINPUT66), .B(n589), .Z(n590) );
  NOR2_X1 U672 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n629), .A2(G53), .ZN(n592) );
  NAND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(G299) );
  NOR2_X1 U675 ( .A1(G286), .A2(n594), .ZN(n596) );
  NOR2_X1 U676 ( .A1(G868), .A2(G299), .ZN(n595) );
  NOR2_X1 U677 ( .A1(n596), .A2(n595), .ZN(G297) );
  NAND2_X1 U678 ( .A1(n597), .A2(G559), .ZN(n598) );
  NAND2_X1 U679 ( .A1(n598), .A2(n963), .ZN(n599) );
  XNOR2_X1 U680 ( .A(n599), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n949), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n963), .A2(G868), .ZN(n600) );
  NOR2_X1 U683 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G67), .A2(n633), .ZN(n604) );
  NAND2_X1 U686 ( .A1(G55), .A2(n629), .ZN(n603) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G93), .A2(n618), .ZN(n606) );
  NAND2_X1 U689 ( .A1(G80), .A2(n622), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(n642) );
  NAND2_X1 U692 ( .A1(G559), .A2(n963), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n609), .B(n949), .ZN(n648) );
  NOR2_X1 U694 ( .A1(G860), .A2(n648), .ZN(n610) );
  XOR2_X1 U695 ( .A(KEYINPUT81), .B(n610), .Z(n611) );
  XNOR2_X1 U696 ( .A(n642), .B(n611), .ZN(G145) );
  NAND2_X1 U697 ( .A1(G88), .A2(n618), .ZN(n613) );
  NAND2_X1 U698 ( .A1(G75), .A2(n622), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U700 ( .A1(G62), .A2(n633), .ZN(n615) );
  NAND2_X1 U701 ( .A1(G50), .A2(n629), .ZN(n614) );
  NAND2_X1 U702 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U703 ( .A1(n617), .A2(n616), .ZN(G166) );
  INV_X1 U704 ( .A(G166), .ZN(G303) );
  NAND2_X1 U705 ( .A1(n629), .A2(G48), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G61), .A2(n633), .ZN(n620) );
  NAND2_X1 U707 ( .A1(G86), .A2(n618), .ZN(n619) );
  NAND2_X1 U708 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U709 ( .A(KEYINPUT84), .B(n621), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n622), .A2(G73), .ZN(n623) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U712 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U714 ( .A(KEYINPUT85), .B(n628), .Z(G305) );
  NAND2_X1 U715 ( .A1(G49), .A2(n629), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U719 ( .A(KEYINPUT82), .B(n634), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n635), .A2(G87), .ZN(n636) );
  XOR2_X1 U721 ( .A(KEYINPUT83), .B(n636), .Z(n637) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(G288) );
  NOR2_X1 U723 ( .A1(G868), .A2(n642), .ZN(n639) );
  XOR2_X1 U724 ( .A(n639), .B(KEYINPUT88), .Z(n651) );
  XNOR2_X1 U725 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n641) );
  XNOR2_X1 U726 ( .A(G290), .B(KEYINPUT19), .ZN(n640) );
  XNOR2_X1 U727 ( .A(n641), .B(n640), .ZN(n643) );
  XOR2_X1 U728 ( .A(n643), .B(n642), .Z(n645) );
  INV_X1 U729 ( .A(G299), .ZN(n950) );
  XOR2_X1 U730 ( .A(G303), .B(n950), .Z(n644) );
  XNOR2_X1 U731 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U732 ( .A(n646), .B(G305), .ZN(n647) );
  XNOR2_X1 U733 ( .A(n647), .B(G288), .ZN(n893) );
  XNOR2_X1 U734 ( .A(n893), .B(n648), .ZN(n649) );
  NAND2_X1 U735 ( .A1(G868), .A2(n649), .ZN(n650) );
  NAND2_X1 U736 ( .A1(n651), .A2(n650), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n652) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n652), .Z(n653) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n653), .ZN(n654) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n654), .ZN(n655) );
  NAND2_X1 U741 ( .A1(n655), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U743 ( .A(KEYINPUT67), .B(G132), .ZN(G219) );
  NOR2_X1 U744 ( .A1(G238), .A2(G236), .ZN(n656) );
  NAND2_X1 U745 ( .A1(G69), .A2(n656), .ZN(n657) );
  NOR2_X1 U746 ( .A1(n657), .A2(G237), .ZN(n658) );
  XNOR2_X1 U747 ( .A(n658), .B(KEYINPUT89), .ZN(n818) );
  NAND2_X1 U748 ( .A1(n818), .A2(G567), .ZN(n663) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n659) );
  XOR2_X1 U750 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U751 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U752 ( .A1(G96), .A2(n661), .ZN(n819) );
  NAND2_X1 U753 ( .A1(n819), .A2(G2106), .ZN(n662) );
  NAND2_X1 U754 ( .A1(n663), .A2(n662), .ZN(n851) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n664) );
  NOR2_X1 U756 ( .A1(n851), .A2(n664), .ZN(n817) );
  NAND2_X1 U757 ( .A1(n817), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(n880), .A2(G113), .ZN(n667) );
  NAND2_X1 U759 ( .A1(G101), .A2(n876), .ZN(n665) );
  XOR2_X1 U760 ( .A(KEYINPUT23), .B(n665), .Z(n666) );
  NAND2_X1 U761 ( .A1(n667), .A2(n666), .ZN(n673) );
  NAND2_X1 U762 ( .A1(G137), .A2(n877), .ZN(n669) );
  NAND2_X1 U763 ( .A1(G125), .A2(n881), .ZN(n668) );
  NAND2_X1 U764 ( .A1(n669), .A2(n668), .ZN(n671) );
  NOR2_X1 U765 ( .A1(n673), .A2(n671), .ZN(G160) );
  INV_X1 U766 ( .A(G40), .ZN(n670) );
  OR2_X1 U767 ( .A1(n671), .A2(n670), .ZN(n672) );
  INV_X1 U768 ( .A(n763), .ZN(n674) );
  XNOR2_X2 U769 ( .A(n676), .B(n675), .ZN(n693) );
  NOR2_X1 U770 ( .A1(n721), .A2(G2084), .ZN(n710) );
  NAND2_X1 U771 ( .A1(G8), .A2(n710), .ZN(n720) );
  NOR2_X1 U772 ( .A1(G1966), .A2(n759), .ZN(n718) );
  XOR2_X1 U773 ( .A(KEYINPUT25), .B(G2078), .Z(n934) );
  NOR2_X1 U774 ( .A1(n721), .A2(n934), .ZN(n677) );
  XNOR2_X1 U775 ( .A(n677), .B(KEYINPUT95), .ZN(n679) );
  INV_X1 U776 ( .A(G1961), .ZN(n835) );
  NAND2_X1 U777 ( .A1(n721), .A2(n835), .ZN(n678) );
  NAND2_X1 U778 ( .A1(n679), .A2(n678), .ZN(n709) );
  NAND2_X1 U779 ( .A1(n709), .A2(G171), .ZN(n708) );
  INV_X1 U780 ( .A(KEYINPUT96), .ZN(n685) );
  INV_X1 U781 ( .A(KEYINPUT27), .ZN(n680) );
  XNOR2_X1 U782 ( .A(n681), .B(n680), .ZN(n683) );
  NAND2_X1 U783 ( .A1(n721), .A2(G1956), .ZN(n682) );
  NAND2_X1 U784 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U785 ( .A(n685), .B(n684), .ZN(n688) );
  XNOR2_X1 U786 ( .A(n687), .B(n686), .ZN(n705) );
  NAND2_X1 U787 ( .A1(n950), .A2(n688), .ZN(n703) );
  NAND2_X1 U788 ( .A1(n693), .A2(G1996), .ZN(n689) );
  XNOR2_X1 U789 ( .A(n689), .B(KEYINPUT26), .ZN(n691) );
  NAND2_X1 U790 ( .A1(n721), .A2(G1341), .ZN(n690) );
  NAND2_X1 U791 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U792 ( .A1(n949), .A2(n692), .ZN(n697) );
  NAND2_X1 U793 ( .A1(G2067), .A2(n693), .ZN(n695) );
  NAND2_X1 U794 ( .A1(n721), .A2(G1348), .ZN(n694) );
  NAND2_X1 U795 ( .A1(n695), .A2(n694), .ZN(n698) );
  NOR2_X1 U796 ( .A1(n699), .A2(n698), .ZN(n696) );
  OR2_X1 U797 ( .A1(n697), .A2(n696), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U802 ( .A(KEYINPUT29), .B(n706), .Z(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n726) );
  NOR2_X1 U804 ( .A1(G171), .A2(n709), .ZN(n715) );
  NOR2_X1 U805 ( .A1(n718), .A2(n710), .ZN(n711) );
  NAND2_X1 U806 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U807 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U808 ( .A1(G168), .A2(n713), .ZN(n714) );
  NOR2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U810 ( .A(n716), .B(KEYINPUT31), .Z(n727) );
  AND2_X1 U811 ( .A1(n726), .A2(n727), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n738) );
  NOR2_X1 U814 ( .A1(n721), .A2(G2090), .ZN(n722) );
  XOR2_X1 U815 ( .A(KEYINPUT97), .B(n722), .Z(n724) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n759), .ZN(n723) );
  NOR2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n725), .A2(G303), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n733) );
  INV_X1 U820 ( .A(n729), .ZN(n730) );
  OR2_X1 U821 ( .A1(n730), .A2(G286), .ZN(n731) );
  AND2_X1 U822 ( .A1(G8), .A2(n731), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n736) );
  XOR2_X1 U824 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n734) );
  XNOR2_X1 U825 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n748) );
  NOR2_X1 U827 ( .A1(G2090), .A2(G303), .ZN(n739) );
  NAND2_X1 U828 ( .A1(G8), .A2(n739), .ZN(n740) );
  NAND2_X1 U829 ( .A1(n748), .A2(n740), .ZN(n741) );
  XOR2_X1 U830 ( .A(KEYINPUT101), .B(n741), .Z(n742) );
  NAND2_X1 U831 ( .A1(n742), .A2(n759), .ZN(n744) );
  XNOR2_X1 U832 ( .A(G1981), .B(G305), .ZN(n971) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n956) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U835 ( .A1(G288), .A2(G1976), .ZN(n745) );
  XOR2_X1 U836 ( .A(n745), .B(KEYINPUT100), .Z(n955) );
  INV_X1 U837 ( .A(n955), .ZN(n746) );
  NOR2_X1 U838 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U840 ( .A1(n956), .A2(n750), .ZN(n751) );
  NOR2_X1 U841 ( .A1(n751), .A2(n759), .ZN(n752) );
  NOR2_X1 U842 ( .A1(KEYINPUT33), .A2(n752), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n971), .A2(n753), .ZN(n756) );
  NOR2_X1 U844 ( .A1(n759), .A2(n955), .ZN(n754) );
  NAND2_X1 U845 ( .A1(KEYINPUT33), .A2(n754), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n760) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XOR2_X1 U848 ( .A(n757), .B(KEYINPUT24), .Z(n758) );
  NAND2_X1 U849 ( .A1(n760), .A2(n510), .ZN(n761) );
  NOR2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n797) );
  NOR2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n809) );
  NAND2_X1 U852 ( .A1(G104), .A2(n876), .ZN(n766) );
  NAND2_X1 U853 ( .A1(G140), .A2(n877), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U855 ( .A(KEYINPUT34), .B(n767), .ZN(n773) );
  NAND2_X1 U856 ( .A1(n880), .A2(G116), .ZN(n768) );
  XOR2_X1 U857 ( .A(KEYINPUT91), .B(n768), .Z(n770) );
  NAND2_X1 U858 ( .A1(n881), .A2(G128), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  XOR2_X1 U860 ( .A(n771), .B(KEYINPUT35), .Z(n772) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U862 ( .A(KEYINPUT36), .B(n774), .Z(n775) );
  XOR2_X1 U863 ( .A(KEYINPUT92), .B(n775), .Z(n890) );
  XNOR2_X1 U864 ( .A(G2067), .B(KEYINPUT37), .ZN(n806) );
  NOR2_X1 U865 ( .A1(n890), .A2(n806), .ZN(n985) );
  NAND2_X1 U866 ( .A1(n809), .A2(n985), .ZN(n804) );
  NAND2_X1 U867 ( .A1(G95), .A2(n876), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G107), .A2(n880), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G119), .A2(n881), .ZN(n778) );
  XNOR2_X1 U871 ( .A(KEYINPUT93), .B(n778), .ZN(n779) );
  NOR2_X1 U872 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n877), .A2(G131), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n859) );
  NAND2_X1 U875 ( .A1(G1991), .A2(n859), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G117), .A2(n880), .ZN(n784) );
  NAND2_X1 U877 ( .A1(G129), .A2(n881), .ZN(n783) );
  NAND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n876), .A2(G105), .ZN(n785) );
  XOR2_X1 U880 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U881 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n877), .A2(G141), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n873) );
  NAND2_X1 U884 ( .A1(G1996), .A2(n873), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n992) );
  NAND2_X1 U886 ( .A1(n992), .A2(n809), .ZN(n792) );
  XNOR2_X1 U887 ( .A(n792), .B(KEYINPUT94), .ZN(n794) );
  XNOR2_X1 U888 ( .A(G1986), .B(G290), .ZN(n952) );
  NAND2_X1 U889 ( .A1(n952), .A2(n809), .ZN(n793) );
  AND2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n804), .A2(n795), .ZN(n796) );
  XNOR2_X1 U892 ( .A(n798), .B(KEYINPUT103), .ZN(n811) );
  NOR2_X1 U893 ( .A1(n873), .A2(G1996), .ZN(n799) );
  XNOR2_X1 U894 ( .A(n799), .B(KEYINPUT104), .ZN(n1000) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n859), .ZN(n988) );
  NOR2_X1 U896 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n988), .A2(n800), .ZN(n801) );
  NOR2_X1 U898 ( .A1(n992), .A2(n801), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n1000), .A2(n802), .ZN(n803) );
  XNOR2_X1 U900 ( .A(n803), .B(KEYINPUT39), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n890), .A2(n806), .ZN(n984) );
  NAND2_X1 U903 ( .A1(n807), .A2(n984), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n813) );
  XOR2_X1 U906 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n812) );
  XNOR2_X1 U907 ( .A(n813), .B(n812), .ZN(G329) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n814), .ZN(G217) );
  INV_X1 U909 ( .A(n814), .ZN(G223) );
  AND2_X1 U910 ( .A1(G15), .A2(G2), .ZN(n815) );
  NAND2_X1 U911 ( .A1(G661), .A2(n815), .ZN(G259) );
  NAND2_X1 U912 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U913 ( .A1(n817), .A2(n816), .ZN(G188) );
  XOR2_X1 U914 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  INV_X1 U916 ( .A(G96), .ZN(G221) );
  NOR2_X1 U917 ( .A1(n819), .A2(n818), .ZN(G325) );
  INV_X1 U918 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U919 ( .A(G1348), .B(G2454), .ZN(n820) );
  XNOR2_X1 U920 ( .A(n820), .B(G2430), .ZN(n821) );
  XNOR2_X1 U921 ( .A(n821), .B(G1341), .ZN(n827) );
  XOR2_X1 U922 ( .A(G2443), .B(G2427), .Z(n823) );
  XNOR2_X1 U923 ( .A(G2438), .B(G2446), .ZN(n822) );
  XNOR2_X1 U924 ( .A(n823), .B(n822), .ZN(n825) );
  XOR2_X1 U925 ( .A(G2451), .B(G2435), .Z(n824) );
  XNOR2_X1 U926 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U927 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U928 ( .A1(n828), .A2(G14), .ZN(n829) );
  XNOR2_X1 U929 ( .A(KEYINPUT106), .B(n829), .ZN(n900) );
  XNOR2_X1 U930 ( .A(n900), .B(KEYINPUT107), .ZN(G401) );
  XOR2_X1 U931 ( .A(KEYINPUT111), .B(G1956), .Z(n831) );
  XNOR2_X1 U932 ( .A(G1996), .B(G1991), .ZN(n830) );
  XNOR2_X1 U933 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U934 ( .A(n832), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U935 ( .A(G1971), .B(G1966), .ZN(n833) );
  XNOR2_X1 U936 ( .A(n834), .B(n833), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n835), .B(G1976), .ZN(n837) );
  XNOR2_X1 U938 ( .A(G1986), .B(G1981), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U940 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U941 ( .A(G2474), .B(KEYINPUT110), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(G229) );
  XOR2_X1 U943 ( .A(G2678), .B(G2084), .Z(n843) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U946 ( .A(n844), .B(G2100), .Z(n846) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2072), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U949 ( .A(G2096), .B(KEYINPUT109), .Z(n848) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U952 ( .A(n850), .B(n849), .Z(G227) );
  INV_X1 U953 ( .A(n851), .ZN(G319) );
  NAND2_X1 U954 ( .A1(G124), .A2(n881), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n852), .B(KEYINPUT44), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n876), .A2(G100), .ZN(n853) );
  NAND2_X1 U957 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G136), .A2(n877), .ZN(n856) );
  NAND2_X1 U959 ( .A1(G112), .A2(n880), .ZN(n855) );
  NAND2_X1 U960 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U961 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U962 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n859), .B(KEYINPUT46), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n871) );
  NAND2_X1 U965 ( .A1(G118), .A2(n880), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G130), .A2(n881), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n876), .A2(G106), .ZN(n864) );
  XNOR2_X1 U969 ( .A(n864), .B(KEYINPUT112), .ZN(n866) );
  NAND2_X1 U970 ( .A1(G142), .A2(n877), .ZN(n865) );
  NAND2_X1 U971 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U972 ( .A(n867), .B(KEYINPUT45), .Z(n868) );
  NOR2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U974 ( .A(n871), .B(n870), .Z(n872) );
  XNOR2_X1 U975 ( .A(n990), .B(n872), .ZN(n875) );
  XNOR2_X1 U976 ( .A(n873), .B(G162), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n887) );
  NAND2_X1 U978 ( .A1(G103), .A2(n876), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G139), .A2(n877), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U981 ( .A1(G115), .A2(n880), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G127), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n995) );
  XOR2_X1 U986 ( .A(n887), .B(n995), .Z(n889) );
  XNOR2_X1 U987 ( .A(G164), .B(G160), .ZN(n888) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U990 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n893), .B(n949), .ZN(n894) );
  XOR2_X1 U992 ( .A(n894), .B(n963), .Z(n896) );
  XNOR2_X1 U993 ( .A(G171), .B(G286), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U995 ( .A1(G37), .A2(n897), .ZN(G397) );
  XNOR2_X1 U996 ( .A(KEYINPUT114), .B(KEYINPUT49), .ZN(n899) );
  NOR2_X1 U997 ( .A1(G229), .A2(G227), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n902) );
  NAND2_X1 U999 ( .A1(G319), .A2(n900), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(n904), .A2(n903), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1004 ( .A(KEYINPUT121), .B(G16), .Z(n930) );
  XOR2_X1 U1005 ( .A(G5), .B(G1961), .Z(n919) );
  XNOR2_X1 U1006 ( .A(G1966), .B(G21), .ZN(n917) );
  XNOR2_X1 U1007 ( .A(KEYINPUT59), .B(G1348), .ZN(n905) );
  XNOR2_X1 U1008 ( .A(n905), .B(G4), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(G1956), .B(G20), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(G1341), .B(G19), .ZN(n906) );
  XNOR2_X1 U1011 ( .A(n906), .B(KEYINPUT122), .ZN(n908) );
  XNOR2_X1 U1012 ( .A(G6), .B(G1981), .ZN(n907) );
  NOR2_X1 U1013 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1014 ( .A(KEYINPUT123), .B(n909), .ZN(n910) );
  NOR2_X1 U1015 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1016 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1017 ( .A(KEYINPUT60), .B(n914), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(KEYINPUT124), .B(n915), .ZN(n916) );
  NOR2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(n927) );
  XNOR2_X1 U1021 ( .A(G1986), .B(G24), .ZN(n921) );
  XNOR2_X1 U1022 ( .A(G23), .B(G1976), .ZN(n920) );
  NOR2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(G1971), .B(KEYINPUT125), .ZN(n922) );
  XNOR2_X1 U1025 ( .A(n922), .B(G22), .ZN(n923) );
  NAND2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(KEYINPUT58), .B(n925), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1029 ( .A(KEYINPUT61), .B(n928), .Z(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n982) );
  XOR2_X1 U1031 ( .A(G1991), .B(G25), .Z(n931) );
  NAND2_X1 U1032 ( .A1(n931), .A2(G28), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G1996), .B(G32), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(G33), .B(G2072), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(G2067), .B(G26), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G27), .B(n934), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1041 ( .A(KEYINPUT53), .B(n941), .Z(n944) );
  XOR2_X1 U1042 ( .A(KEYINPUT54), .B(G34), .Z(n942) );
  XNOR2_X1 U1043 ( .A(G2084), .B(n942), .ZN(n943) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(G35), .B(G2090), .ZN(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1047 ( .A(KEYINPUT55), .B(n947), .Z(n948) );
  NOR2_X1 U1048 ( .A1(G29), .A2(n948), .ZN(n979) );
  XNOR2_X1 U1049 ( .A(n949), .B(G1341), .ZN(n968) );
  XOR2_X1 U1050 ( .A(G1971), .B(G303), .Z(n954) );
  XOR2_X1 U1051 ( .A(G1956), .B(n950), .Z(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n959) );
  XOR2_X1 U1054 ( .A(KEYINPUT117), .B(n955), .Z(n957) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(n960), .B(KEYINPUT118), .ZN(n962) );
  XOR2_X1 U1058 ( .A(G301), .B(G1961), .Z(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1060 ( .A(G1348), .B(n963), .Z(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1062 ( .A(KEYINPUT119), .B(n966), .ZN(n967) );
  NOR2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1064 ( .A(KEYINPUT120), .B(n969), .Z(n974) );
  XOR2_X1 U1065 ( .A(G168), .B(G1966), .Z(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(KEYINPUT57), .B(n972), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1069 ( .A(G16), .B(KEYINPUT56), .Z(n975) );
  XNOR2_X1 U1070 ( .A(KEYINPUT116), .B(n975), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n980), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n983), .B(KEYINPUT126), .ZN(n1011) );
  INV_X1 U1076 ( .A(n984), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n994) );
  XOR2_X1 U1078 ( .A(G160), .B(G2084), .Z(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n1005) );
  XOR2_X1 U1083 ( .A(G2072), .B(n995), .Z(n997) );
  XOR2_X1 U1084 ( .A(G164), .B(G2078), .Z(n996) );
  NOR2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(KEYINPUT50), .B(n998), .ZN(n1003) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT51), .B(n1001), .Z(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(KEYINPUT52), .B(n1006), .Z(n1007) );
  NOR2_X1 U1093 ( .A1(KEYINPUT55), .A2(n1007), .ZN(n1008) );
  XNOR2_X1 U1094 ( .A(KEYINPUT115), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(G29), .ZN(n1010) );
  NAND2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1097 ( .A(KEYINPUT62), .B(n1012), .ZN(G150) );
  INV_X1 U1098 ( .A(G150), .ZN(G311) );
endmodule

