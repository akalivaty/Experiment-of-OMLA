

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U549 ( .A(n732), .ZN(n516) );
  AND2_X2 U550 ( .A1(n574), .A2(G2105), .ZN(n885) );
  NOR2_X2 U551 ( .A1(G2105), .A2(n574), .ZN(n890) );
  NOR2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n569) );
  XOR2_X1 U553 ( .A(KEYINPUT88), .B(n687), .Z(n517) );
  NOR2_X2 U554 ( .A1(n694), .A2(n693), .ZN(G164) );
  AND2_X1 U555 ( .A1(n780), .A2(n779), .ZN(n518) );
  OR2_X1 U556 ( .A1(n767), .A2(n778), .ZN(n519) );
  AND2_X1 U557 ( .A1(n1003), .A2(n830), .ZN(n520) );
  NAND2_X1 U558 ( .A1(n516), .A2(G1956), .ZN(n698) );
  INV_X1 U559 ( .A(KEYINPUT103), .ZN(n748) );
  INV_X1 U560 ( .A(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U561 ( .A1(n519), .A2(n935), .ZN(n768) );
  NOR2_X1 U562 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U563 ( .A1(n818), .A2(n520), .ZN(n819) );
  NOR2_X1 U564 ( .A1(G651), .A2(n648), .ZN(n647) );
  NOR2_X1 U565 ( .A1(G651), .A2(G543), .ZN(n521) );
  XOR2_X1 U566 ( .A(KEYINPUT65), .B(n521), .Z(n639) );
  NAND2_X1 U567 ( .A1(G89), .A2(n639), .ZN(n522) );
  XOR2_X1 U568 ( .A(KEYINPUT75), .B(n522), .Z(n523) );
  XNOR2_X1 U569 ( .A(n523), .B(KEYINPUT4), .ZN(n525) );
  XOR2_X1 U570 ( .A(KEYINPUT0), .B(G543), .Z(n648) );
  INV_X1 U571 ( .A(G651), .ZN(n527) );
  NOR2_X1 U572 ( .A1(n648), .A2(n527), .ZN(n636) );
  NAND2_X1 U573 ( .A1(G76), .A2(n636), .ZN(n524) );
  NAND2_X1 U574 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U575 ( .A(n526), .B(KEYINPUT5), .ZN(n533) );
  NOR2_X1 U576 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n528), .Z(n652) );
  NAND2_X1 U578 ( .A1(G63), .A2(n652), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G51), .A2(n647), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U581 ( .A(KEYINPUT6), .B(n531), .Z(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U583 ( .A(n534), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U584 ( .A(G168), .B(KEYINPUT8), .Z(n535) );
  XNOR2_X1 U585 ( .A(KEYINPUT76), .B(n535), .ZN(G286) );
  NAND2_X1 U586 ( .A1(n647), .A2(G53), .ZN(n542) );
  NAND2_X1 U587 ( .A1(G65), .A2(n652), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G78), .A2(n636), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n639), .A2(G91), .ZN(n538) );
  XOR2_X1 U591 ( .A(KEYINPUT70), .B(n538), .Z(n539) );
  NOR2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U593 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U594 ( .A(KEYINPUT71), .B(n543), .Z(G299) );
  NAND2_X1 U595 ( .A1(G85), .A2(n639), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G72), .A2(n636), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U598 ( .A1(G60), .A2(n652), .ZN(n547) );
  NAND2_X1 U599 ( .A1(G47), .A2(n647), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  OR2_X1 U601 ( .A1(n549), .A2(n548), .ZN(G290) );
  XOR2_X1 U602 ( .A(G2438), .B(G2435), .Z(n551) );
  XNOR2_X1 U603 ( .A(G2430), .B(G2454), .ZN(n550) );
  XNOR2_X1 U604 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U605 ( .A(n552), .B(KEYINPUT106), .Z(n554) );
  XNOR2_X1 U606 ( .A(G1348), .B(G1341), .ZN(n553) );
  XNOR2_X1 U607 ( .A(n554), .B(n553), .ZN(n558) );
  XOR2_X1 U608 ( .A(G2446), .B(KEYINPUT107), .Z(n556) );
  XNOR2_X1 U609 ( .A(G2451), .B(G2427), .ZN(n555) );
  XNOR2_X1 U610 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U611 ( .A(n558), .B(n557), .Z(n560) );
  XNOR2_X1 U612 ( .A(KEYINPUT105), .B(G2443), .ZN(n559) );
  XNOR2_X1 U613 ( .A(n560), .B(n559), .ZN(n561) );
  AND2_X1 U614 ( .A1(n561), .A2(G14), .ZN(G401) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G57), .ZN(G237) );
  NAND2_X1 U618 ( .A1(G62), .A2(n652), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G88), .A2(n639), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U621 ( .A1(G75), .A2(n636), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G50), .A2(n647), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U625 ( .A(KEYINPUT80), .B(n568), .Z(G303) );
  XOR2_X1 U626 ( .A(KEYINPUT66), .B(n569), .Z(n570) );
  XNOR2_X1 U627 ( .A(n570), .B(KEYINPUT17), .ZN(n689) );
  BUF_X1 U628 ( .A(n689), .Z(n893) );
  NAND2_X1 U629 ( .A1(G137), .A2(n893), .ZN(n573) );
  INV_X1 U630 ( .A(G2104), .ZN(n574) );
  NAND2_X1 U631 ( .A1(G101), .A2(n890), .ZN(n571) );
  XOR2_X1 U632 ( .A(KEYINPUT23), .B(n571), .Z(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U634 ( .A1(G125), .A2(n885), .ZN(n576) );
  AND2_X2 U635 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U636 ( .A1(G113), .A2(n886), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U638 ( .A1(n578), .A2(n577), .ZN(G160) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n834) );
  NAND2_X1 U642 ( .A1(n834), .A2(G567), .ZN(n580) );
  XNOR2_X1 U643 ( .A(n580), .B(KEYINPUT11), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT73), .B(n581), .ZN(G234) );
  NAND2_X1 U645 ( .A1(G56), .A2(n652), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n582), .Z(n588) );
  NAND2_X1 U647 ( .A1(n639), .A2(G81), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U649 ( .A1(G68), .A2(n636), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n586), .Z(n587) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n647), .A2(G43), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n930) );
  INV_X1 U655 ( .A(G860), .ZN(n613) );
  OR2_X1 U656 ( .A1(n930), .A2(n613), .ZN(G153) );
  NAND2_X1 U657 ( .A1(n636), .A2(G77), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n591), .B(KEYINPUT68), .ZN(n593) );
  NAND2_X1 U659 ( .A1(G90), .A2(n639), .ZN(n592) );
  NAND2_X1 U660 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U661 ( .A(n594), .B(KEYINPUT9), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G64), .A2(n652), .ZN(n596) );
  NAND2_X1 U663 ( .A1(G52), .A2(n647), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U665 ( .A(KEYINPUT67), .B(n597), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT69), .ZN(G171) );
  INV_X1 U668 ( .A(G171), .ZN(G301) );
  NAND2_X1 U669 ( .A1(G868), .A2(G301), .ZN(n601) );
  XNOR2_X1 U670 ( .A(n601), .B(KEYINPUT74), .ZN(n610) );
  INV_X1 U671 ( .A(G868), .ZN(n667) );
  NAND2_X1 U672 ( .A1(G66), .A2(n652), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G92), .A2(n639), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G79), .A2(n636), .ZN(n605) );
  NAND2_X1 U676 ( .A1(G54), .A2(n647), .ZN(n604) );
  NAND2_X1 U677 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U679 ( .A(KEYINPUT15), .B(n608), .Z(n925) );
  INV_X1 U680 ( .A(n925), .ZN(n904) );
  NAND2_X1 U681 ( .A1(n667), .A2(n904), .ZN(n609) );
  NAND2_X1 U682 ( .A1(n610), .A2(n609), .ZN(G284) );
  NAND2_X1 U683 ( .A1(G868), .A2(G286), .ZN(n612) );
  NAND2_X1 U684 ( .A1(G299), .A2(n667), .ZN(n611) );
  NAND2_X1 U685 ( .A1(n612), .A2(n611), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n613), .A2(G559), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n614), .A2(n925), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n930), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n925), .A2(G868), .ZN(n616) );
  NOR2_X1 U691 ( .A1(G559), .A2(n616), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(G282) );
  NAND2_X1 U693 ( .A1(n885), .A2(G123), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n619), .B(KEYINPUT18), .ZN(n621) );
  NAND2_X1 U695 ( .A1(G111), .A2(n886), .ZN(n620) );
  NAND2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U697 ( .A1(G99), .A2(n890), .ZN(n623) );
  NAND2_X1 U698 ( .A1(G135), .A2(n893), .ZN(n622) );
  NAND2_X1 U699 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n996) );
  XNOR2_X1 U701 ( .A(G2096), .B(n996), .ZN(n627) );
  INV_X1 U702 ( .A(G2100), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(G156) );
  NAND2_X1 U704 ( .A1(n925), .A2(G559), .ZN(n663) );
  XNOR2_X1 U705 ( .A(n930), .B(n663), .ZN(n628) );
  NOR2_X1 U706 ( .A1(n628), .A2(G860), .ZN(n635) );
  NAND2_X1 U707 ( .A1(G67), .A2(n652), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G93), .A2(n639), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G80), .A2(n636), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G55), .A2(n647), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  OR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n666) );
  XOR2_X1 U714 ( .A(n635), .B(n666), .Z(G145) );
  XOR2_X1 U715 ( .A(KEYINPUT2), .B(KEYINPUT79), .Z(n638) );
  NAND2_X1 U716 ( .A1(G73), .A2(n636), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n638), .B(n637), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G86), .A2(n639), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G48), .A2(n647), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n652), .A2(G61), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT78), .B(n642), .Z(n643) );
  NOR2_X1 U723 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U725 ( .A1(G651), .A2(G74), .ZN(n654) );
  NAND2_X1 U726 ( .A1(G49), .A2(n647), .ZN(n650) );
  NAND2_X1 U727 ( .A1(G87), .A2(n648), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U729 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U731 ( .A(KEYINPUT77), .B(n655), .Z(G288) );
  XNOR2_X1 U732 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n657) );
  INV_X1 U733 ( .A(G299), .ZN(n914) );
  XNOR2_X1 U734 ( .A(G290), .B(n914), .ZN(n656) );
  XNOR2_X1 U735 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U736 ( .A(n666), .B(n658), .Z(n660) );
  XNOR2_X1 U737 ( .A(n930), .B(G303), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(G305), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n662), .B(G288), .ZN(n906) );
  XNOR2_X1 U741 ( .A(KEYINPUT82), .B(n663), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n906), .B(n664), .ZN(n665) );
  NAND2_X1 U743 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U745 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n673), .A2(G2072), .ZN(n674) );
  XOR2_X1 U751 ( .A(KEYINPUT83), .B(n674), .Z(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U753 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G108), .A2(n676), .ZN(n840) );
  NAND2_X1 U757 ( .A1(G567), .A2(n840), .ZN(n683) );
  NOR2_X1 U758 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U759 ( .A(KEYINPUT84), .B(n677), .Z(n678) );
  XNOR2_X1 U760 ( .A(n678), .B(KEYINPUT22), .ZN(n679) );
  NOR2_X1 U761 ( .A1(G218), .A2(n679), .ZN(n680) );
  XOR2_X1 U762 ( .A(KEYINPUT85), .B(n680), .Z(n681) );
  NAND2_X1 U763 ( .A1(G96), .A2(n681), .ZN(n839) );
  NAND2_X1 U764 ( .A1(G2106), .A2(n839), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n683), .A2(n682), .ZN(n841) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n684) );
  XNOR2_X1 U767 ( .A(KEYINPUT86), .B(n684), .ZN(n685) );
  NOR2_X1 U768 ( .A1(n841), .A2(n685), .ZN(n837) );
  NAND2_X1 U769 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G126), .A2(n885), .ZN(n686) );
  XNOR2_X1 U771 ( .A(n686), .B(KEYINPUT87), .ZN(n688) );
  NAND2_X1 U772 ( .A1(G114), .A2(n886), .ZN(n687) );
  NOR2_X1 U773 ( .A1(n688), .A2(n517), .ZN(n691) );
  NAND2_X1 U774 ( .A1(n689), .A2(G138), .ZN(n690) );
  NAND2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n694) );
  NAND2_X1 U776 ( .A1(G102), .A2(n890), .ZN(n692) );
  XNOR2_X1 U777 ( .A(KEYINPUT89), .B(n692), .ZN(n693) );
  NOR2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n917) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n785) );
  NOR2_X1 U780 ( .A1(G1384), .A2(G164), .ZN(n783) );
  INV_X1 U781 ( .A(KEYINPUT64), .ZN(n782) );
  XNOR2_X1 U782 ( .A(n783), .B(n782), .ZN(n695) );
  NOR2_X2 U783 ( .A1(n785), .A2(n695), .ZN(n732) );
  NAND2_X1 U784 ( .A1(n732), .A2(G2072), .ZN(n697) );
  INV_X1 U785 ( .A(KEYINPUT27), .ZN(n696) );
  XNOR2_X1 U786 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U788 ( .A(KEYINPUT98), .B(n700), .Z(n703) );
  NOR2_X1 U789 ( .A1(n703), .A2(n914), .ZN(n702) );
  INV_X1 U790 ( .A(KEYINPUT28), .ZN(n701) );
  XNOR2_X1 U791 ( .A(n702), .B(n701), .ZN(n725) );
  NAND2_X1 U792 ( .A1(n914), .A2(n703), .ZN(n723) );
  AND2_X1 U793 ( .A1(n516), .A2(G1348), .ZN(n705) );
  NAND2_X1 U794 ( .A1(KEYINPUT100), .A2(n705), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n704), .A2(KEYINPUT99), .ZN(n712) );
  INV_X1 U796 ( .A(n705), .ZN(n708) );
  NAND2_X1 U797 ( .A1(G2067), .A2(n732), .ZN(n706) );
  XNOR2_X1 U798 ( .A(KEYINPUT100), .B(n706), .ZN(n707) );
  NAND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n710) );
  INV_X1 U800 ( .A(KEYINPUT99), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n719) );
  OR2_X1 U803 ( .A1(n904), .A2(n719), .ZN(n718) );
  INV_X1 U804 ( .A(G1996), .ZN(n972) );
  OR2_X1 U805 ( .A1(n516), .A2(n972), .ZN(n713) );
  XNOR2_X1 U806 ( .A(n713), .B(KEYINPUT26), .ZN(n715) );
  NAND2_X1 U807 ( .A1(n516), .A2(G1341), .ZN(n714) );
  NAND2_X1 U808 ( .A1(n715), .A2(n714), .ZN(n716) );
  OR2_X1 U809 ( .A1(n930), .A2(n716), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U811 ( .A1(n904), .A2(n719), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U815 ( .A(n726), .B(KEYINPUT29), .Z(n731) );
  XNOR2_X1 U816 ( .A(KEYINPUT25), .B(G2078), .ZN(n971) );
  NOR2_X1 U817 ( .A1(n516), .A2(n971), .ZN(n728) );
  INV_X1 U818 ( .A(G1961), .ZN(n942) );
  NOR2_X1 U819 ( .A1(n732), .A2(n942), .ZN(n727) );
  NOR2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n736) );
  AND2_X1 U821 ( .A1(G171), .A2(n736), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n729), .B(KEYINPUT97), .ZN(n730) );
  NAND2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n742) );
  NAND2_X2 U824 ( .A1(G8), .A2(n516), .ZN(n778) );
  NOR2_X1 U825 ( .A1(G1966), .A2(n778), .ZN(n756) );
  NOR2_X1 U826 ( .A1(G2084), .A2(n516), .ZN(n754) );
  NOR2_X1 U827 ( .A1(n756), .A2(n754), .ZN(n733) );
  NAND2_X1 U828 ( .A1(G8), .A2(n733), .ZN(n734) );
  XNOR2_X1 U829 ( .A(KEYINPUT30), .B(n734), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n735), .A2(G168), .ZN(n738) );
  NOR2_X1 U831 ( .A1(G171), .A2(n736), .ZN(n737) );
  NOR2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U833 ( .A(n739), .B(KEYINPUT101), .ZN(n740) );
  XNOR2_X1 U834 ( .A(n740), .B(KEYINPUT31), .ZN(n741) );
  NAND2_X1 U835 ( .A1(n742), .A2(n741), .ZN(n753) );
  NAND2_X1 U836 ( .A1(n753), .A2(G286), .ZN(n747) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n778), .ZN(n744) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n516), .ZN(n743) );
  NOR2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U840 ( .A1(n745), .A2(G303), .ZN(n746) );
  NAND2_X1 U841 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U842 ( .A(n749), .B(n748), .ZN(n750) );
  NAND2_X1 U843 ( .A1(G8), .A2(n750), .ZN(n752) );
  XNOR2_X1 U844 ( .A(n752), .B(n751), .ZN(n760) );
  NAND2_X1 U845 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U846 ( .A1(n753), .A2(n755), .ZN(n757) );
  NOR2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U848 ( .A(n758), .B(KEYINPUT102), .ZN(n759) );
  NOR2_X2 U849 ( .A1(n760), .A2(n759), .ZN(n771) );
  NOR2_X1 U850 ( .A1(n917), .A2(n771), .ZN(n763) );
  NOR2_X1 U851 ( .A1(G303), .A2(G1971), .ZN(n761) );
  XOR2_X1 U852 ( .A(KEYINPUT104), .B(n761), .Z(n762) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n923) );
  NAND2_X1 U855 ( .A1(n764), .A2(n923), .ZN(n765) );
  NOR2_X1 U856 ( .A1(n765), .A2(n778), .ZN(n766) );
  NOR2_X1 U857 ( .A1(KEYINPUT33), .A2(n766), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n917), .A2(KEYINPUT33), .ZN(n767) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n935) );
  INV_X1 U860 ( .A(n770), .ZN(n781) );
  INV_X1 U861 ( .A(n771), .ZN(n774) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n775), .A2(n778), .ZN(n780) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U867 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  OR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n781), .A2(n518), .ZN(n820) );
  XNOR2_X1 U870 ( .A(G1986), .B(G290), .ZN(n916) );
  XOR2_X1 U871 ( .A(n783), .B(n782), .Z(n784) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n830) );
  NAND2_X1 U873 ( .A1(n916), .A2(n830), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(KEYINPUT90), .ZN(n798) );
  NAND2_X1 U875 ( .A1(G104), .A2(n890), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G140), .A2(n893), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n789), .ZN(n795) );
  NAND2_X1 U879 ( .A1(n885), .A2(G128), .ZN(n790) );
  XOR2_X1 U880 ( .A(KEYINPUT91), .B(n790), .Z(n792) );
  NAND2_X1 U881 ( .A1(n886), .A2(G116), .ZN(n791) );
  NAND2_X1 U882 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U883 ( .A(n793), .B(KEYINPUT35), .Z(n794) );
  NOR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U885 ( .A(KEYINPUT36), .B(n796), .Z(n797) );
  XOR2_X1 U886 ( .A(KEYINPUT92), .B(n797), .Z(n900) );
  XNOR2_X1 U887 ( .A(G2067), .B(KEYINPUT37), .ZN(n827) );
  NOR2_X1 U888 ( .A1(n900), .A2(n827), .ZN(n999) );
  NAND2_X1 U889 ( .A1(n830), .A2(n999), .ZN(n825) );
  NAND2_X1 U890 ( .A1(n798), .A2(n825), .ZN(n818) );
  NAND2_X1 U891 ( .A1(G119), .A2(n885), .ZN(n800) );
  NAND2_X1 U892 ( .A1(G131), .A2(n893), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G107), .A2(n886), .ZN(n801) );
  XNOR2_X1 U895 ( .A(KEYINPUT93), .B(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n890), .A2(G95), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n879) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n879), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n806), .B(KEYINPUT94), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G129), .A2(n885), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G117), .A2(n886), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n890), .A2(G105), .ZN(n809) );
  XOR2_X1 U905 ( .A(KEYINPUT38), .B(n809), .Z(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U907 ( .A(KEYINPUT95), .B(n812), .Z(n814) );
  NAND2_X1 U908 ( .A1(G141), .A2(n893), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n878) );
  NAND2_X1 U910 ( .A1(G1996), .A2(n878), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT96), .B(n817), .ZN(n1003) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n832) );
  NOR2_X1 U914 ( .A1(G1996), .A2(n878), .ZN(n994) );
  NOR2_X1 U915 ( .A1(G1986), .A2(G290), .ZN(n821) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n879), .ZN(n997) );
  NOR2_X1 U917 ( .A1(n821), .A2(n997), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n520), .A2(n822), .ZN(n823) );
  NOR2_X1 U919 ( .A1(n994), .A2(n823), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n824), .B(KEYINPUT39), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n900), .A2(n827), .ZN(n1008) );
  NAND2_X1 U923 ( .A1(n828), .A2(n1008), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U926 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  XNOR2_X1 U931 ( .A(KEYINPUT108), .B(n836), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U939 ( .A(KEYINPUT109), .B(n841), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2474), .B(G1956), .Z(n843) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n844), .B(KEYINPUT112), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1971), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(G1976), .B(G1981), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1961), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U950 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(G229) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n854) );
  XNOR2_X1 U953 ( .A(G2090), .B(KEYINPUT42), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U955 ( .A(n855), .B(G2678), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U958 ( .A(KEYINPUT110), .B(G2100), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U962 ( .A1(G124), .A2(n885), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n862), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n893), .A2(G136), .ZN(n863) );
  XOR2_X1 U965 ( .A(KEYINPUT113), .B(n863), .Z(n864) );
  NAND2_X1 U966 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G100), .A2(n890), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G112), .A2(n886), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U970 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G130), .A2(n885), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G118), .A2(n886), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G106), .A2(n890), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G142), .A2(n893), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U977 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT114), .B(n875), .ZN(n876) );
  NOR2_X1 U979 ( .A1(n877), .A2(n876), .ZN(n882) );
  XNOR2_X1 U980 ( .A(G160), .B(n878), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U982 ( .A(n882), .B(n881), .Z(n884) );
  XNOR2_X1 U983 ( .A(G164), .B(G162), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n902) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n898) );
  NAND2_X1 U986 ( .A1(G127), .A2(n885), .ZN(n888) );
  NAND2_X1 U987 ( .A1(G115), .A2(n886), .ZN(n887) );
  NAND2_X1 U988 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n889), .B(KEYINPUT47), .ZN(n892) );
  NAND2_X1 U990 ( .A1(G103), .A2(n890), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n896) );
  NAND2_X1 U992 ( .A1(G139), .A2(n893), .ZN(n894) );
  XNOR2_X1 U993 ( .A(KEYINPUT115), .B(n894), .ZN(n895) );
  NOR2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n988) );
  XNOR2_X1 U995 ( .A(n996), .B(n988), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U999 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(G171), .B(n904), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n905), .B(G286), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n908), .ZN(G397) );
  NOR2_X1 U1004 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n910), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n911) );
  AND2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n913), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G303), .ZN(G166) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1013 ( .A(G16), .B(KEYINPUT56), .ZN(n941) );
  XNOR2_X1 U1014 ( .A(n914), .B(G1956), .ZN(n915) );
  XNOR2_X1 U1015 ( .A(n915), .B(KEYINPUT122), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n922) );
  XOR2_X1 U1018 ( .A(G1971), .B(G303), .Z(n920) );
  XNOR2_X1 U1019 ( .A(KEYINPUT123), .B(n920), .ZN(n921) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n924) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n934) );
  XNOR2_X1 U1022 ( .A(n925), .B(G1348), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(G171), .B(G1961), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT121), .B(n928), .ZN(n932) );
  XOR2_X1 U1026 ( .A(G1341), .B(KEYINPUT124), .Z(n929) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n931) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n939) );
  XNOR2_X1 U1030 ( .A(G1966), .B(G168), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(n937), .B(KEYINPUT57), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n1020) );
  XNOR2_X1 U1035 ( .A(G5), .B(n942), .ZN(n956) );
  XNOR2_X1 U1036 ( .A(KEYINPUT59), .B(G1348), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n943), .B(G4), .ZN(n948) );
  XOR2_X1 U1038 ( .A(G1956), .B(KEYINPUT125), .Z(n944) );
  XNOR2_X1 U1039 ( .A(G20), .B(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(G6), .B(G1981), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(KEYINPUT126), .B(G1341), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(G19), .B(n949), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1046 ( .A(KEYINPUT60), .B(n952), .Z(n954) );
  XNOR2_X1 U1047 ( .A(G1966), .B(G21), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n963) );
  XNOR2_X1 U1050 ( .A(G1986), .B(G24), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G1971), .B(G22), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n960) );
  XOR2_X1 U1053 ( .A(G1976), .B(G23), .Z(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT58), .B(n961), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT61), .B(n964), .Z(n965) );
  NOR2_X1 U1058 ( .A1(G16), .A2(n965), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT127), .B(n966), .ZN(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(G11), .ZN(n1018) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G26), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(G33), .B(G2072), .ZN(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n978) );
  XOR2_X1 U1064 ( .A(G1991), .B(G25), .Z(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(G28), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(n971), .B(G27), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n972), .B(G32), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n979), .B(KEYINPUT53), .ZN(n982) );
  XOR2_X1 U1072 ( .A(G2084), .B(KEYINPUT54), .Z(n980) );
  XNOR2_X1 U1073 ( .A(G34), .B(n980), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(G35), .B(G2090), .ZN(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1077 ( .A(KEYINPUT120), .B(n985), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(G29), .A2(n986), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(n987), .B(KEYINPUT55), .ZN(n1016) );
  XNOR2_X1 U1080 ( .A(G2072), .B(n988), .ZN(n989) );
  XNOR2_X1 U1081 ( .A(n989), .B(KEYINPUT119), .ZN(n991) );
  XOR2_X1 U1082 ( .A(G2078), .B(G164), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT50), .B(n992), .ZN(n1012) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n995), .Z(n1006) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(G160), .B(G2084), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT116), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT117), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT118), .B(n1010), .Z(n1011) );
  NAND2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(KEYINPUT52), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1100 ( .A1(G29), .A2(n1014), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1104 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1105 ( .A(G311), .ZN(G150) );
endmodule

