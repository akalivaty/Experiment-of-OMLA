

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XNOR2_X1 U323 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U324 ( .A(n433), .B(KEYINPUT119), .ZN(n434) );
  XOR2_X1 U325 ( .A(KEYINPUT28), .B(n467), .Z(n536) );
  XOR2_X1 U326 ( .A(G120GAT), .B(G106GAT), .Z(n291) );
  INV_X1 U327 ( .A(KEYINPUT54), .ZN(n433) );
  XNOR2_X1 U328 ( .A(n405), .B(n291), .ZN(n392) );
  XNOR2_X1 U329 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n430) );
  XNOR2_X1 U330 ( .A(n393), .B(n392), .ZN(n397) );
  XNOR2_X1 U331 ( .A(n431), .B(n430), .ZN(n531) );
  XOR2_X1 U332 ( .A(KEYINPUT89), .B(n475), .Z(n520) );
  XNOR2_X1 U333 ( .A(n457), .B(G190GAT), .ZN(n458) );
  XNOR2_X1 U334 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U335 ( .A(G36GAT), .B(G190GAT), .Z(n352) );
  XOR2_X1 U336 ( .A(G99GAT), .B(G85GAT), .Z(n398) );
  XOR2_X1 U337 ( .A(n352), .B(n398), .Z(n293) );
  XOR2_X1 U338 ( .A(G50GAT), .B(G106GAT), .Z(n438) );
  XOR2_X1 U339 ( .A(G29GAT), .B(G134GAT), .Z(n330) );
  XNOR2_X1 U340 ( .A(n438), .B(n330), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n299) );
  INV_X1 U342 ( .A(G92GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n295), .B(KEYINPUT7), .ZN(n381) );
  XOR2_X1 U345 ( .A(G92GAT), .B(n381), .Z(n297) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U348 ( .A(n299), .B(n298), .Z(n307) );
  XOR2_X1 U349 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n301) );
  XNOR2_X1 U350 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U352 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n303) );
  XNOR2_X1 U353 ( .A(G162GAT), .B(KEYINPUT11), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n559) );
  INV_X1 U357 ( .A(KEYINPUT120), .ZN(n456) );
  XOR2_X1 U358 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n309) );
  XNOR2_X1 U359 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U361 ( .A(n310), .B(KEYINPUT82), .Z(n312) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(KEYINPUT83), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n362) );
  XOR2_X1 U364 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n314) );
  XNOR2_X1 U365 ( .A(G15GAT), .B(G183GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n362), .B(n315), .ZN(n328) );
  XOR2_X1 U368 ( .A(G99GAT), .B(G134GAT), .Z(n317) );
  XNOR2_X1 U369 ( .A(G43GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n326) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n318), .B(G120GAT), .ZN(n333) );
  XOR2_X1 U373 ( .A(G71GAT), .B(n333), .Z(n320) );
  NAND2_X1 U374 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U376 ( .A(G127GAT), .B(G176GAT), .Z(n322) );
  XNOR2_X1 U377 ( .A(KEYINPUT81), .B(KEYINPUT20), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U379 ( .A(n324), .B(n323), .Z(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n533) );
  INV_X1 U382 ( .A(KEYINPUT55), .ZN(n453) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(G127GAT), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n329), .B(G57GAT), .ZN(n413) );
  XOR2_X1 U385 ( .A(n413), .B(G85GAT), .Z(n332) );
  XNOR2_X1 U386 ( .A(G148GAT), .B(n330), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n337) );
  XOR2_X1 U388 ( .A(n333), .B(KEYINPUT5), .Z(n335) );
  NAND2_X1 U389 ( .A1(G225GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U391 ( .A(n337), .B(n336), .Z(n346) );
  XNOR2_X1 U392 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n338), .B(KEYINPUT3), .ZN(n339) );
  XOR2_X1 U394 ( .A(n339), .B(KEYINPUT86), .Z(n341) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(G162GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n451) );
  XOR2_X1 U397 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n343) );
  XNOR2_X1 U398 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n451), .B(n344), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n475) );
  NAND2_X1 U402 ( .A1(G64GAT), .A2(n294), .ZN(n349) );
  INV_X1 U403 ( .A(G64GAT), .ZN(n347) );
  NAND2_X1 U404 ( .A1(n347), .A2(G92GAT), .ZN(n348) );
  NAND2_X1 U405 ( .A1(n349), .A2(n348), .ZN(n351) );
  XNOR2_X1 U406 ( .A(G176GAT), .B(G204GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n389) );
  XOR2_X1 U408 ( .A(n352), .B(n389), .Z(n354) );
  NAND2_X1 U409 ( .A1(G226GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n366) );
  XOR2_X1 U411 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n356) );
  XNOR2_X1 U412 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n359) );
  XOR2_X1 U414 ( .A(KEYINPUT75), .B(G211GAT), .Z(n358) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(G183GAT), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n412) );
  XOR2_X1 U417 ( .A(n359), .B(n412), .Z(n364) );
  XOR2_X1 U418 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n361) );
  XNOR2_X1 U419 ( .A(G197GAT), .B(G218GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n361), .B(n360), .ZN(n437) );
  XNOR2_X1 U421 ( .A(n362), .B(n437), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n522) );
  XNOR2_X1 U424 ( .A(n522), .B(KEYINPUT118), .ZN(n432) );
  XOR2_X1 U425 ( .A(G141GAT), .B(G113GAT), .Z(n368) );
  XNOR2_X1 U426 ( .A(G169GAT), .B(G29GAT), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U428 ( .A(KEYINPUT67), .B(G8GAT), .Z(n370) );
  XNOR2_X1 U429 ( .A(G197GAT), .B(G1GAT), .ZN(n369) );
  XNOR2_X1 U430 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U431 ( .A(n372), .B(n371), .Z(n379) );
  INV_X1 U432 ( .A(G50GAT), .ZN(n374) );
  XNOR2_X1 U433 ( .A(G15GAT), .B(G22GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n373), .B(KEYINPUT69), .ZN(n404) );
  XNOR2_X1 U435 ( .A(n374), .B(n404), .ZN(n376) );
  NAND2_X1 U436 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U438 ( .A(G36GAT), .B(n377), .ZN(n378) );
  XNOR2_X1 U439 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n380), .B(KEYINPUT30), .ZN(n383) );
  XOR2_X1 U441 ( .A(n381), .B(KEYINPUT29), .Z(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U443 ( .A(KEYINPUT65), .B(KEYINPUT70), .Z(n385) );
  XNOR2_X1 U444 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X2 U446 ( .A(n387), .B(n386), .ZN(n575) );
  INV_X1 U447 ( .A(KEYINPUT32), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n391) );
  NAND2_X1 U449 ( .A1(G230GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n393) );
  XOR2_X1 U451 ( .A(G71GAT), .B(KEYINPUT13), .Z(n405) );
  XOR2_X1 U452 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n395) );
  XNOR2_X1 U453 ( .A(G57GAT), .B(KEYINPUT31), .ZN(n394) );
  XOR2_X1 U454 ( .A(n395), .B(n394), .Z(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n400) );
  XOR2_X1 U456 ( .A(G148GAT), .B(G78GAT), .Z(n439) );
  XNOR2_X1 U457 ( .A(n439), .B(n398), .ZN(n399) );
  XNOR2_X1 U458 ( .A(n400), .B(n399), .ZN(n579) );
  XNOR2_X1 U459 ( .A(n579), .B(KEYINPUT41), .ZN(n564) );
  NAND2_X1 U460 ( .A1(n575), .A2(n564), .ZN(n401) );
  XNOR2_X1 U461 ( .A(KEYINPUT46), .B(n401), .ZN(n420) );
  XOR2_X1 U462 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n403) );
  XNOR2_X1 U463 ( .A(G155GAT), .B(G78GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n417) );
  XOR2_X1 U465 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U466 ( .A1(G231GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U468 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n409) );
  XNOR2_X1 U469 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U471 ( .A(n411), .B(n410), .Z(n415) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U474 ( .A(n417), .B(n416), .Z(n493) );
  INV_X1 U475 ( .A(n493), .ZN(n582) );
  XNOR2_X1 U476 ( .A(KEYINPUT109), .B(n582), .ZN(n570) );
  INV_X1 U477 ( .A(n559), .ZN(n418) );
  AND2_X1 U478 ( .A1(n570), .A2(n418), .ZN(n419) );
  AND2_X1 U479 ( .A1(n420), .A2(n419), .ZN(n422) );
  XNOR2_X1 U480 ( .A(KEYINPUT47), .B(KEYINPUT110), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n429) );
  INV_X1 U482 ( .A(KEYINPUT36), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n559), .B(KEYINPUT102), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n590) );
  NOR2_X1 U485 ( .A1(n493), .A2(n590), .ZN(n425) );
  XOR2_X1 U486 ( .A(KEYINPUT45), .B(n425), .Z(n426) );
  NOR2_X1 U487 ( .A1(n575), .A2(n426), .ZN(n427) );
  NAND2_X1 U488 ( .A1(n427), .A2(n579), .ZN(n428) );
  NAND2_X1 U489 ( .A1(n429), .A2(n428), .ZN(n431) );
  NAND2_X1 U490 ( .A1(n432), .A2(n531), .ZN(n435) );
  NOR2_X1 U491 ( .A1(n520), .A2(n436), .ZN(n574) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U494 ( .A(G204GAT), .B(KEYINPUT22), .Z(n442) );
  NAND2_X1 U495 ( .A1(G228GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n449) );
  XOR2_X1 U498 ( .A(G211GAT), .B(KEYINPUT24), .Z(n446) );
  XNOR2_X1 U499 ( .A(KEYINPUT23), .B(KEYINPUT87), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(G22GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n467) );
  NAND2_X1 U504 ( .A1(n574), .A2(n467), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n454) );
  NOR2_X1 U506 ( .A1(n533), .A2(n454), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n569) );
  INV_X1 U508 ( .A(n569), .ZN(n563) );
  NAND2_X1 U509 ( .A1(n559), .A2(n563), .ZN(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT99), .Z(n482) );
  NAND2_X1 U512 ( .A1(n579), .A2(n575), .ZN(n495) );
  XNOR2_X1 U513 ( .A(KEYINPUT78), .B(KEYINPUT16), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n559), .A2(n493), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n461), .B(n460), .ZN(n480) );
  XNOR2_X1 U516 ( .A(KEYINPUT27), .B(n522), .ZN(n470) );
  NAND2_X1 U517 ( .A1(n520), .A2(n470), .ZN(n530) );
  INV_X1 U518 ( .A(n533), .ZN(n524) );
  OR2_X1 U519 ( .A1(n536), .A2(n524), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n530), .A2(n462), .ZN(n478) );
  NAND2_X1 U521 ( .A1(n522), .A2(n524), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n463), .A2(n467), .ZN(n464) );
  XNOR2_X1 U523 ( .A(n464), .B(KEYINPUT25), .ZN(n466) );
  XOR2_X1 U524 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n465) );
  XNOR2_X1 U525 ( .A(n466), .B(n465), .ZN(n473) );
  NOR2_X1 U526 ( .A1(n524), .A2(n467), .ZN(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n573) );
  NAND2_X1 U529 ( .A1(n470), .A2(n573), .ZN(n471) );
  XNOR2_X1 U530 ( .A(KEYINPUT95), .B(n471), .ZN(n472) );
  NOR2_X1 U531 ( .A1(n473), .A2(n472), .ZN(n474) );
  NOR2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n476), .B(KEYINPUT98), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n491) );
  INV_X1 U535 ( .A(n491), .ZN(n479) );
  NAND2_X1 U536 ( .A1(n480), .A2(n479), .ZN(n507) );
  NOR2_X1 U537 ( .A1(n495), .A2(n507), .ZN(n489) );
  NAND2_X1 U538 ( .A1(n489), .A2(n520), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U541 ( .A1(n522), .A2(n489), .ZN(n484) );
  XNOR2_X1 U542 ( .A(n484), .B(KEYINPUT100), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G8GAT), .B(n485), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n487) );
  NAND2_X1 U545 ( .A1(n489), .A2(n524), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U547 ( .A(G15GAT), .B(n488), .Z(G1326GAT) );
  NAND2_X1 U548 ( .A1(n536), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n490), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  NOR2_X1 U551 ( .A1(n491), .A2(n590), .ZN(n492) );
  NAND2_X1 U552 ( .A1(n493), .A2(n492), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT37), .B(n494), .Z(n519) );
  NOR2_X1 U554 ( .A1(n519), .A2(n495), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT38), .B(n496), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n520), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n522), .A2(n504), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n504), .A2(n524), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n504), .A2(n536), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n509) );
  INV_X1 U568 ( .A(n575), .ZN(n506) );
  NAND2_X1 U569 ( .A1(n506), .A2(n564), .ZN(n518) );
  NOR2_X1 U570 ( .A1(n518), .A2(n507), .ZN(n514) );
  NAND2_X1 U571 ( .A1(n514), .A2(n520), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n522), .A2(n514), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n524), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(KEYINPUT106), .ZN(n513) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U580 ( .A1(n514), .A2(n536), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n520), .A2(n526), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n522), .A2(n526), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n526), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n528) );
  NAND2_X1 U591 ( .A1(n526), .A2(n536), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U593 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  INV_X1 U594 ( .A(n530), .ZN(n532) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n549) );
  NOR2_X1 U596 ( .A1(n533), .A2(n549), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(KEYINPUT111), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n575), .A2(n545), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U602 ( .A1(n545), .A2(n564), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  INV_X1 U605 ( .A(n545), .ZN(n541) );
  NOR2_X1 U606 ( .A1(n570), .A2(n541), .ZN(n543) );
  XNOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n559), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n548), .ZN(G1343GAT) );
  XOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT115), .Z(n552) );
  INV_X1 U615 ( .A(n573), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n560), .A2(n575), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U621 ( .A1(n560), .A2(n564), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT117), .Z(n558) );
  NAND2_X1 U625 ( .A1(n560), .A2(n582), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n575), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(n571), .Z(n572) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(n572), .ZN(G1350GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n589) );
  INV_X1 U640 ( .A(n589), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n575), .A2(n583), .ZN(n578) );
  XOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT60), .Z(n576) );
  XNOR2_X1 U643 ( .A(KEYINPUT59), .B(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  OR2_X1 U646 ( .A1(n589), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n585) );
  NAND2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n592) );
  NOR2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U656 ( .A(n592), .B(n591), .Z(G1355GAT) );
endmodule

