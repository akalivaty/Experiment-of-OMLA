//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n541, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n462), .A2(new_n464), .A3(G137), .A4(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n461), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n467), .B1(new_n466), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n462), .A2(new_n464), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n472), .B1(G2105), .B2(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n474), .A2(new_n465), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n462), .A2(new_n464), .A3(G138), .A4(new_n465), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G138), .A4(new_n465), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT5), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G62), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT68), .B(G651), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT6), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(G543), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(new_n502), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n508), .A2(new_n514), .A3(new_n510), .ZN(new_n515));
  OAI221_X1 g090(.A(new_n507), .B1(new_n511), .B2(new_n512), .C1(new_n513), .C2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  INV_X1    g092(.A(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G89), .ZN(new_n519));
  INV_X1    g094(.A(new_n511), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT69), .B(G51), .Z(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n519), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  AOI22_X1  g102(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n505), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n518), .A2(G90), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n520), .A2(G52), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  AOI22_X1  g108(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n505), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n518), .A2(G81), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n520), .A2(G43), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G188));
  NAND3_X1  g120(.A1(new_n520), .A2(KEYINPUT9), .A3(G53), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(G91), .ZN(new_n547));
  INV_X1    g122(.A(G78), .ZN(new_n548));
  OR3_X1    g123(.A1(new_n548), .A2(new_n498), .A3(KEYINPUT70), .ZN(new_n549));
  OAI21_X1  g124(.A(KEYINPUT70), .B1(new_n548), .B2(new_n498), .ZN(new_n550));
  INV_X1    g125(.A(G65), .ZN(new_n551));
  OAI211_X1 g126(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n502), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n511), .B2(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n546), .A2(new_n547), .A3(new_n553), .A4(new_n556), .ZN(G299));
  OAI21_X1  g132(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n558));
  INV_X1    g133(.A(G49), .ZN(new_n559));
  INV_X1    g134(.A(G87), .ZN(new_n560));
  OAI221_X1 g135(.A(new_n558), .B1(new_n511), .B2(new_n559), .C1(new_n560), .C2(new_n515), .ZN(G288));
  NAND4_X1  g136(.A1(new_n508), .A2(new_n514), .A3(G86), .A4(new_n510), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT71), .ZN(new_n565));
  INV_X1    g140(.A(G61), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n502), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n499), .A2(new_n501), .A3(KEYINPUT71), .A4(G61), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(new_n506), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n564), .B1(new_n571), .B2(KEYINPUT72), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n520), .A2(G48), .B1(new_n562), .B2(new_n563), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n575), .A3(new_n506), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n505), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n520), .A2(G47), .ZN(new_n580));
  XNOR2_X1  g155(.A(KEYINPUT74), .B(G85), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n518), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT75), .B(KEYINPUT10), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n515), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G651), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n520), .A2(G54), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n586), .B1(new_n515), .B2(new_n585), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n587), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n584), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n584), .B1(new_n594), .B2(G868), .ZN(G321));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  XOR2_X1   g172(.A(G299), .B(KEYINPUT76), .Z(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G297));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(G868), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n538), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n593), .A2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n493), .A2(new_n468), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT77), .B(KEYINPUT12), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT78), .B(G2100), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n478), .ZN(new_n614));
  INV_X1    g189(.A(G123), .ZN(new_n615));
  OR3_X1    g190(.A1(new_n614), .A2(KEYINPUT79), .A3(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(KEYINPUT79), .B1(new_n614), .B2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n480), .A2(G135), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n465), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n616), .A2(new_n617), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2096), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT80), .ZN(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  INV_X1    g200(.A(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  OAI21_X1  g203(.A(KEYINPUT14), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT82), .Z(new_n630));
  NAND2_X1  g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT83), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n636), .B(new_n638), .Z(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n636), .B(new_n638), .ZN(new_n642));
  INV_X1    g217(.A(new_n640), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n644), .A3(G14), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n647), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2100), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n649), .A2(new_n650), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n654), .B(new_n657), .Z(G227));
  XNOR2_X1  g233(.A(G1971), .B(G1976), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT20), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n666), .B1(new_n660), .B2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n665), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT85), .B(G1981), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1986), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n676), .B(new_n678), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  INV_X1    g255(.A(KEYINPUT95), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G24), .ZN(new_n683));
  INV_X1    g258(.A(G290), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1986), .ZN(new_n686));
  AND2_X1   g261(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n478), .A2(G119), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n480), .A2(G131), .ZN(new_n689));
  OAI21_X1  g264(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n465), .A2(G107), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n688), .B(new_n689), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  MUX2_X1   g267(.A(G25), .B(new_n692), .S(G29), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT35), .B(G1991), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n686), .A2(new_n687), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G16), .A2(G22), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G166), .B2(G16), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT87), .B(G1971), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n682), .A2(G23), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n558), .B1(new_n515), .B2(new_n560), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G49), .B2(new_n520), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n702), .B1(new_n704), .B2(new_n682), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT33), .B(G1976), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n574), .A2(G16), .A3(new_n576), .ZN(new_n709));
  OR2_X1    g284(.A1(G6), .A2(G16), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT32), .B(G1981), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n710), .ZN(new_n713));
  INV_X1    g288(.A(new_n711), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n708), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n708), .A2(new_n717), .A3(new_n712), .A4(new_n715), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n697), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n725), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g303(.A1(G160), .A2(G29), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT24), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n725), .B1(new_n730), .B2(G34), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n730), .A2(G34), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n732), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n728), .A2(G2090), .B1(G2084), .B2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n728), .ZN(new_n739));
  INV_X1    g314(.A(G2090), .ZN(new_n740));
  OAI21_X1  g315(.A(KEYINPUT94), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n728), .A2(new_n742), .A3(G2090), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n738), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n480), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n478), .A2(G129), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n468), .A2(G105), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT26), .Z(new_n749));
  NAND4_X1  g324(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(new_n725), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G32), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n751), .A2(KEYINPUT93), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(KEYINPUT93), .B2(new_n751), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT27), .B(G1996), .Z(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n758));
  OAI22_X1  g333(.A1(new_n621), .A2(new_n725), .B1(new_n758), .B2(G11), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n754), .A2(new_n756), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n737), .A2(G2084), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(G28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(G28), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n764), .A2(new_n765), .A3(new_n725), .ZN(new_n766));
  AND4_X1   g341(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n766), .ZN(new_n767));
  AND3_X1   g342(.A1(new_n744), .A2(new_n757), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n539), .A2(new_n682), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n682), .B2(G19), .ZN(new_n770));
  INV_X1    g345(.A(G1341), .ZN(new_n771));
  NAND2_X1  g346(.A1(G168), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G16), .B2(G21), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  OAI22_X1  g349(.A1(new_n770), .A2(new_n771), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n682), .A2(KEYINPUT23), .A3(G20), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT23), .ZN(new_n777));
  INV_X1    g352(.A(G20), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G16), .ZN(new_n779));
  INV_X1    g354(.A(G299), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n776), .B(new_n779), .C1(new_n780), .C2(new_n682), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1956), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n775), .B(new_n782), .C1(new_n771), .C2(new_n770), .ZN(new_n783));
  NOR2_X1   g358(.A1(G27), .A2(G29), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G164), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G2078), .Z(new_n786));
  NAND2_X1  g361(.A1(G171), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G5), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(G1961), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n682), .A2(G4), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n594), .B2(new_n682), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1348), .ZN(new_n793));
  AOI211_X1 g368(.A(new_n790), .B(new_n793), .C1(new_n774), .C2(new_n773), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n768), .A2(new_n783), .A3(new_n786), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n724), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n725), .A2(G26), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n478), .A2(G128), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT89), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n480), .A2(G140), .ZN(new_n800));
  OR2_X1    g375(.A1(G104), .A2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n801), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n797), .B1(new_n805), .B2(new_n725), .ZN(new_n806));
  MUX2_X1   g381(.A(new_n797), .B(new_n806), .S(KEYINPUT28), .Z(new_n807));
  INV_X1    g382(.A(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n788), .A2(new_n789), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n721), .A2(new_n723), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n796), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n468), .A2(G103), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT25), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n480), .A2(G139), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n814), .A2(KEYINPUT90), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(KEYINPUT90), .B1(new_n814), .B2(new_n815), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n818));
  OAI22_X1  g393(.A1(new_n816), .A2(new_n817), .B1(new_n465), .B2(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G33), .B(new_n819), .S(G29), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT91), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G2072), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n681), .B1(new_n812), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n811), .ZN(new_n824));
  INV_X1    g399(.A(new_n810), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n824), .A2(new_n724), .A3(new_n825), .A4(new_n795), .ZN(new_n826));
  INV_X1    g401(.A(new_n822), .ZN(new_n827));
  NAND4_X1  g402(.A1(new_n826), .A2(KEYINPUT95), .A3(new_n827), .A4(new_n809), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(new_n828), .ZN(G311));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n827), .A3(new_n809), .ZN(G150));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n502), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT96), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n506), .ZN(new_n835));
  AOI22_X1  g410(.A1(G55), .A2(new_n520), .B1(new_n518), .B2(G93), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G860), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT97), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n538), .A2(new_n836), .A3(new_n835), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n538), .B1(new_n836), .B2(new_n835), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT39), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n593), .A2(new_n601), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n840), .B1(new_n848), .B2(G860), .ZN(G145));
  NAND2_X1  g424(.A1(new_n480), .A2(G142), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT98), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(KEYINPUT98), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n852), .B(new_n853), .C1(G118), .C2(new_n465), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n478), .A2(G130), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n850), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n750), .B(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT99), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n610), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n692), .B(G164), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G160), .B(G162), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n621), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n819), .B(new_n804), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n861), .A2(new_n865), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n844), .B(new_n605), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n593), .B(G299), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT101), .B1(new_n780), .B2(new_n593), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n594), .A2(G299), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n780), .A2(new_n593), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n878), .B1(new_n881), .B2(KEYINPUT101), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n877), .B1(new_n882), .B2(KEYINPUT41), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n875), .B1(new_n872), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n874), .B1(new_n884), .B2(new_n871), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n704), .B(G303), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(G305), .ZN(new_n889));
  XNOR2_X1  g464(.A(G303), .B(G288), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n576), .A3(new_n574), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n891), .A3(new_n684), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n684), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  OAI211_X1 g470(.A(KEYINPUT42), .B(new_n874), .C1(new_n884), .C2(new_n871), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n887), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n887), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(G868), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n837), .A2(new_n603), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(G295));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n900), .ZN(G331));
  NAND2_X1  g477(.A1(G168), .A2(G301), .ZN(new_n903));
  NAND2_X1  g478(.A1(G171), .A2(G286), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n843), .B2(new_n842), .ZN(new_n906));
  INV_X1    g481(.A(new_n843), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n907), .A2(new_n841), .A3(new_n904), .A4(new_n903), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n906), .A2(new_n881), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n878), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n873), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n913), .A2(new_n914), .B1(new_n873), .B2(new_n876), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n906), .A2(new_n908), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n910), .B(new_n894), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n906), .A2(new_n908), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n909), .B1(new_n883), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(KEYINPUT104), .A3(new_n894), .ZN(new_n922));
  INV_X1    g497(.A(new_n894), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n915), .A2(new_n916), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n909), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n919), .A2(new_n867), .A3(new_n922), .A4(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n910), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n873), .A2(new_n876), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n919), .A2(new_n932), .A3(new_n867), .A4(new_n922), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n933), .A2(new_n927), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n928), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n933), .A2(new_n936), .A3(KEYINPUT43), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n919), .A2(new_n867), .A3(new_n922), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n927), .A3(new_n932), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n935), .B1(new_n942), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g518(.A1(new_n492), .A2(new_n495), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n486), .A2(new_n489), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n476), .A2(G2105), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(G40), .C1(new_n470), .C2(new_n471), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n804), .B(G2067), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n750), .B(G1996), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n692), .A2(new_n694), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n692), .A2(new_n694), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1986), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n684), .ZN(new_n961));
  NOR2_X1   g536(.A1(G290), .A2(G1986), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n952), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n944), .A2(new_n945), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI211_X1 g544(.A(KEYINPUT107), .B(G1384), .C1(new_n944), .C2(new_n945), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n951), .B1(new_n947), .B2(KEYINPUT50), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(G164), .B2(G1384), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n967), .A2(new_n966), .A3(new_n968), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n977), .A2(KEYINPUT108), .A3(new_n965), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n974), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT118), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT118), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n973), .A2(new_n981), .A3(new_n974), .A4(new_n978), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n789), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n975), .A2(new_n976), .A3(new_n948), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n951), .B1(KEYINPUT45), .B2(new_n946), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(G2078), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n949), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n986), .B1(new_n989), .B2(G2078), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n983), .A2(new_n988), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n993), .A2(G171), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n951), .B(KEYINPUT126), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n946), .A2(KEYINPUT45), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n949), .A3(new_n996), .A4(new_n987), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n983), .A2(new_n991), .A3(new_n992), .A4(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G171), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n964), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  INV_X1    g576(.A(G8), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n984), .A2(new_n985), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT112), .B1(new_n1003), .B2(new_n774), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n1006));
  AOI211_X1 g581(.A(new_n1006), .B(G1966), .C1(new_n984), .C2(new_n985), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G2084), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n973), .A2(new_n1010), .A3(new_n974), .A4(new_n978), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1002), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G286), .A2(G8), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT123), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT124), .B(new_n1001), .C1(new_n1012), .C2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1011), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1016), .B2(G8), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT124), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1014), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n951), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n977), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n704), .A2(G1976), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1026), .A2(KEYINPUT109), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G288), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1002), .B1(new_n977), .B2(new_n1022), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1981), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n572), .A2(new_n1035), .A3(new_n576), .A4(new_n573), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n520), .A2(G48), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(new_n571), .A3(new_n562), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(G1981), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(KEYINPUT110), .A2(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1036), .B(new_n1039), .C1(KEYINPUT110), .C2(KEYINPUT49), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1032), .A3(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1034), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n973), .A2(new_n740), .A3(new_n974), .A4(new_n978), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT106), .B(G1971), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n989), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G303), .A2(G8), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT55), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(G8), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1022), .A2(new_n965), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1023), .A2(KEYINPUT111), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n946), .A2(new_n965), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT111), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(new_n1022), .C1(new_n977), .C2(new_n965), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(new_n740), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1002), .B1(new_n1059), .B2(new_n1048), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1045), .B(new_n1053), .C1(new_n1052), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n998), .A2(G171), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(KEYINPUT54), .C1(G171), .C2(new_n993), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1000), .A2(new_n1021), .A3(new_n1062), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1055), .A2(new_n1056), .A3(new_n1058), .ZN(new_n1066));
  INV_X1    g641(.A(G1956), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT56), .B(G2072), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n985), .A2(new_n949), .A3(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(new_n1070), .B(KEYINPUT115), .Z(new_n1071));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n1072));
  XNOR2_X1  g647(.A(G299), .B(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1068), .A2(new_n1071), .A3(new_n1076), .A4(new_n1073), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1348), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n980), .A2(new_n1080), .A3(new_n982), .ZN(new_n1081));
  XOR2_X1   g656(.A(new_n1023), .B(KEYINPUT117), .Z(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n808), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n593), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1073), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT119), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  NOR3_X1   g664(.A1(new_n1088), .A2(new_n1078), .A3(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT60), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n594), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1081), .A2(new_n1083), .A3(KEYINPUT60), .A4(new_n593), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1074), .B1(new_n1085), .B2(KEYINPUT122), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1068), .A2(new_n1071), .A3(new_n1102), .A4(new_n1073), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(KEYINPUT61), .A3(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1023), .B(KEYINPUT117), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(G1341), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1996), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n985), .A2(new_n949), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n538), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT59), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1111), .B(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1098), .A2(new_n1100), .A3(new_n1104), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1065), .B1(new_n1091), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1015), .A2(new_n1019), .A3(new_n1118), .A4(new_n1020), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1117), .A2(new_n1062), .A3(new_n994), .A4(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1053), .A2(new_n1044), .A3(new_n1034), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1059), .A2(new_n1048), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1052), .B1(new_n1122), .B2(G8), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1016), .A2(G8), .A3(G168), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT113), .B1(new_n1125), .B2(KEYINPUT63), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1049), .A2(G8), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1051), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1127), .A2(KEYINPUT114), .A3(KEYINPUT63), .A4(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1045), .A2(new_n1012), .A3(G168), .A4(new_n1053), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(KEYINPUT63), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT113), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1135), .B(new_n1136), .C1(new_n1061), .C2(new_n1124), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1126), .A2(new_n1130), .A3(new_n1134), .A4(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1044), .A2(new_n1030), .A3(new_n704), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n1036), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1053), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1140), .A2(new_n1032), .B1(new_n1141), .B2(new_n1045), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1120), .A2(new_n1138), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n963), .B1(new_n1116), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n952), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n955), .A2(new_n958), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n805), .A2(new_n808), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n952), .B1(new_n953), .B2(new_n750), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT46), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1145), .B2(G1996), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n952), .A2(KEYINPUT46), .A3(new_n1109), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1149), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1153), .B(KEYINPUT47), .Z(new_n1154));
  OAI21_X1  g729(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n952), .A2(new_n962), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n1156), .B(KEYINPUT48), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1148), .B(new_n1154), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1144), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g734(.A1(new_n940), .A2(KEYINPUT105), .A3(new_n927), .A4(new_n932), .ZN(new_n1161));
  AOI21_X1  g735(.A(new_n936), .B1(new_n926), .B2(KEYINPUT43), .ZN(new_n1162));
  NOR2_X1   g736(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n1163));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g738(.A(G227), .ZN(new_n1165));
  NAND3_X1  g739(.A1(new_n645), .A2(G319), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n1166), .A2(KEYINPUT127), .ZN(new_n1167));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n645), .A2(new_n1168), .A3(G319), .A4(new_n1165), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  AND2_X1   g744(.A1(new_n869), .A2(new_n679), .ZN(new_n1171));
  AND3_X1   g745(.A1(new_n1164), .A2(new_n1170), .A3(new_n1171), .ZN(G308));
  NAND3_X1  g746(.A1(new_n1164), .A2(new_n1170), .A3(new_n1171), .ZN(G225));
endmodule


