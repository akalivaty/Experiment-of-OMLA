//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n563, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n602, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND3_X1   g037(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(KEYINPUT69), .B2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n471), .ZN(new_n481));
  NAND3_X1  g056(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n462), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT70), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n479), .B(new_n485), .C1(G136), .C2(new_n486), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT71), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G114), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n489), .B1(new_n494), .B2(new_n462), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n481), .A2(new_n482), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT3), .B(G2104), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n495), .B(new_n496), .C1(new_n501), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  XOR2_X1   g089(.A(KEYINPUT72), .B(G88), .Z(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n512), .A2(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  NAND2_X1  g095(.A1(new_n513), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(new_n522), .B1(new_n507), .B2(new_n508), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G51), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n516), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n511), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n514), .A2(new_n531), .B1(new_n516), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AOI22_X1  g109(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n511), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n514), .A2(new_n537), .B1(new_n516), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  XNOR2_X1  g120(.A(KEYINPUT73), .B(G65), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n509), .A2(new_n546), .B1(G78), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G91), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n547), .A2(new_n511), .B1(new_n548), .B2(new_n514), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT9), .B1(new_n516), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(KEYINPUT6), .A2(G651), .ZN(new_n554));
  NAND2_X1  g129(.A1(KEYINPUT6), .A2(G651), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(new_n557), .A3(G53), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n550), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G74), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n507), .A2(new_n563), .A3(new_n508), .ZN(new_n564));
  AOI22_X1  g139(.A1(G49), .A2(new_n556), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n509), .A2(new_n513), .A3(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G288));
  NAND2_X1  g142(.A1(G73), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  AND2_X1   g145(.A1(KEYINPUT5), .A2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(KEYINPUT5), .A2(G543), .ZN(new_n572));
  OAI211_X1 g147(.A(KEYINPUT74), .B(G61), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT74), .B1(new_n509), .B2(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n507), .A2(new_n508), .B1(new_n554), .B2(new_n555), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G86), .B1(new_n556), .B2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n511), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n514), .A2(new_n582), .B1(new_n516), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n581), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT76), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n511), .B1(new_n589), .B2(new_n516), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT77), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  OAI221_X1 g167(.A(new_n592), .B1(new_n516), .B2(new_n589), .C1(new_n588), .C2(new_n511), .ZN(new_n593));
  AND3_X1   g168(.A1(new_n509), .A2(new_n513), .A3(G92), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(KEYINPUT10), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n591), .A2(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n587), .B1(G868), .B2(new_n597), .ZN(G321));
  XOR2_X1   g173(.A(G321), .B(KEYINPUT78), .Z(G284));
  MUX2_X1   g174(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g175(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g176(.A(KEYINPUT79), .B(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n597), .B1(G860), .B2(new_n602), .ZN(G148));
  NAND2_X1  g178(.A1(new_n597), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g182(.A1(new_n469), .A2(G2105), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n502), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(G2100), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n486), .A2(G135), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n483), .A2(G123), .ZN(new_n614));
  OR2_X1    g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n615), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NAND2_X1  g193(.A1(new_n612), .A2(new_n618), .ZN(G156));
  XOR2_X1   g194(.A(KEYINPUT15), .B(G2435), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2438), .ZN(new_n621));
  XOR2_X1   g196(.A(G2427), .B(G2430), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT82), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n621), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(G1341), .B(G1348), .Z(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2443), .B(G2446), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT81), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n630), .A2(new_n634), .ZN(new_n636));
  AND3_X1   g211(.A1(new_n635), .A2(G14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT83), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(G2072), .A2(G2078), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n442), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n642), .A2(KEYINPUT84), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(KEYINPUT84), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n648), .A3(new_n644), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n642), .B(KEYINPUT17), .ZN(new_n650));
  OAI211_X1 g225(.A(new_n649), .B(new_n640), .C1(new_n650), .C2(new_n644), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n644), .A3(new_n639), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n646), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2096), .B(G2100), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  AND2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT20), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n658), .A2(new_n659), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n657), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n657), .B2(new_n663), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1981), .B(G1986), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT86), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(G229));
  OR2_X1    g249(.A1(G6), .A2(G16), .ZN(new_n675));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(G305), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT32), .B(G1981), .Z(new_n678));
  OR2_X1    g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(G23), .ZN(new_n680));
  INV_X1    g255(.A(G288), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n676), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT89), .Z(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT33), .B(G1976), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI22_X1  g260(.A1(new_n683), .A2(new_n684), .B1(new_n677), .B2(new_n678), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n676), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n676), .ZN(new_n688));
  INV_X1    g263(.A(G1971), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AND4_X1   g265(.A1(new_n679), .A2(new_n685), .A3(new_n686), .A4(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G24), .ZN(new_n695));
  XOR2_X1   g270(.A(G290), .B(KEYINPUT88), .Z(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1986), .ZN(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G25), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n486), .A2(G131), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT87), .Z(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G107), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G2105), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n483), .B2(G119), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n700), .B1(new_n708), .B2(new_n699), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  XOR2_X1   g285(.A(new_n709), .B(new_n710), .Z(new_n711));
  NOR2_X1   g286(.A1(new_n698), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n693), .A2(new_n694), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n713), .A2(KEYINPUT90), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT90), .B(KEYINPUT36), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n699), .A2(G35), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G162), .B2(new_n699), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G2090), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n719), .B(new_n721), .Z(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT26), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(G105), .B2(new_n608), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n486), .A2(G141), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n483), .A2(G129), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G32), .B(new_n730), .S(G29), .Z(new_n731));
  XOR2_X1   g306(.A(KEYINPUT27), .B(G1996), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G164), .A2(G29), .ZN(new_n734));
  OR2_X1    g309(.A1(G27), .A2(G29), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  AND2_X1   g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n699), .B1(KEYINPUT24), .B2(G34), .ZN(new_n740));
  OAI22_X1  g315(.A1(G160), .A2(new_n699), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n737), .A2(G2078), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G4), .A2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n597), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(G1348), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n745), .B(new_n746), .Z(new_n747));
  OR4_X1    g322(.A1(new_n722), .A2(new_n733), .A3(new_n743), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n676), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n676), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT94), .Z(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n754));
  AND3_X1   g329(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n486), .A2(G139), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n502), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n756), .B(new_n757), .C1(new_n462), .C2(new_n758), .ZN(new_n759));
  MUX2_X1   g334(.A(G33), .B(new_n759), .S(G29), .Z(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G2072), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n751), .A2(new_n752), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n699), .A2(G26), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT28), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n486), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n483), .A2(G128), .ZN(new_n766));
  OR2_X1    g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n764), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2067), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n753), .A2(new_n761), .A3(new_n762), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n617), .A2(new_n699), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT93), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n676), .A2(G21), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G168), .B2(new_n676), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G28), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT30), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n779), .B2(KEYINPUT30), .ZN(new_n781));
  OR2_X1    g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  NAND2_X1  g357(.A1(KEYINPUT31), .A2(G11), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n676), .A2(G19), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n540), .B2(new_n676), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n778), .B(new_n784), .C1(G1341), .C2(new_n786), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n774), .B(new_n787), .C1(G1341), .C2(new_n786), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n676), .A2(G20), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT23), .Z(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G299), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT96), .B(G1956), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n737), .A2(G2078), .B1(new_n738), .B2(new_n742), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n788), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n748), .A2(new_n772), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n715), .A2(new_n717), .A3(new_n796), .ZN(G311));
  NAND3_X1  g372(.A1(new_n715), .A2(new_n717), .A3(new_n796), .ZN(G150));
  AOI22_X1  g373(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n511), .ZN(new_n800));
  INV_X1    g375(.A(G93), .ZN(new_n801));
  INV_X1    g376(.A(G55), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n514), .A2(new_n801), .B1(new_n516), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G860), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT37), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n804), .B(KEYINPUT97), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(new_n540), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT97), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n804), .B(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n540), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n597), .A2(G559), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT98), .Z(new_n820));
  OAI21_X1  g395(.A(new_n805), .B1(new_n817), .B2(new_n818), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n807), .B1(new_n820), .B2(new_n821), .ZN(G145));
  XNOR2_X1  g397(.A(G162), .B(G160), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(new_n617), .Z(new_n824));
  AOI22_X1  g399(.A1(G130), .A2(new_n483), .B1(new_n486), .B2(G142), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT100), .ZN(new_n827));
  INV_X1    g402(.A(G118), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n826), .A2(new_n827), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n827), .B2(new_n826), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT101), .ZN(new_n832));
  INV_X1    g407(.A(new_n610), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  OR3_X1    g410(.A1(new_n834), .A2(new_n835), .A3(new_n707), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n707), .B1(new_n834), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n759), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(new_n730), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n730), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n505), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n769), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n841), .A2(new_n505), .A3(new_n842), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n846), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n769), .B1(new_n848), .B2(new_n843), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n838), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n847), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n853), .A2(new_n836), .A3(new_n837), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n838), .B1(new_n849), .B2(new_n847), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n856), .A2(new_n851), .A3(new_n850), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n824), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n824), .A3(new_n850), .ZN(new_n859));
  INV_X1    g434(.A(G37), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT40), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(G395));
  XNOR2_X1  g439(.A(new_n597), .B(G299), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(KEYINPUT41), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n814), .B(new_n604), .ZN(new_n869));
  MUX2_X1   g444(.A(new_n868), .B(new_n865), .S(new_n869), .Z(new_n870));
  XNOR2_X1  g445(.A(G288), .B(KEYINPUT103), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(G290), .Z(new_n872));
  XNOR2_X1  g447(.A(G303), .B(G305), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(KEYINPUT104), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT42), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n870), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G868), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(G868), .B2(new_n804), .ZN(G295));
  OAI21_X1  g457(.A(new_n881), .B1(G868), .B2(new_n804), .ZN(G331));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n875), .A2(new_n877), .ZN(new_n885));
  XNOR2_X1  g460(.A(G286), .B(G171), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n809), .A2(new_n813), .A3(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n809), .B2(new_n813), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(KEYINPUT106), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n888), .A2(new_n865), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n887), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n866), .B(new_n867), .C1(new_n893), .C2(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n885), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(new_n860), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n878), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n884), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n895), .A2(new_n860), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n868), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n890), .A2(new_n865), .A3(new_n887), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n885), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n900), .A2(new_n904), .A3(KEYINPUT43), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n896), .A2(new_n884), .A3(new_n898), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n900), .B2(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT44), .ZN(new_n910));
  OAI22_X1  g485(.A1(new_n906), .A2(new_n907), .B1(new_n908), .B2(new_n910), .ZN(G397));
  NAND2_X1  g486(.A1(new_n708), .A2(new_n710), .ZN(new_n912));
  INV_X1    g487(.A(G1996), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n730), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G2067), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n769), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI22_X1  g492(.A1(new_n912), .A2(new_n917), .B1(G2067), .B2(new_n769), .ZN(new_n918));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n500), .B1(new_n463), .B2(new_n464), .ZN(new_n920));
  AOI22_X1  g495(.A1(new_n920), .A2(KEYINPUT4), .B1(new_n502), .B2(new_n503), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n462), .B1(new_n491), .B2(new_n493), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n496), .B1(new_n922), .B2(new_n488), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n919), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT107), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n505), .A2(new_n926), .A3(new_n919), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n473), .A2(new_n474), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(G2105), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n466), .B1(new_n486), .B2(G137), .ZN(new_n932));
  XOR2_X1   g507(.A(KEYINPUT108), .B(G40), .Z(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n918), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n707), .B(new_n710), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT110), .Z(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n939), .B2(new_n917), .ZN(new_n940));
  INV_X1    g515(.A(new_n936), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n941), .A2(G1986), .A3(G290), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n940), .B1(KEYINPUT48), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(KEYINPUT48), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n916), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n936), .B1(new_n730), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n936), .A2(new_n913), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n951), .B(KEYINPUT47), .Z(new_n952));
  NOR2_X1   g527(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(KEYINPUT121), .B(KEYINPUT51), .Z(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT119), .B1(G168), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT119), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n957), .B(G8), .C1(new_n523), .C2(new_n527), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT122), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n935), .B1(new_n924), .B2(KEYINPUT50), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n966), .B(new_n919), .C1(new_n921), .C2(new_n923), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n738), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT45), .B1(new_n505), .B2(new_n919), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n928), .A2(G1384), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(new_n921), .B2(new_n923), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n468), .A2(new_n475), .A3(new_n933), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n777), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n968), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G8), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n954), .B1(new_n964), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n955), .B1(new_n968), .B2(new_n974), .ZN(new_n978));
  OR2_X1    g553(.A1(new_n959), .A2(KEYINPUT51), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(KEYINPUT120), .A3(new_n959), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT120), .B1(new_n975), .B2(new_n959), .ZN(new_n983));
  OAI22_X1  g558(.A1(new_n977), .A2(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n564), .A2(G651), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n513), .A2(G49), .A3(G543), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n566), .A2(new_n987), .A3(new_n988), .A4(G1976), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n565), .A2(KEYINPUT112), .A3(G1976), .A4(new_n566), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n972), .A2(new_n505), .A3(new_n919), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(G288), .B2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n993), .A2(G8), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n924), .B2(new_n935), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n991), .A2(new_n992), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT52), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n576), .A2(new_n1003), .A3(new_n578), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n576), .B2(new_n578), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT113), .B(new_n1002), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT113), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n998), .B1(new_n1007), .B2(KEYINPUT49), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1001), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n689), .B1(new_n969), .B2(new_n973), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n924), .A2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(G2090), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n972), .A4(new_n967), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G8), .ZN(new_n1015));
  OAI21_X1  g590(.A(G8), .B1(new_n512), .B2(new_n518), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  AND4_X1   g596(.A1(new_n1021), .A2(new_n1014), .A3(G8), .A4(new_n1018), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n955), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1009), .B(new_n1020), .C1(new_n1022), .C2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n935), .B1(new_n505), .B2(new_n970), .ZN(new_n1026));
  INV_X1    g601(.A(G2078), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n924), .A2(new_n928), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(KEYINPUT123), .A2(KEYINPUT53), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1011), .A2(new_n972), .A3(new_n967), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n752), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1030), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G171), .ZN(new_n1037));
  NOR4_X1   g612(.A1(new_n985), .A2(new_n986), .A3(new_n1025), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1014), .A2(G8), .A3(new_n1018), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT111), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1023), .A2(new_n1021), .A3(new_n1018), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1009), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n998), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n681), .A2(new_n995), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1044), .B1(new_n1008), .B2(new_n1006), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(new_n1004), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT114), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1042), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n976), .A2(G286), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1052), .B1(new_n1025), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1009), .A2(new_n1020), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1057), .A2(KEYINPUT63), .A3(new_n1058), .A4(new_n1053), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1025), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1029), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1027), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n475), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n971), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n468), .B(KEYINPUT124), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n929), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1063), .A2(new_n1069), .A3(G301), .A4(new_n1033), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(G171), .B1(new_n1029), .B2(new_n1062), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(KEYINPUT125), .A3(new_n1033), .A4(new_n1069), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1074), .A3(new_n1037), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT126), .B1(new_n1036), .B2(G171), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1063), .A2(new_n1069), .A3(new_n1033), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1079), .B2(G171), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT126), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(G301), .A4(new_n1031), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1078), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1061), .A2(new_n1077), .A3(new_n984), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1032), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1026), .A2(new_n1028), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n559), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(new_n1093), .B2(new_n549), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n550), .A2(new_n559), .A3(new_n1091), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1348), .B1(new_n965), .B2(new_n967), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n994), .A2(G2067), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n597), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(KEYINPUT60), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1026), .A2(new_n913), .A3(new_n1028), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n994), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1104), .B1(new_n1108), .B2(new_n540), .ZN(new_n1109));
  AOI211_X1 g684(.A(KEYINPUT59), .B(new_n812), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1097), .B(new_n1103), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n597), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1096), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1096), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1090), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1093), .A2(new_n549), .A3(new_n1092), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1091), .B1(new_n550), .B2(new_n559), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT116), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1094), .A2(new_n1130), .A3(new_n1095), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1117), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT117), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1117), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1114), .A3(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1116), .A2(new_n1126), .B1(new_n1120), .B2(new_n1137), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1051), .B(new_n1060), .C1(new_n1085), .C2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1137), .A2(new_n1120), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT60), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1103), .A2(new_n1097), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT61), .B1(new_n1148), .B2(KEYINPUT118), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1119), .B1(new_n1149), .B2(new_n1123), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1142), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1084), .A2(new_n1058), .A3(new_n1057), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n963), .A2(new_n978), .ZN(new_n1153));
  OAI22_X1  g728(.A1(new_n1153), .A2(new_n954), .B1(new_n978), .B2(new_n979), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n982), .A2(new_n983), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1154), .A2(new_n1155), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1151), .A2(new_n1152), .A3(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1157), .A2(KEYINPUT127), .A3(new_n1060), .A4(new_n1051), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1038), .B1(new_n1141), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n936), .A2(G1986), .A3(G290), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n942), .A2(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT109), .Z(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n940), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n953), .B1(new_n1159), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g739(.A1(new_n637), .A2(new_n460), .A3(G227), .ZN(new_n1166));
  NOR2_X1   g740(.A1(G229), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g741(.A(new_n1167), .B1(new_n858), .B2(new_n861), .ZN(new_n1168));
  NOR2_X1   g742(.A1(new_n1168), .A2(new_n906), .ZN(G308));
  OAI221_X1 g743(.A(new_n1167), .B1(new_n858), .B2(new_n861), .C1(new_n899), .C2(new_n905), .ZN(G225));
endmodule


