//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1131, new_n1132;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(KEYINPUT66), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n475), .A2(KEYINPUT67), .A3(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G137), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT68), .Z(G160));
  AOI21_X1  g060(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n463), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(G136), .B2(new_n481), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT69), .ZN(G162));
  NAND2_X1  g067(.A1(new_n463), .A2(G138), .ZN(new_n493));
  OR2_X1    g068(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n470), .A3(new_n466), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT70), .A2(G114), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT70), .A2(G114), .ZN(new_n503));
  OAI21_X1  g078(.A(G2105), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(G126), .A2(new_n486), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n500), .A2(KEYINPUT72), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT72), .B1(new_n500), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT73), .B1(new_n511), .B2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(new_n514), .A3(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(new_n515), .B1(KEYINPUT5), .B2(new_n511), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(G543), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT74), .Z(new_n526));
  AOI21_X1  g101(.A(new_n523), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n522), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n530), .B(new_n532), .C1(new_n533), .C2(new_n521), .ZN(new_n534));
  INV_X1    g109(.A(new_n518), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(G89), .B2(new_n535), .ZN(G168));
  AOI22_X1  g111(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n523), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT75), .B(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n518), .A2(new_n539), .B1(new_n521), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AND2_X1   g117(.A1(new_n516), .A2(G56), .ZN(new_n543));
  AND2_X1   g118(.A1(G68), .A2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n546), .ZN(new_n548));
  INV_X1    g123(.A(new_n521), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n535), .A2(G81), .B1(G43), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n516), .A2(G65), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n523), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n516), .A2(G91), .A3(new_n517), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT77), .B(KEYINPUT9), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n549), .A2(G53), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n521), .A2(new_n565), .B1(KEYINPUT77), .B2(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n562), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  XOR2_X1   g144(.A(G168), .B(KEYINPUT78), .Z(G286));
  NAND2_X1  g145(.A1(new_n535), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n549), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  OR3_X1    g151(.A1(new_n575), .A2(new_n576), .A3(new_n523), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n521), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n549), .A2(KEYINPUT80), .A3(G48), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n580), .A2(new_n581), .B1(new_n535), .B2(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n576), .B1(new_n575), .B2(new_n523), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n577), .A2(new_n582), .A3(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n535), .A2(G85), .B1(G47), .B2(new_n549), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n523), .B2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n535), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  NAND2_X1  g165(.A1(new_n516), .A2(G66), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT81), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n523), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(G54), .B2(new_n549), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n588), .B1(new_n597), .B2(G868), .ZN(G321));
  NOR2_X1   g174(.A1(G299), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G286), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  AOI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n597), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g184(.A1(new_n466), .A2(new_n470), .A3(new_n475), .ZN(new_n610));
  XOR2_X1   g185(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n611));
  XNOR2_X1  g186(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT13), .Z(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(G2100), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(G2100), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n481), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n486), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n463), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT83), .B(G2096), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n614), .A2(new_n615), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT84), .Z(G156));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT85), .B(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT86), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT87), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1961), .B(G1966), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n656), .A2(new_n658), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n661), .A3(new_n659), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n666), .C1(new_n661), .C2(new_n665), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1981), .B(G1986), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G229));
  MUX2_X1   g248(.A(G6), .B(G305), .S(G16), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT89), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT32), .B(G1981), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT90), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G22), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(G1971), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(G23), .ZN(new_n685));
  INV_X1    g260(.A(G288), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n678), .A2(new_n679), .A3(new_n684), .A4(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT91), .Z(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  MUX2_X1   g269(.A(G24), .B(G290), .S(G16), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n481), .A2(G131), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n486), .A2(G119), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n463), .A2(G107), .ZN(new_n699));
  OAI21_X1  g274(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n697), .B(new_n698), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT88), .Z(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n696), .B(new_n706), .C1(KEYINPUT92), .C2(KEYINPUT36), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n693), .A2(new_n694), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(G4), .A2(G16), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n597), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT93), .B(G1348), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G2078), .ZN(new_n716));
  NAND2_X1  g291(.A1(G164), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G27), .B2(G29), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n715), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G29), .A2(G33), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT97), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT25), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n481), .A2(G139), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT98), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n723), .A2(KEYINPUT98), .A3(new_n724), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n466), .A2(new_n470), .A3(G127), .ZN(new_n729));
  INV_X1    g304(.A(G115), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n474), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n727), .A2(new_n728), .B1(G2105), .B2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n721), .B1(new_n732), .B2(G29), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n733), .A2(G2072), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G2072), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G35), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G162), .B2(G29), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT29), .B(G2090), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n734), .B(new_n739), .C1(new_n737), .C2(new_n738), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n680), .A2(G21), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G168), .B2(new_n680), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1966), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n718), .A2(new_n716), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G26), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT28), .Z(new_n747));
  OAI21_X1  g322(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n748));
  INV_X1    g323(.A(G116), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT95), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n481), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n486), .A2(G128), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n747), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT96), .B(G2067), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT30), .B(G28), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n760), .B1(new_n745), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n620), .B2(new_n745), .ZN(new_n763));
  NOR4_X1   g338(.A1(new_n743), .A2(new_n744), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n719), .A2(new_n740), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G19), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n552), .B2(G16), .ZN(new_n767));
  XOR2_X1   g342(.A(KEYINPUT94), .B(G1341), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n680), .A2(G20), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT100), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G299), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n680), .A2(G5), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G171), .B2(new_n680), .ZN(new_n776));
  INV_X1    g351(.A(G1961), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(G29), .A2(G32), .ZN(new_n779));
  NAND3_X1  g354(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT26), .Z(new_n781));
  NAND2_X1  g356(.A1(new_n481), .A2(G141), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n486), .A2(G129), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n475), .A2(G105), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n781), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT99), .Z(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n779), .B1(new_n787), .B2(G29), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n769), .A2(new_n774), .A3(new_n778), .A4(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G34), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(KEYINPUT24), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n792), .A2(KEYINPUT24), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n745), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G160), .B2(new_n745), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2084), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n765), .A2(new_n791), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n710), .A2(new_n711), .A3(new_n798), .ZN(G150));
  INV_X1    g374(.A(G150), .ZN(G311));
  AOI22_X1  g375(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(new_n523), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT103), .B(G93), .ZN(new_n803));
  INV_X1    g378(.A(G55), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n518), .A2(new_n803), .B1(new_n804), .B2(new_n521), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n551), .B(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n596), .A2(new_n604), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT102), .B(KEYINPUT104), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT39), .ZN(new_n815));
  AOI21_X1  g390(.A(G860), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n807), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  NAND2_X1  g395(.A1(new_n786), .A2(new_n732), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n785), .B2(new_n732), .ZN(new_n822));
  OAI211_X1 g397(.A(G126), .B(G2105), .C1(new_n468), .C2(new_n469), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n824));
  INV_X1    g399(.A(G114), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n463), .B1(new_n826), .B2(new_n501), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n823), .B1(new_n827), .B2(new_n505), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n499), .B2(new_n497), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n755), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n822), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n481), .A2(G142), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n486), .A2(G130), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n463), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n832), .B(new_n833), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n701), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT105), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n612), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT106), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n831), .A2(new_n839), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n841), .B(new_n842), .Z(new_n843));
  XNOR2_X1  g418(.A(G160), .B(new_n620), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G162), .Z(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n842), .A3(new_n840), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT40), .Z(G395));
  XOR2_X1   g426(.A(new_n596), .B(G299), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT107), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n852), .B(KEYINPUT41), .Z(new_n854));
  XOR2_X1   g429(.A(new_n606), .B(new_n808), .Z(new_n855));
  MUX2_X1   g430(.A(new_n853), .B(new_n854), .S(new_n855), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT42), .ZN(new_n857));
  XNOR2_X1  g432(.A(G305), .B(G290), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n686), .B(G303), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G868), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(G868), .B2(new_n806), .ZN(G295));
  OAI21_X1  g438(.A(new_n862), .B1(G868), .B2(new_n806), .ZN(G331));
  NOR2_X1   g439(.A1(G168), .A2(G171), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n601), .B2(G171), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(new_n808), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n854), .ZN(new_n868));
  INV_X1    g443(.A(new_n852), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n869), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n848), .B1(new_n870), .B2(new_n860), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n860), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT43), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n875));
  INV_X1    g450(.A(new_n860), .ZN(new_n876));
  INV_X1    g451(.A(new_n867), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n853), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n878), .B2(new_n868), .ZN(new_n879));
  NOR3_X1   g454(.A1(new_n871), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(KEYINPUT44), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n871), .A2(KEYINPUT43), .A3(new_n879), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n872), .A2(new_n873), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(KEYINPUT43), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n884), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g460(.A(KEYINPUT127), .ZN(new_n886));
  AOI21_X1  g461(.A(G1384), .B1(new_n500), .B2(new_n507), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n471), .A2(new_n472), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(G2105), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(G40), .A3(new_n482), .A4(new_n480), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT109), .Z(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n755), .B(G2067), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n898), .B1(G1996), .B2(new_n785), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n894), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(G1996), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n787), .ZN(new_n903));
  XOR2_X1   g478(.A(new_n903), .B(KEYINPUT108), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n701), .B(new_n705), .ZN(new_n905));
  AOI211_X1 g480(.A(new_n900), .B(new_n904), .C1(new_n895), .C2(new_n905), .ZN(new_n906));
  NOR3_X1   g481(.A1(new_n901), .A2(G1986), .A3(G290), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(KEYINPUT48), .Z(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n902), .B(KEYINPUT46), .Z(new_n910));
  OAI21_X1  g485(.A(new_n895), .B1(new_n785), .B2(new_n898), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n912), .B(KEYINPUT47), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n756), .A2(G2067), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n904), .A2(new_n900), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n702), .A2(new_n705), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(new_n896), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n914), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G8), .ZN(new_n921));
  INV_X1    g496(.A(new_n893), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n922), .B2(new_n887), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n686), .A2(G1976), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT111), .B(G1976), .Z(new_n925));
  AOI21_X1  g500(.A(KEYINPUT52), .B1(G288), .B2(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n924), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(KEYINPUT52), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT49), .ZN(new_n930));
  NAND2_X1  g505(.A1(G305), .A2(G1981), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(G305), .A2(G1981), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n933), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(KEYINPUT49), .A3(new_n931), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n936), .A3(new_n923), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n500), .A2(new_n507), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT72), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n829), .A2(KEYINPUT72), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n944));
  NOR4_X1   g519(.A1(new_n829), .A2(new_n944), .A3(new_n889), .A4(G1384), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT110), .B1(new_n887), .B2(KEYINPUT45), .ZN(new_n946));
  OAI22_X1  g521(.A1(new_n943), .A2(KEYINPUT45), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n922), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n683), .ZN(new_n950));
  AOI211_X1 g525(.A(KEYINPUT50), .B(G1384), .C1(new_n500), .C2(new_n507), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(new_n893), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n952), .B1(new_n943), .B2(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(G2090), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n921), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G303), .A2(G8), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT55), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n938), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n949), .B2(G2078), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(KEYINPUT117), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT117), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n952), .B(new_n964), .C1(new_n943), .C2(new_n953), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n777), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n893), .B1(new_n889), .B2(new_n888), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n508), .B2(new_n509), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n967), .B1(new_n889), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n716), .A2(KEYINPUT53), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n962), .B(new_n966), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n893), .B1(KEYINPUT50), .B2(new_n888), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(KEYINPUT50), .B2(new_n969), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(G2090), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n949), .B2(new_n683), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n958), .B1(new_n976), .B2(new_n921), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n960), .A2(G171), .A3(new_n972), .A4(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1966), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n970), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n980), .A2(KEYINPUT113), .ZN(new_n981));
  INV_X1    g556(.A(G2084), .ZN(new_n982));
  INV_X1    g557(.A(new_n954), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n980), .A2(KEYINPUT113), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G168), .ZN(new_n986));
  OAI21_X1  g561(.A(G8), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G168), .B1(new_n981), .B2(new_n984), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT51), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n990), .B(G8), .C1(new_n985), .C2(new_n986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n978), .B1(new_n992), .B2(KEYINPUT62), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(new_n994), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n956), .A2(new_n959), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n601), .A2(G8), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n981), .B2(new_n984), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n997), .A2(new_n960), .A3(KEYINPUT63), .A4(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n960), .A2(new_n977), .A3(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(KEYINPUT63), .ZN(new_n1002));
  AND4_X1   g577(.A1(new_n959), .A2(new_n956), .A3(new_n937), .A4(new_n929), .ZN(new_n1003));
  NOR2_X1   g578(.A1(G288), .A2(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n933), .B1(new_n937), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1007));
  INV_X1    g582(.A(new_n923), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n1006), .B2(KEYINPUT112), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1003), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1002), .A2(new_n1010), .A3(KEYINPUT114), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT114), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n996), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n939), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(new_n944), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n887), .A2(KEYINPUT110), .A3(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1017), .A2(new_n967), .A3(KEYINPUT53), .A4(new_n716), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n962), .A2(new_n966), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(G171), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(G171), .B2(new_n972), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT126), .B(KEYINPUT54), .Z(new_n1022));
  OR2_X1    g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1019), .A2(G171), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1024), .B(KEYINPUT54), .C1(G171), .C2(new_n972), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1025), .A2(new_n977), .A3(new_n960), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n992), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1348), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n963), .A2(new_n1028), .A3(new_n965), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n922), .A2(new_n887), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(G2067), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(KEYINPUT60), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(KEYINPUT124), .A3(new_n596), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n596), .B1(new_n1032), .B2(KEYINPUT124), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1034), .A2(new_n1035), .B1(KEYINPUT124), .B2(new_n1032), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(KEYINPUT60), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OR3_X1    g614(.A1(new_n560), .A2(KEYINPUT115), .A3(new_n561), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT115), .B1(new_n560), .B2(new_n561), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n567), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT116), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n562), .A2(KEYINPUT57), .A3(new_n567), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1047), .A3(new_n1043), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1956), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n974), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT56), .B(G2072), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n948), .A2(new_n922), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1049), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT61), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1049), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1053), .A2(new_n1051), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT61), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1054), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1036), .A2(new_n1039), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT58), .B(G1341), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1030), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT119), .B(G1996), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n893), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n947), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n969), .A2(new_n889), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(new_n1017), .A3(new_n1068), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT120), .A3(new_n1066), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n551), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1064), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT59), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1074), .A2(KEYINPUT120), .A3(new_n1066), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT120), .B1(new_n1074), .B2(new_n1066), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n552), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(KEYINPUT121), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1078), .B1(new_n1080), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1077), .B1(new_n1083), .B2(KEYINPUT121), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1064), .A3(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1086), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1063), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1060), .B1(new_n1037), .B2(new_n596), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1054), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT118), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1027), .B1(new_n1096), .B2(KEYINPUT125), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1092), .A2(new_n1098), .A3(new_n1095), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1013), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  XOR2_X1   g675(.A(G290), .B(G1986), .Z(new_n1101));
  OAI21_X1  g676(.A(new_n906), .B1(new_n901), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n886), .B(new_n920), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1057), .A2(new_n1062), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1032), .A2(KEYINPUT124), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1032), .A2(KEYINPUT124), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n597), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(new_n1107), .B2(new_n1033), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1108), .B2(new_n1038), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1080), .A2(new_n1084), .A3(KEYINPUT122), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1077), .B(new_n552), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT122), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT123), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1085), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1109), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1095), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT125), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1027), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1099), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1002), .A2(new_n1010), .A3(KEYINPUT114), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1123), .A2(new_n1124), .B1(new_n995), .B2(new_n993), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1102), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n920), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT127), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1103), .A2(new_n1128), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g704(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1131));
  OR3_X1    g705(.A1(new_n850), .A2(G229), .A3(new_n1131), .ZN(new_n1132));
  NOR2_X1   g706(.A1(new_n1132), .A2(new_n884), .ZN(G308));
  INV_X1    g707(.A(G308), .ZN(G225));
endmodule


