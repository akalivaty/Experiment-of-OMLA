

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734;

  AND2_X1 U369 ( .A1(n680), .A2(n557), .ZN(n558) );
  NOR2_X1 U370 ( .A1(n628), .A2(n630), .ZN(n471) );
  OR2_X1 U371 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U372 ( .A(n392), .B(n391), .ZN(n561) );
  INV_X1 U373 ( .A(n542), .ZN(n517) );
  XNOR2_X1 U374 ( .A(n421), .B(G472), .ZN(n547) );
  XNOR2_X1 U375 ( .A(n383), .B(n382), .ZN(n542) );
  XNOR2_X1 U376 ( .A(n446), .B(n433), .ZN(n722) );
  XOR2_X1 U377 ( .A(KEYINPUT23), .B(n346), .Z(n378) );
  XNOR2_X1 U378 ( .A(n402), .B(n401), .ZN(n714) );
  BUF_X1 U379 ( .A(G128), .Z(n346) );
  XNOR2_X1 U380 ( .A(n395), .B(G134), .ZN(n446) );
  XNOR2_X1 U381 ( .A(G110), .B(G107), .ZN(n387) );
  INV_X1 U382 ( .A(G953), .ZN(n724) );
  NOR2_X2 U383 ( .A1(n590), .A2(n589), .ZN(n347) );
  NOR2_X2 U384 ( .A1(n512), .A2(n734), .ZN(n513) );
  AND2_X2 U385 ( .A1(n516), .A2(n515), .ZN(n723) );
  AND2_X1 U386 ( .A1(n705), .A2(n584), .ZN(n351) );
  XNOR2_X2 U387 ( .A(n583), .B(n582), .ZN(n705) );
  NOR2_X2 U388 ( .A1(n590), .A2(n589), .ZN(n672) );
  NOR2_X1 U389 ( .A1(n579), .A2(n681), .ZN(n580) );
  BUF_X2 U390 ( .A(n556), .Z(n680) );
  NOR2_X2 U391 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U392 ( .A1(n731), .A2(n733), .ZN(n477) );
  XNOR2_X1 U393 ( .A(n722), .B(G146), .ZN(n416) );
  XNOR2_X1 U394 ( .A(n387), .B(n386), .ZN(n400) );
  BUF_X1 U395 ( .A(n354), .Z(n348) );
  BUF_X1 U396 ( .A(n547), .Z(n349) );
  NOR2_X2 U397 ( .A1(n621), .A2(n617), .ZN(n589) );
  XNOR2_X1 U398 ( .A(n547), .B(n486), .ZN(n354) );
  XOR2_X1 U399 ( .A(KEYINPUT4), .B(KEYINPUT69), .Z(n720) );
  XNOR2_X1 U400 ( .A(n367), .B(G125), .ZN(n394) );
  INV_X1 U401 ( .A(G146), .ZN(n367) );
  XNOR2_X1 U402 ( .A(n394), .B(n368), .ZN(n429) );
  INV_X1 U403 ( .A(KEYINPUT10), .ZN(n368) );
  XOR2_X1 U404 ( .A(G140), .B(G137), .Z(n384) );
  XNOR2_X1 U405 ( .A(n407), .B(n710), .ZN(n418) );
  XNOR2_X1 U406 ( .A(n468), .B(KEYINPUT102), .ZN(n628) );
  NOR2_X1 U407 ( .A1(n467), .A2(n466), .ZN(n482) );
  XNOR2_X1 U408 ( .A(n429), .B(n432), .ZN(n434) );
  XNOR2_X1 U409 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U410 ( .A(n429), .B(n369), .ZN(n719) );
  BUF_X1 U411 ( .A(n479), .Z(n496) );
  XNOR2_X1 U412 ( .A(n425), .B(n424), .ZN(n495) );
  XNOR2_X1 U413 ( .A(KEYINPUT30), .B(KEYINPUT105), .ZN(n424) );
  XNOR2_X1 U414 ( .A(n444), .B(n443), .ZN(n500) );
  XNOR2_X1 U415 ( .A(n400), .B(n404), .ZN(n388) );
  XNOR2_X1 U416 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U417 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U418 ( .A(n719), .B(n372), .Z(n350) );
  XNOR2_X1 U419 ( .A(n546), .B(n545), .ZN(n664) );
  NOR2_X1 U420 ( .A1(n586), .A2(n585), .ZN(n352) );
  NOR2_X1 U421 ( .A1(n352), .A2(n588), .ZN(n353) );
  NOR2_X1 U422 ( .A1(n354), .A2(n560), .ZN(n518) );
  NOR2_X1 U423 ( .A1(n488), .A2(n348), .ZN(n489) );
  NAND2_X1 U424 ( .A1(n541), .A2(n348), .ZN(n573) );
  AND2_X2 U425 ( .A1(n355), .A2(n353), .ZN(n590) );
  NAND2_X1 U426 ( .A1(n351), .A2(n723), .ZN(n355) );
  NAND2_X1 U427 ( .A1(n533), .A2(n532), .ZN(n535) );
  XOR2_X1 U428 ( .A(n433), .B(KEYINPUT12), .Z(n356) );
  XOR2_X1 U429 ( .A(KEYINPUT67), .B(KEYINPUT19), .Z(n357) );
  XOR2_X1 U430 ( .A(n384), .B(KEYINPUT79), .Z(n358) );
  AND2_X1 U431 ( .A1(n502), .A2(n692), .ZN(n503) );
  INV_X1 U432 ( .A(n384), .ZN(n369) );
  BUF_X1 U433 ( .A(n624), .Z(n654) );
  XNOR2_X1 U434 ( .A(n434), .B(n356), .ZN(n441) );
  XNOR2_X1 U435 ( .A(n412), .B(n411), .ZN(n479) );
  XNOR2_X1 U436 ( .A(n350), .B(n379), .ZN(n601) );
  INV_X1 U437 ( .A(KEYINPUT108), .ZN(n459) );
  XNOR2_X1 U438 ( .A(n442), .B(G475), .ZN(n443) );
  INV_X1 U439 ( .A(KEYINPUT113), .ZN(n473) );
  XNOR2_X1 U440 ( .A(n462), .B(n461), .ZN(n731) );
  XNOR2_X1 U441 ( .A(n476), .B(n475), .ZN(n733) );
  XNOR2_X1 U442 ( .A(KEYINPUT15), .B(G902), .ZN(n586) );
  NAND2_X1 U443 ( .A1(n586), .A2(G234), .ZN(n359) );
  XNOR2_X1 U444 ( .A(n359), .B(KEYINPUT20), .ZN(n380) );
  AND2_X1 U445 ( .A1(n380), .A2(G221), .ZN(n360) );
  XNOR2_X1 U446 ( .A(n360), .B(KEYINPUT21), .ZN(n634) );
  INV_X1 U447 ( .A(n634), .ZN(n538) );
  NAND2_X1 U448 ( .A1(G234), .A2(G237), .ZN(n361) );
  XNOR2_X1 U449 ( .A(n361), .B(KEYINPUT14), .ZN(n362) );
  XNOR2_X1 U450 ( .A(KEYINPUT76), .B(n362), .ZN(n363) );
  NAND2_X1 U451 ( .A1(G952), .A2(n363), .ZN(n652) );
  NOR2_X1 U452 ( .A1(n652), .A2(G953), .ZN(n523) );
  AND2_X1 U453 ( .A1(n363), .A2(G953), .ZN(n364) );
  NAND2_X1 U454 ( .A1(G902), .A2(n364), .ZN(n522) );
  NOR2_X1 U455 ( .A1(n522), .A2(G900), .ZN(n365) );
  NOR2_X1 U456 ( .A1(n523), .A2(n365), .ZN(n366) );
  NOR2_X1 U457 ( .A1(n538), .A2(n366), .ZN(n463) );
  XOR2_X1 U458 ( .A(KEYINPUT24), .B(KEYINPUT81), .Z(n371) );
  XNOR2_X1 U459 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n370) );
  XNOR2_X1 U460 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U461 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n374) );
  NAND2_X1 U462 ( .A1(G234), .A2(n724), .ZN(n373) );
  XNOR2_X1 U463 ( .A(n374), .B(n373), .ZN(n445) );
  NAND2_X1 U464 ( .A1(G221), .A2(n445), .ZN(n376) );
  XNOR2_X1 U465 ( .A(G110), .B(G119), .ZN(n375) );
  XNOR2_X1 U466 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U467 ( .A(n378), .B(n377), .ZN(n379) );
  INV_X1 U468 ( .A(G902), .ZN(n456) );
  NAND2_X1 U469 ( .A1(n601), .A2(n456), .ZN(n383) );
  NAND2_X1 U470 ( .A1(G217), .A2(n380), .ZN(n381) );
  XNOR2_X1 U471 ( .A(KEYINPUT25), .B(n381), .ZN(n382) );
  XNOR2_X2 U472 ( .A(G143), .B(G128), .ZN(n395) );
  XOR2_X1 U473 ( .A(KEYINPUT71), .B(G131), .Z(n433) );
  NAND2_X1 U474 ( .A1(G227), .A2(n724), .ZN(n385) );
  XNOR2_X1 U475 ( .A(n358), .B(n385), .ZN(n389) );
  INV_X1 U476 ( .A(G104), .ZN(n386) );
  XNOR2_X1 U477 ( .A(n720), .B(G101), .ZN(n404) );
  XNOR2_X1 U478 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U479 ( .A(n416), .B(n390), .ZN(n607) );
  NAND2_X1 U480 ( .A1(n607), .A2(n456), .ZN(n392) );
  XOR2_X1 U481 ( .A(KEYINPUT73), .B(G469), .Z(n391) );
  AND2_X1 U482 ( .A1(n517), .A2(n561), .ZN(n393) );
  AND2_X1 U483 ( .A1(n463), .A2(n393), .ZN(n494) );
  XNOR2_X1 U484 ( .A(n395), .B(n394), .ZN(n399) );
  XNOR2_X1 U485 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n397) );
  NAND2_X1 U486 ( .A1(n724), .A2(G224), .ZN(n396) );
  XNOR2_X1 U487 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U488 ( .A(n399), .B(n398), .ZN(n403) );
  INV_X1 U489 ( .A(n400), .ZN(n402) );
  XNOR2_X1 U490 ( .A(KEYINPUT16), .B(G122), .ZN(n401) );
  XNOR2_X1 U491 ( .A(n714), .B(n403), .ZN(n408) );
  INV_X1 U492 ( .A(n404), .ZN(n407) );
  XOR2_X1 U493 ( .A(G113), .B(G116), .Z(n406) );
  XNOR2_X1 U494 ( .A(G119), .B(KEYINPUT3), .ZN(n405) );
  XNOR2_X1 U495 ( .A(n406), .B(n405), .ZN(n710) );
  XNOR2_X1 U496 ( .A(n408), .B(n418), .ZN(n593) );
  NAND2_X1 U497 ( .A1(n593), .A2(n586), .ZN(n412) );
  NOR2_X1 U498 ( .A1(G237), .A2(G902), .ZN(n409) );
  XNOR2_X1 U499 ( .A(n409), .B(KEYINPUT78), .ZN(n423) );
  INV_X1 U500 ( .A(G210), .ZN(n410) );
  OR2_X1 U501 ( .A1(n423), .A2(n410), .ZN(n411) );
  XOR2_X1 U502 ( .A(KEYINPUT77), .B(KEYINPUT38), .Z(n413) );
  XNOR2_X1 U503 ( .A(n496), .B(n413), .ZN(n626) );
  AND2_X1 U504 ( .A1(n494), .A2(n626), .ZN(n426) );
  XNOR2_X1 U505 ( .A(G137), .B(KEYINPUT92), .ZN(n414) );
  XOR2_X1 U506 ( .A(n414), .B(KEYINPUT5), .Z(n415) );
  XNOR2_X1 U507 ( .A(n416), .B(n415), .ZN(n420) );
  NOR2_X1 U508 ( .A1(G953), .A2(G237), .ZN(n435) );
  NAND2_X1 U509 ( .A1(n435), .A2(G210), .ZN(n417) );
  XNOR2_X1 U510 ( .A(n420), .B(n419), .ZN(n673) );
  NAND2_X1 U511 ( .A1(n673), .A2(n456), .ZN(n421) );
  INV_X1 U512 ( .A(G214), .ZN(n422) );
  OR2_X1 U513 ( .A1(n423), .A2(n422), .ZN(n625) );
  NAND2_X1 U514 ( .A1(n349), .A2(n625), .ZN(n425) );
  NAND2_X1 U515 ( .A1(n426), .A2(n495), .ZN(n428) );
  XOR2_X1 U516 ( .A(KEYINPUT84), .B(KEYINPUT39), .Z(n427) );
  XNOR2_X1 U517 ( .A(n428), .B(n427), .ZN(n514) );
  XOR2_X1 U518 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n431) );
  XNOR2_X1 U519 ( .A(G140), .B(KEYINPUT95), .ZN(n430) );
  XNOR2_X1 U520 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U521 ( .A(G143), .B(G113), .Z(n439) );
  NAND2_X1 U522 ( .A1(n435), .A2(G214), .ZN(n437) );
  XNOR2_X1 U523 ( .A(G104), .B(G122), .ZN(n436) );
  XNOR2_X1 U524 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U525 ( .A(n439), .B(n438), .Z(n440) );
  XNOR2_X1 U526 ( .A(n441), .B(n440), .ZN(n666) );
  NOR2_X1 U527 ( .A1(G902), .A2(n666), .ZN(n444) );
  XNOR2_X1 U528 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n442) );
  AND2_X1 U529 ( .A1(n445), .A2(G217), .ZN(n448) );
  INV_X1 U530 ( .A(n446), .ZN(n447) );
  XNOR2_X1 U531 ( .A(n448), .B(n447), .ZN(n455) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n450) );
  XNOR2_X1 U533 ( .A(G116), .B(KEYINPUT9), .ZN(n449) );
  XNOR2_X1 U534 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U535 ( .A(n451), .B(KEYINPUT99), .Z(n453) );
  XNOR2_X1 U536 ( .A(G107), .B(G122), .ZN(n452) );
  XNOR2_X1 U537 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U538 ( .A(n455), .B(n454), .ZN(n612) );
  NAND2_X1 U539 ( .A1(n612), .A2(n456), .ZN(n457) );
  XNOR2_X1 U540 ( .A(n457), .B(G478), .ZN(n483) );
  NOR2_X1 U541 ( .A1(n500), .A2(n483), .ZN(n458) );
  XNOR2_X1 U542 ( .A(n458), .B(KEYINPUT100), .ZN(n697) );
  INV_X1 U543 ( .A(n697), .ZN(n693) );
  NOR2_X1 U544 ( .A1(n514), .A2(n693), .ZN(n462) );
  XNOR2_X1 U545 ( .A(KEYINPUT109), .B(KEYINPUT40), .ZN(n460) );
  XOR2_X1 U546 ( .A(n463), .B(KEYINPUT72), .Z(n464) );
  NOR2_X1 U547 ( .A1(n517), .A2(n464), .ZN(n487) );
  AND2_X1 U548 ( .A1(n547), .A2(n487), .ZN(n465) );
  XOR2_X1 U549 ( .A(KEYINPUT28), .B(n465), .Z(n467) );
  XNOR2_X1 U550 ( .A(n561), .B(KEYINPUT107), .ZN(n466) );
  INV_X1 U551 ( .A(n483), .ZN(n499) );
  NAND2_X1 U552 ( .A1(n500), .A2(n499), .ZN(n468) );
  NAND2_X1 U553 ( .A1(n626), .A2(n625), .ZN(n630) );
  XOR2_X1 U554 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n469) );
  XNOR2_X1 U555 ( .A(KEYINPUT41), .B(n469), .ZN(n470) );
  XNOR2_X1 U556 ( .A(n471), .B(n470), .ZN(n655) );
  INV_X1 U557 ( .A(n655), .ZN(n472) );
  NAND2_X1 U558 ( .A1(n482), .A2(n472), .ZN(n476) );
  XOR2_X1 U559 ( .A(KEYINPUT42), .B(KEYINPUT112), .Z(n474) );
  XNOR2_X1 U560 ( .A(n477), .B(KEYINPUT46), .ZN(n504) );
  INV_X1 U561 ( .A(n625), .ZN(n478) );
  NOR2_X1 U562 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U563 ( .A(n480), .B(n357), .ZN(n526) );
  INV_X1 U564 ( .A(n526), .ZN(n481) );
  NAND2_X1 U565 ( .A1(n482), .A2(n481), .ZN(n694) );
  AND2_X1 U566 ( .A1(n500), .A2(n483), .ZN(n699) );
  NOR2_X1 U567 ( .A1(n697), .A2(n699), .ZN(n629) );
  NOR2_X1 U568 ( .A1(n694), .A2(n629), .ZN(n484) );
  XOR2_X1 U569 ( .A(KEYINPUT47), .B(n484), .Z(n493) );
  INV_X1 U570 ( .A(KEYINPUT101), .ZN(n485) );
  XNOR2_X1 U571 ( .A(n485), .B(KEYINPUT6), .ZN(n486) );
  NAND2_X1 U572 ( .A1(n487), .A2(n697), .ZN(n488) );
  NAND2_X1 U573 ( .A1(n489), .A2(n625), .ZN(n507) );
  NOR2_X1 U574 ( .A1(n507), .A2(n496), .ZN(n490) );
  XNOR2_X1 U575 ( .A(n490), .B(KEYINPUT36), .ZN(n491) );
  XNOR2_X2 U576 ( .A(n561), .B(KEYINPUT1), .ZN(n639) );
  NAND2_X1 U577 ( .A1(n491), .A2(n639), .ZN(n703) );
  INV_X1 U578 ( .A(n703), .ZN(n492) );
  NOR2_X1 U579 ( .A1(n493), .A2(n492), .ZN(n502) );
  AND2_X1 U580 ( .A1(n495), .A2(n494), .ZN(n497) );
  INV_X1 U581 ( .A(n496), .ZN(n509) );
  NAND2_X1 U582 ( .A1(n497), .A2(n509), .ZN(n498) );
  XOR2_X1 U583 ( .A(KEYINPUT106), .B(n498), .Z(n501) );
  NOR2_X1 U584 ( .A1(n500), .A2(n499), .ZN(n532) );
  NAND2_X1 U585 ( .A1(n501), .A2(n532), .ZN(n692) );
  NAND2_X1 U586 ( .A1(n504), .A2(n503), .ZN(n506) );
  XOR2_X1 U587 ( .A(KEYINPUT83), .B(KEYINPUT48), .Z(n505) );
  XNOR2_X1 U588 ( .A(n506), .B(n505), .ZN(n512) );
  NOR2_X1 U589 ( .A1(n639), .A2(n507), .ZN(n508) );
  XNOR2_X1 U590 ( .A(n508), .B(KEYINPUT43), .ZN(n510) );
  NOR2_X1 U591 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U592 ( .A(n511), .B(KEYINPUT104), .ZN(n734) );
  XNOR2_X1 U593 ( .A(n513), .B(KEYINPUT82), .ZN(n516) );
  INV_X1 U594 ( .A(n699), .ZN(n688) );
  NOR2_X1 U595 ( .A1(n514), .A2(n688), .ZN(n704) );
  INV_X1 U596 ( .A(n704), .ZN(n515) );
  NAND2_X1 U597 ( .A1(n517), .A2(n634), .ZN(n560) );
  NAND2_X1 U598 ( .A1(n518), .A2(n639), .ZN(n521) );
  INV_X1 U599 ( .A(KEYINPUT74), .ZN(n519) );
  XNOR2_X1 U600 ( .A(n519), .B(KEYINPUT33), .ZN(n520) );
  XNOR2_X1 U601 ( .A(n521), .B(n520), .ZN(n624) );
  INV_X1 U602 ( .A(n624), .ZN(n529) );
  NOR2_X1 U603 ( .A1(n522), .A2(G898), .ZN(n524) );
  NOR2_X1 U604 ( .A1(n524), .A2(n523), .ZN(n525) );
  INV_X1 U605 ( .A(KEYINPUT0), .ZN(n527) );
  XNOR2_X2 U606 ( .A(n528), .B(n527), .ZN(n566) );
  NAND2_X1 U607 ( .A1(n529), .A2(n566), .ZN(n531) );
  INV_X1 U608 ( .A(KEYINPUT34), .ZN(n530) );
  XNOR2_X1 U609 ( .A(n531), .B(n530), .ZN(n533) );
  INV_X1 U610 ( .A(KEYINPUT35), .ZN(n534) );
  XNOR2_X2 U611 ( .A(n535), .B(n534), .ZN(n556) );
  INV_X1 U612 ( .A(KEYINPUT44), .ZN(n536) );
  NAND2_X1 U613 ( .A1(n556), .A2(n536), .ZN(n537) );
  XNOR2_X1 U614 ( .A(n537), .B(KEYINPUT68), .ZN(n554) );
  NOR2_X1 U615 ( .A1(n628), .A2(n538), .ZN(n539) );
  NAND2_X1 U616 ( .A1(n566), .A2(n539), .ZN(n540) );
  XNOR2_X1 U617 ( .A(n540), .B(KEYINPUT22), .ZN(n550) );
  INV_X1 U618 ( .A(n550), .ZN(n541) );
  INV_X1 U619 ( .A(n573), .ZN(n544) );
  AND2_X1 U620 ( .A1(n639), .A2(n542), .ZN(n543) );
  NAND2_X1 U621 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U622 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n545) );
  INV_X1 U623 ( .A(n664), .ZN(n552) );
  BUF_X1 U624 ( .A(n349), .Z(n637) );
  OR2_X1 U625 ( .A1(n637), .A2(n517), .ZN(n548) );
  OR2_X1 U626 ( .A1(n548), .A2(n639), .ZN(n549) );
  OR2_X1 U627 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U628 ( .A(n551), .B(KEYINPUT103), .ZN(n600) );
  NAND2_X1 U629 ( .A1(n552), .A2(n557), .ZN(n553) );
  XNOR2_X1 U630 ( .A(n555), .B(KEYINPUT75), .ZN(n581) );
  INV_X1 U631 ( .A(n600), .ZN(n557) );
  NAND2_X1 U632 ( .A1(n558), .A2(n552), .ZN(n559) );
  NAND2_X1 U633 ( .A1(n559), .A2(KEYINPUT44), .ZN(n572) );
  INV_X1 U634 ( .A(n560), .ZN(n640) );
  NAND2_X1 U635 ( .A1(n561), .A2(n640), .ZN(n562) );
  NOR2_X1 U636 ( .A1(n637), .A2(n562), .ZN(n563) );
  NAND2_X1 U637 ( .A1(n566), .A2(n563), .ZN(n564) );
  XNOR2_X1 U638 ( .A(n564), .B(KEYINPUT93), .ZN(n684) );
  AND2_X1 U639 ( .A1(n637), .A2(n640), .ZN(n565) );
  AND2_X1 U640 ( .A1(n639), .A2(n565), .ZN(n646) );
  NAND2_X1 U641 ( .A1(n566), .A2(n646), .ZN(n568) );
  XNOR2_X1 U642 ( .A(KEYINPUT94), .B(KEYINPUT31), .ZN(n567) );
  XNOR2_X1 U643 ( .A(n568), .B(n567), .ZN(n700) );
  OR2_X1 U644 ( .A1(n684), .A2(n700), .ZN(n570) );
  INV_X1 U645 ( .A(n629), .ZN(n569) );
  NAND2_X1 U646 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U647 ( .A1(n572), .A2(n571), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n573), .B(KEYINPUT85), .ZN(n575) );
  INV_X1 U649 ( .A(n639), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n577) );
  INV_X1 U651 ( .A(KEYINPUT86), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n577), .B(n576), .ZN(n578) );
  AND2_X1 U653 ( .A1(n578), .A2(n517), .ZN(n681) );
  NAND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U655 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n582) );
  INV_X1 U656 ( .A(n586), .ZN(n584) );
  NAND2_X1 U657 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n585) );
  INV_X1 U658 ( .A(KEYINPUT2), .ZN(n617) );
  NOR2_X1 U659 ( .A1(n586), .A2(n617), .ZN(n587) );
  NOR2_X1 U660 ( .A1(n587), .A2(KEYINPUT66), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n705), .A2(n723), .ZN(n621) );
  NAND2_X1 U662 ( .A1(n672), .A2(G210), .ZN(n595) );
  XOR2_X1 U663 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT55), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n595), .B(n594), .ZN(n597) );
  NOR2_X1 U667 ( .A1(n724), .A2(G952), .ZN(n596) );
  XNOR2_X1 U668 ( .A(n596), .B(KEYINPUT89), .ZN(n676) );
  NAND2_X1 U669 ( .A1(n597), .A2(n676), .ZN(n599) );
  INV_X1 U670 ( .A(KEYINPUT56), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n599), .B(n598), .ZN(G51) );
  XOR2_X1 U672 ( .A(G110), .B(n600), .Z(G12) );
  BUF_X1 U673 ( .A(n672), .Z(n611) );
  NAND2_X1 U674 ( .A1(n611), .A2(G217), .ZN(n604) );
  XNOR2_X1 U675 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n602) );
  XNOR2_X1 U676 ( .A(n601), .B(n602), .ZN(n603) );
  XNOR2_X1 U677 ( .A(n604), .B(n603), .ZN(n605) );
  INV_X1 U678 ( .A(n676), .ZN(n615) );
  NOR2_X1 U679 ( .A1(n605), .A2(n615), .ZN(G66) );
  NAND2_X1 U680 ( .A1(n611), .A2(G469), .ZN(n609) );
  XNOR2_X1 U681 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n606) );
  XNOR2_X1 U682 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n609), .B(n608), .ZN(n610) );
  NOR2_X1 U684 ( .A1(n610), .A2(n615), .ZN(G54) );
  NAND2_X1 U685 ( .A1(n611), .A2(G478), .ZN(n614) );
  XOR2_X1 U686 ( .A(n612), .B(KEYINPUT122), .Z(n613) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n616), .A2(n615), .ZN(G63) );
  INV_X1 U689 ( .A(KEYINPUT53), .ZN(n663) );
  INV_X1 U690 ( .A(n621), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n617), .A2(KEYINPUT80), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n619), .A2(n618), .ZN(n623) );
  XOR2_X1 U693 ( .A(KEYINPUT2), .B(KEYINPUT80), .Z(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n659) );
  NOR2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n632) );
  NOR2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U699 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U700 ( .A1(n654), .A2(n633), .ZN(n650) );
  NOR2_X1 U701 ( .A1(n517), .A2(n634), .ZN(n635) );
  XOR2_X1 U702 ( .A(KEYINPUT49), .B(n635), .Z(n636) );
  NOR2_X1 U703 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U704 ( .A(KEYINPUT117), .B(n638), .ZN(n643) );
  NOR2_X1 U705 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U706 ( .A(KEYINPUT50), .B(n641), .ZN(n642) );
  NOR2_X1 U707 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U708 ( .A(n644), .B(KEYINPUT118), .ZN(n645) );
  NOR2_X1 U709 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U710 ( .A(KEYINPUT51), .B(n647), .Z(n648) );
  NOR2_X1 U711 ( .A1(n655), .A2(n648), .ZN(n649) );
  NOR2_X1 U712 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U713 ( .A(n651), .B(KEYINPUT52), .ZN(n653) );
  NOR2_X1 U714 ( .A1(n653), .A2(n652), .ZN(n657) );
  NOR2_X1 U715 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U716 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U717 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U718 ( .A(n660), .B(KEYINPUT119), .ZN(n661) );
  NAND2_X1 U719 ( .A1(n661), .A2(n724), .ZN(n662) );
  XNOR2_X1 U720 ( .A(n663), .B(n662), .ZN(G75) );
  XOR2_X1 U721 ( .A(n664), .B(G119), .Z(G21) );
  NAND2_X1 U722 ( .A1(n347), .A2(G475), .ZN(n668) );
  XOR2_X1 U723 ( .A(KEYINPUT87), .B(KEYINPUT59), .Z(n665) );
  XNOR2_X1 U724 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U725 ( .A(n668), .B(n667), .ZN(n669) );
  NAND2_X1 U726 ( .A1(n669), .A2(n676), .ZN(n671) );
  XNOR2_X1 U727 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n670) );
  XNOR2_X1 U728 ( .A(n671), .B(n670), .ZN(G60) );
  NAND2_X1 U729 ( .A1(n347), .A2(G472), .ZN(n675) );
  XNOR2_X1 U730 ( .A(n673), .B(KEYINPUT62), .ZN(n674) );
  XNOR2_X1 U731 ( .A(n675), .B(n674), .ZN(n677) );
  NAND2_X1 U732 ( .A1(n677), .A2(n676), .ZN(n679) );
  XNOR2_X1 U733 ( .A(KEYINPUT88), .B(KEYINPUT63), .ZN(n678) );
  XNOR2_X1 U734 ( .A(n679), .B(n678), .ZN(G57) );
  XNOR2_X1 U735 ( .A(n680), .B(G122), .ZN(G24) );
  XOR2_X1 U736 ( .A(G101), .B(n681), .Z(G3) );
  NAND2_X1 U737 ( .A1(n697), .A2(n684), .ZN(n682) );
  XNOR2_X1 U738 ( .A(n682), .B(KEYINPUT114), .ZN(n683) );
  XNOR2_X1 U739 ( .A(G104), .B(n683), .ZN(G6) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n686) );
  NAND2_X1 U741 ( .A1(n684), .A2(n699), .ZN(n685) );
  XNOR2_X1 U742 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U743 ( .A(G107), .B(n687), .ZN(G9) );
  NOR2_X1 U744 ( .A1(n694), .A2(n688), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n346), .B(KEYINPUT29), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n690), .B(n689), .ZN(G30) );
  XOR2_X1 U747 ( .A(G143), .B(KEYINPUT115), .Z(n691) );
  XNOR2_X1 U748 ( .A(n692), .B(n691), .ZN(G45) );
  NOR2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U750 ( .A(KEYINPUT116), .B(n695), .Z(n696) );
  XNOR2_X1 U751 ( .A(G146), .B(n696), .ZN(G48) );
  NAND2_X1 U752 ( .A1(n700), .A2(n697), .ZN(n698) );
  XNOR2_X1 U753 ( .A(n698), .B(G113), .ZN(G15) );
  NAND2_X1 U754 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U755 ( .A(n701), .B(G116), .ZN(G18) );
  XOR2_X1 U756 ( .A(G125), .B(KEYINPUT37), .Z(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(G27) );
  XOR2_X1 U758 ( .A(G134), .B(n704), .Z(G36) );
  NAND2_X1 U759 ( .A1(n705), .A2(n724), .ZN(n709) );
  NAND2_X1 U760 ( .A1(G953), .A2(G224), .ZN(n706) );
  XNOR2_X1 U761 ( .A(KEYINPUT61), .B(n706), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n707), .A2(G898), .ZN(n708) );
  NAND2_X1 U763 ( .A1(n709), .A2(n708), .ZN(n718) );
  XOR2_X1 U764 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n712) );
  XNOR2_X1 U765 ( .A(G101), .B(n710), .ZN(n711) );
  XNOR2_X1 U766 ( .A(n712), .B(n711), .ZN(n713) );
  XOR2_X1 U767 ( .A(n714), .B(n713), .Z(n716) );
  NOR2_X1 U768 ( .A1(G898), .A2(n724), .ZN(n715) );
  NOR2_X1 U769 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(G69) );
  XNOR2_X1 U771 ( .A(n720), .B(n719), .ZN(n721) );
  XOR2_X1 U772 ( .A(n722), .B(n721), .Z(n726) );
  XOR2_X1 U773 ( .A(n726), .B(n723), .Z(n725) );
  NAND2_X1 U774 ( .A1(n725), .A2(n724), .ZN(n730) );
  XNOR2_X1 U775 ( .A(G227), .B(n726), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n727), .A2(G900), .ZN(n728) );
  NAND2_X1 U777 ( .A1(n728), .A2(G953), .ZN(n729) );
  NAND2_X1 U778 ( .A1(n730), .A2(n729), .ZN(G72) );
  XNOR2_X1 U779 ( .A(n731), .B(G131), .ZN(n732) );
  XNOR2_X1 U780 ( .A(n732), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U781 ( .A(n733), .B(G137), .Z(G39) );
  XOR2_X1 U782 ( .A(G140), .B(n734), .Z(G42) );
endmodule

