//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(G50), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n208), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  NAND3_X1  g0041(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(new_n209), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n202), .A2(G50), .ZN(new_n244));
  OR3_X1    g0044(.A1(new_n244), .A2(KEYINPUT68), .A3(new_n210), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n210), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G150), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT68), .B1(new_n244), .B2(new_n210), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n245), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G58), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n210), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n243), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n210), .A2(G1), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n243), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(new_n265), .B2(G50), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT65), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT65), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G274), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G226), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(new_n270), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n280), .B1(new_n281), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G1698), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G222), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G223), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(G1698), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n291), .B1(new_n215), .B2(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT66), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n277), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n294), .A2(new_n293), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n298), .B1(G77), .B2(new_n289), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n299), .A2(KEYINPUT66), .A3(new_n291), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n285), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n267), .B1(new_n301), .B2(G169), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(new_n301), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n304), .A2(KEYINPUT70), .A3(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(KEYINPUT69), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT70), .B1(new_n304), .B2(G179), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n303), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT73), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n301), .A2(new_n311), .A3(G190), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n260), .A2(KEYINPUT9), .A3(new_n266), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT72), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT9), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n304), .A2(G200), .B1(new_n316), .B2(new_n267), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n313), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n317), .A2(new_n315), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n313), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n308), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G68), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G20), .ZN(new_n325));
  INV_X1    g0125(.A(G50), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n325), .B1(new_n258), .B2(new_n215), .C1(new_n326), .C2(new_n247), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n243), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT11), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n262), .A2(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT12), .B1(new_n333), .B2(G68), .ZN(new_n334));
  INV_X1    g0134(.A(G13), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(G1), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT12), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n334), .B1(new_n325), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT71), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n336), .B2(G20), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n330), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n243), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n264), .A2(new_n324), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n343), .A2(KEYINPUT75), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT75), .B1(new_n343), .B2(new_n344), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n329), .B(new_n339), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT74), .ZN(new_n348));
  INV_X1    g0148(.A(G232), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n294), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n292), .A2(KEYINPUT74), .A3(G232), .A4(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G97), .ZN(new_n353));
  INV_X1    g0153(.A(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n292), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n353), .B1(new_n355), .B2(new_n281), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n277), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G238), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n280), .B1(new_n359), .B2(new_n284), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT13), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n278), .B1(new_n274), .B2(new_n271), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(G238), .B2(new_n283), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n356), .B1(new_n350), .B2(new_n351), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n362), .B(new_n364), .C1(new_n365), .C2(new_n277), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G169), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n368), .A2(KEYINPUT14), .B1(new_n369), .B2(new_n367), .ZN(new_n370));
  INV_X1    g0170(.A(G169), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n371), .B1(new_n361), .B2(new_n366), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT14), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n347), .B1(new_n370), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n347), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n361), .A2(G190), .A3(new_n366), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n361), .B2(new_n366), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT76), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n380), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n377), .A4(new_n376), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n343), .B(G77), .C1(G1), .C2(new_n210), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n342), .A2(new_n215), .ZN(new_n387));
  INV_X1    g0187(.A(new_n243), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n252), .A2(new_n247), .B1(new_n210), .B2(new_n215), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n246), .A2(G20), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n292), .A2(G238), .A3(G1698), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n395), .B1(new_n217), .B2(new_n292), .C1(new_n355), .C2(new_n349), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n282), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n363), .B1(G244), .B2(new_n283), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n371), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n394), .B(new_n400), .C1(G179), .C2(new_n399), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n394), .B1(G200), .B2(new_n399), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n397), .A2(G190), .A3(new_n398), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n375), .A2(new_n385), .A3(new_n401), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n287), .A2(KEYINPUT77), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT77), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT3), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n408), .A3(G33), .ZN(new_n409));
  AOI21_X1  g0209(.A(G20), .B1(new_n409), .B2(new_n286), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT7), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n324), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n286), .ZN(new_n413));
  XNOR2_X1  g0213(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(G33), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT7), .B1(new_n415), .B2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n255), .A2(new_n324), .ZN(new_n418));
  OAI21_X1  g0218(.A(G20), .B1(new_n418), .B2(new_n201), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n248), .A2(G159), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT16), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n411), .A2(G20), .ZN(new_n425));
  AOI21_X1  g0225(.A(G33), .B1(new_n406), .B2(new_n408), .ZN(new_n426));
  INV_X1    g0226(.A(new_n288), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n411), .B1(new_n292), .B2(G20), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n324), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n424), .B1(new_n430), .B2(new_n421), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n431), .A3(new_n243), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n283), .A2(G232), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n280), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(G223), .A2(G1698), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n281), .B2(G1698), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n409), .A3(new_n286), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G33), .A2(G87), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n277), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G200), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n275), .A2(new_n279), .B1(new_n283), .B2(G232), .ZN(new_n441));
  AND2_X1   g0241(.A1(new_n437), .A2(new_n438), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n441), .B(G190), .C1(new_n442), .C2(new_n277), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n257), .A2(new_n265), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n262), .B2(new_n257), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n432), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n421), .B1(new_n412), .B2(new_n416), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n388), .B1(new_n451), .B2(KEYINPUT16), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n446), .B1(new_n452), .B2(new_n431), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(KEYINPUT17), .A3(new_n444), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(KEYINPUT78), .A2(KEYINPUT18), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n432), .A2(new_n447), .ZN(new_n458));
  OAI21_X1  g0258(.A(G169), .B1(new_n434), .B2(new_n439), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n441), .B(G179), .C1(new_n442), .C2(new_n277), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n461), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n453), .A2(new_n464), .A3(KEYINPUT18), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT18), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(new_n458), .B2(new_n461), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT78), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g0269(.A1(new_n323), .A2(new_n405), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OR3_X1    g0271(.A1(new_n262), .A2(KEYINPUT25), .A3(G107), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT25), .B1(new_n262), .B2(G107), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n261), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n262), .A2(new_n474), .A3(new_n209), .A4(new_n242), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n472), .B(new_n473), .C1(new_n217), .C2(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT89), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT5), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT81), .B1(new_n479), .B2(G41), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n268), .A3(KEYINPUT5), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n261), .B(G45), .C1(new_n268), .C2(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n282), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G264), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n484), .B1(new_n480), .B2(new_n482), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n279), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n409), .A2(G250), .A3(new_n354), .A4(new_n286), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G294), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n415), .A2(KEYINPUT90), .A3(G257), .A4(G1698), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT90), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n409), .A2(new_n286), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G257), .A2(G1698), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n492), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n487), .B(new_n489), .C1(new_n498), .C2(new_n277), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(new_n379), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n500), .B1(G190), .B2(new_n499), .ZN(new_n501));
  OR3_X1    g0301(.A1(new_n210), .A2(KEYINPUT23), .A3(G107), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(KEYINPUT88), .B1(KEYINPUT23), .B2(G107), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n502), .A2(KEYINPUT88), .B1(new_n505), .B2(G20), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(G87), .ZN(new_n509));
  NOR4_X1   g0309(.A1(new_n289), .A2(KEYINPUT22), .A3(G20), .A4(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT86), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n415), .A2(new_n511), .A3(new_n210), .A4(G87), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n409), .A2(new_n210), .A3(G87), .A4(new_n286), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT86), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT22), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT87), .A4(KEYINPUT22), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n508), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n243), .B1(new_n519), .B2(KEYINPUT24), .ZN(new_n520));
  INV_X1    g0320(.A(new_n514), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT22), .B1(new_n513), .B2(KEYINPUT86), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n510), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(KEYINPUT24), .A3(new_n507), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n478), .B(new_n501), .C1(new_n520), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n507), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n388), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n477), .B1(new_n531), .B2(new_n526), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n499), .A2(G179), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n499), .A2(new_n371), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n528), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n217), .B1(new_n428), .B2(new_n429), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT6), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n542), .A2(new_n210), .B1(new_n215), .B2(new_n247), .ZN(new_n543));
  OAI211_X1 g0343(.A(KEYINPUT79), .B(new_n243), .C1(new_n537), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n475), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n262), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(G97), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT80), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n545), .B(new_n549), .C1(G97), .C2(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n540), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n538), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(G20), .B1(G77), .B2(new_n248), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n288), .B1(new_n414), .B2(G33), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n289), .A2(new_n210), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n425), .B1(new_n559), .B2(new_n411), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n560), .B2(new_n217), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT79), .B1(new_n561), .B2(new_n243), .ZN(new_n562));
  OR2_X1    g0362(.A1(new_n552), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n409), .A2(G244), .A3(new_n354), .A4(new_n286), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT4), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g0366(.A1(KEYINPUT4), .A2(G244), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n286), .A2(new_n288), .A3(new_n567), .A4(new_n354), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n286), .A2(new_n288), .A3(G250), .A4(G1698), .ZN(new_n569));
  NAND2_X1  g0369(.A1(G33), .A2(G283), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n282), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n480), .A2(new_n482), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(new_n277), .C1(new_n574), .C2(new_n484), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n489), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT82), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n575), .A2(new_n578), .A3(new_n489), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n371), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n575), .A2(new_n578), .A3(new_n489), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n277), .B1(new_n566), .B2(new_n571), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n578), .B1(new_n575), .B2(new_n489), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n369), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n563), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n486), .A2(G270), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n489), .ZN(new_n589));
  NOR2_X1   g0389(.A1(G257), .A2(G1698), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n218), .B2(G1698), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(new_n409), .A3(new_n286), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n289), .A2(G303), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n277), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n593), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n282), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n486), .A2(G270), .B1(new_n279), .B2(new_n488), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n598), .A3(G190), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n331), .A2(new_n600), .A3(new_n332), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n261), .B2(G33), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n388), .B(new_n602), .C1(new_n341), .C2(new_n330), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n242), .A2(new_n209), .B1(G20), .B2(new_n600), .ZN(new_n604));
  INV_X1    g0404(.A(G97), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n570), .B(new_n210), .C1(G33), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT20), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n604), .A2(KEYINPUT20), .A3(new_n606), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n601), .B(new_n603), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n595), .A2(new_n599), .A3(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n609), .B(G169), .C1(new_n589), .C2(new_n594), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n589), .A2(new_n594), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(G179), .A3(new_n609), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n597), .A2(new_n598), .ZN(new_n618));
  INV_X1    g0418(.A(new_n614), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(G169), .A3(new_n619), .A4(new_n609), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n611), .A2(new_n615), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n391), .B(KEYINPUT84), .ZN(new_n622));
  INV_X1    g0422(.A(new_n475), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n333), .A2(new_n392), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n415), .A2(new_n210), .A3(G68), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT19), .B1(new_n390), .B2(G97), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT19), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n210), .B1(new_n353), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n554), .A2(new_n509), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n624), .B(new_n626), .C1(new_n633), .C2(new_n388), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n277), .B(G250), .C1(G1), .C2(new_n269), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n277), .A2(new_n261), .A3(G45), .A4(G274), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(G238), .A2(G1698), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n216), .B2(G1698), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n415), .A2(new_n640), .B1(G33), .B2(G116), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n638), .B1(new_n641), .B2(new_n277), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n371), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n638), .B(new_n369), .C1(new_n641), .C2(new_n277), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n634), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n388), .B1(new_n627), .B2(new_n632), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n475), .A2(new_n509), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n646), .A2(new_n625), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(G200), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n638), .B(G190), .C1(new_n641), .C2(new_n277), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n621), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n573), .A2(new_n577), .A3(new_n309), .A4(new_n579), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n585), .B2(G200), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT83), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n552), .A2(new_n562), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n656), .B1(new_n655), .B2(new_n657), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n587), .B(new_n653), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n471), .A2(new_n536), .A3(new_n660), .ZN(G372));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n587), .B2(new_n652), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n637), .A2(KEYINPUT91), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT91), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n664), .B1(new_n635), .B2(new_n636), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n663), .A2(new_n665), .B1(new_n641), .B2(new_n277), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n371), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n634), .A3(new_n644), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(G200), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n648), .A3(new_n650), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n586), .A2(new_n581), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT26), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .A4(new_n563), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n662), .A2(new_n675), .A3(new_n668), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n582), .A2(new_n584), .ZN(new_n677));
  AOI21_X1  g0477(.A(G200), .B1(new_n677), .B2(new_n573), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n309), .A2(new_n573), .A3(new_n577), .A4(new_n579), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n657), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT83), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n528), .A3(new_n587), .A4(new_n672), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n529), .A2(new_n530), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n685), .A2(new_n243), .A3(new_n526), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n535), .B1(new_n686), .B2(new_n478), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n615), .A2(new_n617), .A3(new_n620), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n676), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n470), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n308), .ZN(new_n692));
  INV_X1    g0492(.A(new_n467), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n458), .A2(new_n466), .A3(new_n461), .ZN(new_n694));
  INV_X1    g0494(.A(new_n367), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n695), .A2(G179), .B1(new_n372), .B2(new_n373), .ZN(new_n696));
  INV_X1    g0496(.A(new_n374), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n376), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT92), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n401), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n401), .A2(new_n699), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n698), .B1(new_n385), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(new_n693), .B(new_n694), .C1(new_n703), .C2(new_n455), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n318), .A2(KEYINPUT10), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n321), .A2(new_n320), .A3(new_n313), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n692), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n691), .A2(new_n708), .ZN(G369));
  INV_X1    g0509(.A(new_n687), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n336), .A2(new_n210), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(KEYINPUT27), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(G213), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(G343), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n532), .A2(new_n717), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n710), .A2(new_n717), .B1(new_n536), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n717), .A2(new_n610), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n688), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n621), .B2(new_n720), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G330), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n687), .A2(new_n717), .ZN(new_n726));
  INV_X1    g0526(.A(new_n536), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n688), .A2(new_n717), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n725), .A2(new_n726), .A3(new_n729), .ZN(G399));
  INV_X1    g0530(.A(new_n206), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n631), .A2(G116), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(G1), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(new_n213), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n690), .A2(new_n717), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT26), .B1(new_n587), .B2(new_n671), .ZN(new_n743));
  INV_X1    g0543(.A(new_n652), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n673), .A3(new_n674), .A4(new_n563), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n743), .A2(new_n745), .A3(new_n668), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n684), .B2(new_n689), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(KEYINPUT29), .A3(new_n717), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n738), .A2(KEYINPUT95), .A3(new_n739), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n742), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT93), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n487), .B1(new_n498), .B2(new_n277), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n618), .A2(new_n642), .A3(new_n369), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(new_n585), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT30), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n616), .A2(G179), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(new_n752), .A3(new_n642), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(KEYINPUT93), .A3(KEYINPUT30), .A4(new_n585), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  AND4_X1   g0561(.A1(new_n369), .A2(new_n580), .A3(new_n618), .A4(new_n666), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n762), .A2(new_n499), .B1(new_n755), .B2(new_n756), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT31), .B1(new_n764), .B2(new_n716), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT31), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n766), .B(new_n717), .C1(new_n761), .C2(new_n763), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT94), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n660), .A2(new_n716), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n727), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n683), .A2(new_n587), .A3(new_n653), .A4(new_n717), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n772), .A2(new_n536), .A3(KEYINPUT94), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n768), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G330), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n750), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n737), .B1(new_n778), .B2(G1), .ZN(G364));
  NOR2_X1   g0579(.A1(new_n722), .A2(G330), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT97), .Z(new_n781));
  NOR2_X1   g0581(.A1(new_n335), .A2(G20), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n261), .B1(new_n782), .B2(G45), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n732), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n781), .A2(new_n723), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n209), .B1(G20), .B2(new_n371), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n240), .A2(G45), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n415), .A2(new_n731), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n793), .B(new_n794), .C1(G45), .C2(new_n213), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n292), .A2(new_n206), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(G116), .B2(new_n206), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT98), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n792), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n210), .A2(new_n369), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G190), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n210), .A2(G179), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(new_n309), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n804), .A2(G68), .B1(new_n807), .B2(G107), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n309), .A2(G179), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n210), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G97), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n805), .A2(G190), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G87), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n808), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G190), .A2(G200), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n805), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT32), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n803), .A2(new_n309), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n820), .B1(new_n822), .B2(new_n326), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n818), .A2(KEYINPUT32), .A3(new_n819), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n802), .A2(new_n817), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n802), .A2(G190), .A3(new_n379), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n292), .B1(new_n825), .B2(new_n215), .C1(new_n255), .C2(new_n826), .ZN(new_n827));
  NOR4_X1   g0627(.A1(new_n816), .A2(new_n823), .A3(new_n824), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n826), .ZN(new_n829));
  INV_X1    g0629(.A(new_n818), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n829), .A2(G322), .B1(new_n830), .B2(G329), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n289), .C1(new_n832), .C2(new_n825), .ZN(new_n833));
  INV_X1    g0633(.A(G317), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(KEYINPUT33), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n834), .A2(KEYINPUT33), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n804), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n821), .A2(G326), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n837), .B(new_n838), .C1(new_n839), .C2(new_n810), .ZN(new_n840));
  INV_X1    g0640(.A(G283), .ZN(new_n841));
  INV_X1    g0641(.A(G303), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n806), .A2(new_n841), .B1(new_n813), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n833), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n828), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n786), .B(new_n801), .C1(new_n791), .C2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n790), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n722), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n787), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G396));
  NAND2_X1  g0650(.A1(new_n394), .A2(new_n716), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n404), .A2(new_n401), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT101), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n700), .A2(new_n394), .A3(new_n701), .A4(new_n716), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n404), .A2(new_n401), .A3(new_n855), .A4(new_n851), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n738), .B(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G330), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n770), .A2(new_n727), .A3(new_n769), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT94), .B1(new_n772), .B2(new_n536), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n862), .B2(new_n768), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n858), .A2(new_n863), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n785), .B(new_n864), .C1(KEYINPUT102), .C2(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(KEYINPUT102), .B2(new_n865), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n791), .A2(new_n788), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT99), .Z(new_n869));
  OAI21_X1  g0669(.A(new_n785), .B1(new_n869), .B2(G77), .ZN(new_n870));
  INV_X1    g0670(.A(new_n804), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n871), .A2(new_n841), .B1(new_n217), .B2(new_n813), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G87), .B2(new_n807), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n826), .A2(new_n839), .B1(new_n818), .B2(new_n832), .ZN(new_n874));
  INV_X1    g0674(.A(new_n825), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n292), .B(new_n874), .C1(G116), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n821), .A2(G303), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n873), .A2(new_n812), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n829), .A2(G143), .B1(new_n875), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n822), .B2(new_n880), .C1(new_n881), .C2(new_n871), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT34), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT100), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n807), .A2(G68), .ZN(new_n885));
  OAI221_X1 g0685(.A(new_n885), .B1(new_n326), .B2(new_n813), .C1(new_n255), .C2(new_n810), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n495), .B(new_n886), .C1(G132), .C2(new_n830), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n883), .A2(KEYINPUT100), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n870), .B1(new_n890), .B2(new_n791), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n857), .B2(new_n789), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n867), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(G384));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n448), .B1(new_n453), .B2(new_n464), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT107), .B1(new_n453), .B2(new_n714), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT107), .ZN(new_n898));
  INV_X1    g0698(.A(new_n714), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n458), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n896), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n902));
  INV_X1    g0702(.A(KEYINPUT106), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n451), .A2(KEYINPUT16), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n446), .B1(new_n904), .B2(new_n452), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n903), .B1(new_n905), .B2(new_n714), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n423), .A2(new_n243), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n451), .A2(KEYINPUT16), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n447), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT106), .A3(new_n899), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n461), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n906), .A2(new_n910), .A3(new_n448), .A4(new_n911), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n901), .A2(new_n902), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n906), .A2(new_n910), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n463), .B2(new_n468), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n895), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n901), .A2(new_n902), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n906), .A2(new_n910), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT78), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n693), .B2(new_n694), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n458), .A2(new_n461), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n456), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(new_n450), .A3(new_n454), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n920), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n926), .A3(KEYINPUT38), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n916), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n347), .A2(new_n716), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n929), .B(KEYINPUT105), .Z(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n381), .A2(new_n384), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n931), .B1(new_n932), .B2(new_n698), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n375), .A2(new_n385), .A3(new_n930), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n857), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n774), .A2(new_n928), .A3(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT109), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n941), .A3(new_n938), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n693), .A2(new_n694), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n900), .B(new_n897), .C1(new_n944), .C2(new_n455), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n901), .A2(new_n902), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n901), .A2(new_n902), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n895), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n938), .B1(new_n949), .B2(new_n927), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n935), .B1(new_n862), .B2(new_n768), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n943), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n470), .A2(new_n774), .ZN(new_n954));
  OAI21_X1  g0754(.A(G330), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n698), .A2(new_n717), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n916), .A2(new_n927), .A3(KEYINPUT39), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n948), .A2(new_n895), .ZN(new_n960));
  INV_X1    g0760(.A(new_n927), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n958), .B(new_n959), .C1(new_n962), .C2(KEYINPUT39), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n933), .A2(new_n934), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n690), .A2(new_n717), .A3(new_n857), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n401), .A2(new_n716), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT104), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n964), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n928), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n944), .A2(new_n714), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n963), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n742), .A2(new_n470), .A3(new_n748), .A4(new_n749), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n708), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n971), .B(new_n973), .Z(new_n974));
  NOR2_X1   g0774(.A1(new_n956), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n956), .A2(new_n974), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n261), .B2(new_n782), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n975), .B1(new_n977), .B2(KEYINPUT110), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(KEYINPUT110), .B2(new_n977), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n542), .B(KEYINPUT103), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT35), .ZN(new_n981));
  OAI211_X1 g0781(.A(G116), .B(new_n211), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(new_n981), .B2(new_n980), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT36), .Z(new_n984));
  NOR3_X1   g0784(.A1(new_n213), .A2(new_n215), .A3(new_n418), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n324), .A2(G50), .ZN(new_n986));
  OAI211_X1 g0786(.A(G1), .B(new_n335), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n979), .A2(new_n984), .A3(new_n987), .ZN(G367));
  OAI21_X1  g0788(.A(new_n729), .B1(new_n719), .B2(new_n728), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n723), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n729), .A2(new_n726), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n683), .B(new_n587), .C1(new_n657), .C2(new_n717), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n673), .A2(new_n563), .A3(new_n716), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT44), .Z(new_n998));
  NOR2_X1   g0798(.A1(new_n992), .A2(new_n996), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(new_n725), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n777), .B1(new_n991), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n732), .B(KEYINPUT41), .Z(new_n1004));
  OAI21_X1  g0804(.A(new_n783), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n995), .A2(new_n727), .A3(new_n728), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n683), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n587), .B1(new_n710), .B2(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1006), .A2(KEYINPUT42), .B1(new_n717), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(KEYINPUT42), .B2(new_n1006), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT43), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n648), .A2(new_n717), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n672), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n1012), .A2(new_n668), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1010), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1011), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1017), .B(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n725), .A2(new_n996), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1005), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1016), .A2(new_n790), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n794), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n792), .B1(new_n206), .B2(new_n391), .C1(new_n1025), .C2(new_n232), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n785), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n826), .A2(new_n881), .B1(new_n825), .B2(new_n326), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n289), .B(new_n1028), .C1(G137), .C2(new_n830), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n813), .A2(new_n255), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n810), .A2(new_n324), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(G159), .C2(new_n804), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n806), .A2(new_n215), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G143), .B2(new_n821), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1029), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n822), .A2(new_n832), .B1(new_n217), .B2(new_n810), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G294), .B2(new_n804), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n826), .A2(new_n842), .B1(new_n825), .B2(new_n841), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G317), .B2(new_n830), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n415), .B1(G97), .B2(new_n807), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n813), .A2(new_n600), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT46), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1035), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1027), .B1(new_n1045), .B2(new_n791), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1024), .A2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1023), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(G387));
  NOR2_X1   g0849(.A1(new_n777), .A2(new_n990), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(new_n733), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n778), .B2(new_n991), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n719), .A2(new_n847), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n252), .A2(G50), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT50), .ZN(new_n1055));
  AOI21_X1  g0855(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n734), .A3(new_n1056), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1057), .B(new_n794), .C1(new_n229), .C2(new_n269), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n797), .A2(new_n734), .B1(G107), .B2(new_n206), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT111), .Z(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(KEYINPUT112), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n792), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT112), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n785), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n829), .A2(G317), .B1(new_n875), .B2(G303), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n821), .A2(G322), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(new_n832), .C2(new_n871), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n841), .B2(new_n810), .C1(new_n839), .C2(new_n813), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1072), .A2(KEYINPUT49), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n806), .A2(new_n600), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n415), .B(new_n1075), .C1(G326), .C2(new_n830), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n822), .A2(new_n819), .B1(new_n813), .B2(new_n215), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n495), .B(new_n1078), .C1(G97), .C2(new_n807), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n257), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n804), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n622), .A2(new_n811), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n825), .A2(new_n324), .B1(new_n818), .B2(new_n881), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G50), .B2(new_n829), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1077), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1064), .B1(new_n1086), .B2(new_n791), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n991), .A2(new_n784), .B1(new_n1053), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1052), .A2(new_n1088), .ZN(G393));
  NOR2_X1   g0889(.A1(new_n1050), .A2(new_n1002), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT113), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n733), .B1(new_n1050), .B2(new_n1002), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n996), .A2(new_n790), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n237), .A2(new_n1025), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n792), .B1(new_n605), .B2(new_n206), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n785), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n822), .A2(new_n881), .B1(new_n819), .B2(new_n826), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n825), .A2(new_n252), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n495), .B(new_n1100), .C1(G143), .C2(new_n830), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n810), .A2(new_n215), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n806), .A2(new_n509), .B1(new_n813), .B2(new_n324), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(G50), .C2(new_n804), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G317), .A2(new_n821), .B1(new_n829), .B2(G311), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n871), .A2(new_n842), .B1(new_n600), .B2(new_n810), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n292), .B1(new_n830), .B2(G322), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n839), .B2(new_n825), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n806), .A2(new_n217), .B1(new_n813), .B2(new_n841), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1108), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1105), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1097), .B1(new_n1113), .B2(new_n791), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1002), .A2(new_n784), .B1(new_n1094), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1093), .A2(new_n1115), .ZN(G390));
  INV_X1    g0916(.A(new_n964), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n863), .A2(new_n857), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT39), .B1(new_n949), .B2(new_n927), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n959), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1120), .A2(new_n1121), .B1(new_n968), .B2(new_n958), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT115), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n747), .A2(new_n717), .A3(new_n857), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT114), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n967), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1124), .B2(new_n967), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n964), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1122), .B(new_n1123), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1124), .A2(new_n967), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(KEYINPUT114), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1124), .A2(new_n1125), .A3(new_n967), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1117), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1129), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1123), .B1(new_n1137), .B2(new_n1122), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1119), .B1(new_n1131), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1122), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT115), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1118), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n863), .A2(new_n470), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n972), .A2(new_n708), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n857), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n964), .B1(new_n775), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1118), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n965), .A2(new_n967), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1146), .B(new_n1118), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1144), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1139), .A2(new_n1142), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT116), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1151), .B(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1138), .A2(new_n1119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1141), .A2(new_n1130), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n1119), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n732), .B(new_n1152), .C1(new_n1154), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n784), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n788), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n785), .B1(new_n869), .B2(new_n1080), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n830), .A2(G125), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n289), .B(new_n1162), .C1(G132), .C2(new_n829), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(G159), .A2(new_n811), .B1(new_n821), .B2(G128), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT117), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n875), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n804), .A2(G137), .B1(new_n807), .B2(G50), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1163), .A2(new_n1164), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n813), .A2(new_n881), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1171));
  XNOR2_X1  g0971(.A(new_n1170), .B(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n826), .A2(new_n600), .B1(new_n818), .B2(new_n839), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n292), .B(new_n1173), .C1(G97), .C2(new_n875), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n815), .A3(new_n885), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1102), .B1(G283), .B2(new_n821), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n217), .B2(new_n871), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1169), .A2(new_n1172), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1161), .B1(new_n1178), .B2(new_n791), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1160), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1158), .A2(new_n1159), .A3(new_n1180), .ZN(G378));
  XOR2_X1   g0981(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n267), .A2(new_n899), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT120), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n707), .A2(new_n308), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n707), .B2(new_n308), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1183), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1189), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n1187), .A3(new_n1182), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n788), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n415), .A2(G41), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G50), .B(new_n1195), .C1(new_n246), .C2(new_n268), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n871), .A2(new_n605), .B1(new_n822), .B2(new_n600), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n806), .A2(new_n255), .B1(new_n813), .B2(new_n215), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n622), .A2(new_n875), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n826), .A2(new_n217), .B1(new_n818), .B2(new_n841), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1201), .A2(new_n1031), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1195), .A4(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT58), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1196), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(G128), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n826), .A2(new_n1206), .B1(new_n825), .B2(new_n880), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G132), .B2(new_n804), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1166), .A2(new_n814), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G150), .A2(new_n811), .B1(new_n821), .B2(G125), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n807), .A2(G159), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n830), .C2(G124), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1205), .B1(new_n1204), .B2(new_n1203), .C1(new_n1212), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n791), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT119), .Z(new_n1219));
  AOI211_X1 g1019(.A(new_n786), .B(new_n1219), .C1(new_n326), .C2(new_n868), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1194), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT121), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n859), .B1(new_n950), .B2(new_n951), .ZN(new_n1224));
  AOI211_X1 g1024(.A(KEYINPUT109), .B(KEYINPUT40), .C1(new_n951), .C2(new_n928), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n941), .B1(new_n937), .B2(new_n938), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1193), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1193), .B(new_n1224), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1223), .B(new_n971), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1229), .A2(new_n971), .A3(new_n1230), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n971), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1231), .B1(new_n1234), .B2(new_n1223), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1222), .B1(new_n1235), .B2(new_n784), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1144), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1152), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1144), .B1(new_n1157), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n971), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1193), .B1(new_n943), .B2(new_n1224), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1230), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1229), .A2(new_n971), .A3(new_n1230), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT57), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n732), .B1(new_n1241), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1236), .B1(new_n1239), .B2(new_n1249), .ZN(G375));
  INV_X1    g1050(.A(new_n791), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n826), .A2(new_n841), .B1(new_n825), .B2(new_n217), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n292), .B(new_n1252), .C1(G303), .C2(new_n830), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1033), .B1(G116), .B2(new_n804), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n821), .A2(G294), .B1(new_n814), .B2(G97), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1082), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n810), .A2(new_n326), .B1(new_n813), .B2(new_n819), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G132), .B2(new_n821), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1166), .A2(new_n804), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n825), .A2(new_n881), .B1(new_n818), .B2(new_n1206), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(G137), .B2(new_n829), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n495), .B1(G58), .B2(new_n807), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1259), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1251), .B1(new_n1256), .B2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n785), .B1(new_n869), .B2(G68), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n964), .C2(new_n788), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(new_n1240), .B2(new_n784), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1149), .A2(new_n1144), .A3(new_n1150), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1004), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1267), .B1(new_n1154), .B2(new_n1270), .ZN(G381));
  OR4_X1    g1071(.A1(G396), .A2(G393), .A3(G384), .A4(G381), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1272), .A2(G390), .A3(G387), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1180), .B1(new_n1274), .B2(new_n783), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1151), .B(KEYINPUT116), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n733), .B1(new_n1276), .B2(new_n1274), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1275), .B1(new_n1277), .B2(new_n1152), .ZN(new_n1278));
  INV_X1    g1078(.A(G375), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1273), .A2(new_n1278), .A3(new_n1279), .ZN(G407));
  NAND2_X1  g1080(.A1(new_n715), .A2(G213), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT122), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1279), .A2(new_n1278), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G407), .A2(G213), .A3(new_n1283), .ZN(G409));
  XNOR2_X1  g1084(.A(G393), .B(new_n849), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(G390), .A2(new_n1048), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(G390), .A2(new_n1048), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1286), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n1287), .A3(new_n1285), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1236), .C1(new_n1239), .C2(new_n1249), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1233), .A2(KEYINPUT121), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1245), .A2(new_n1223), .A3(new_n1246), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1238), .A2(new_n1269), .A3(new_n1295), .A4(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1222), .B1(new_n1247), .B2(new_n784), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT123), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1278), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1294), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1300), .B1(new_n1299), .B2(new_n1278), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1268), .B1(new_n1151), .B2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1149), .A2(KEYINPUT60), .A3(new_n1150), .A4(new_n1144), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n732), .A3(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(G384), .A2(new_n1309), .A3(new_n1267), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1267), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n893), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NOR4_X1   g1113(.A1(new_n1304), .A2(new_n1305), .A3(new_n1282), .A4(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1313), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1281), .B(new_n1315), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1305), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1316), .A2(KEYINPUT126), .A3(new_n1305), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1314), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  XOR2_X1   g1121(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1322));
  INV_X1    g1122(.A(new_n1281), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(G2897), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1315), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT124), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1313), .A2(G2897), .A3(new_n1282), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1325), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1304), .A2(new_n1282), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1322), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1293), .B1(new_n1321), .B2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1293), .A2(KEYINPUT61), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1316), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1331), .A2(KEYINPUT63), .A3(new_n1315), .ZN(new_n1337));
  OAI22_X1  g1137(.A1(new_n1328), .A2(new_n1329), .B1(new_n1304), .B2(new_n1323), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1334), .A2(new_n1336), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1333), .A2(new_n1339), .ZN(G405));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1290), .A2(new_n1292), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G375), .A2(new_n1278), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1343), .A2(new_n1294), .A3(new_n1313), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1294), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1315), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1342), .A2(new_n1344), .A3(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(KEYINPUT127), .A3(new_n1293), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1293), .A2(KEYINPUT127), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1349), .A2(new_n1344), .A3(new_n1346), .A4(new_n1342), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1348), .A2(new_n1350), .ZN(G402));
endmodule


