//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT65), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(new_n202), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g0018(.A(KEYINPUT66), .B(G238), .Z(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G87), .A2(G250), .ZN(new_n225));
  NAND4_X1  g0025(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n208), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n211), .B(new_n218), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G68), .B(G77), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n216), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n216), .A2(new_n252), .A3(KEYINPUT68), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G20), .B2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n249), .A2(new_n251), .B1(new_n256), .B2(G150), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(new_n204), .B2(new_n216), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n215), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n260), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n265), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(G50), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n268), .A2(new_n269), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n216), .A2(G1), .ZN(new_n273));
  NOR3_X1   g0073(.A1(new_n272), .A2(new_n260), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n271), .B1(new_n274), .B2(G50), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n263), .A2(new_n264), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  AND2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  OAI21_X1  g0082(.A(KEYINPUT67), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n252), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n288), .A3(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n283), .A2(G223), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(G1698), .B1(new_n285), .B2(new_n286), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n291), .A2(G222), .B1(new_n281), .B2(G77), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n278), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  AND2_X1   g0094(.A1(G1), .A2(G13), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(new_n277), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G226), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n278), .A2(new_n297), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n276), .B1(G169), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT10), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n264), .A2(new_n275), .ZN(new_n311));
  AOI21_X1  g0111(.A(KEYINPUT69), .B1(new_n258), .B2(new_n260), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT9), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT9), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n263), .A2(new_n314), .A3(new_n264), .A4(new_n275), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n303), .A2(G190), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n303), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n310), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  AOI211_X1 g0121(.A(KEYINPUT10), .B(new_n319), .C1(new_n313), .C2(new_n315), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n309), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n285), .A2(new_n216), .A3(new_n286), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT7), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n216), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n220), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(G58), .B(G68), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G20), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n253), .A2(new_n255), .ZN(new_n332));
  INV_X1    g0132(.A(G159), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n324), .B1(new_n329), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT7), .B1(new_n281), .B2(new_n216), .ZN(new_n336));
  NOR4_X1   g0136(.A1(new_n279), .A2(new_n280), .A3(new_n326), .A4(G20), .ZN(new_n337));
  OAI21_X1  g0137(.A(G68), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n256), .A2(G159), .B1(new_n330), .B2(G20), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(KEYINPUT16), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n335), .A2(new_n340), .A3(new_n260), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n270), .A2(new_n249), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n260), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n270), .B(new_n344), .C1(G1), .C2(new_n216), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n343), .B1(new_n345), .B2(new_n248), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n299), .B1(new_n233), .B2(new_n301), .ZN(new_n349));
  OR2_X1    g0149(.A1(G223), .A2(G1698), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n300), .A2(G1698), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n350), .B(new_n351), .C1(new_n279), .C2(new_n280), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G87), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT74), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n278), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n357));
  AOI211_X1 g0157(.A(new_n306), .B(new_n349), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n354), .A2(new_n355), .ZN(new_n360));
  INV_X1    g0160(.A(new_n278), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n349), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n358), .A2(new_n364), .A3(KEYINPUT75), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n352), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n367));
  AOI21_X1  g0167(.A(KEYINPUT74), .B1(new_n352), .B2(new_n353), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n367), .A2(new_n368), .A3(new_n278), .ZN(new_n369));
  OAI21_X1  g0169(.A(G169), .B1(new_n369), .B2(new_n349), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n362), .A2(G179), .A3(new_n363), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n348), .B1(new_n365), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT18), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n338), .A2(new_n339), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n344), .B1(new_n376), .B2(new_n324), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n346), .B1(new_n377), .B2(new_n340), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT75), .B1(new_n358), .B2(new_n364), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n366), .A3(new_n371), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT18), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n375), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n318), .B1(new_n369), .B2(new_n349), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n362), .A2(new_n385), .A3(new_n363), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT17), .B1(new_n378), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  AOI211_X1 g0189(.A(G190), .B(new_n349), .C1(new_n356), .C2(new_n357), .ZN(new_n390));
  AOI21_X1  g0190(.A(G200), .B1(new_n362), .B2(new_n363), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(new_n348), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n378), .A2(KEYINPUT76), .A3(new_n387), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n388), .B1(new_n395), .B2(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n383), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT15), .B(G87), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n332), .B2(new_n248), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(new_n260), .B1(new_n274), .B2(G77), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n272), .A2(new_n205), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT72), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n219), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n283), .A2(new_n406), .A3(new_n289), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n291), .A2(G232), .B1(new_n281), .B2(G107), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n278), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G244), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n299), .B1(new_n410), .B2(new_n301), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n405), .B1(G190), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n318), .B2(new_n412), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n306), .A2(new_n412), .B1(new_n402), .B2(new_n404), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n359), .B1(new_n409), .B2(new_n411), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT73), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n414), .A2(KEYINPUT73), .A3(new_n417), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n332), .A2(new_n240), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n250), .A2(new_n205), .B1(new_n216), .B2(G68), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n260), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT11), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n425), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT12), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n270), .A2(new_n428), .A3(G68), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n428), .B2(new_n270), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n220), .B1(new_n345), .B2(KEYINPUT12), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n233), .A2(G1698), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n287), .B(new_n435), .C1(G226), .C2(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G97), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n278), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G238), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n299), .B1(new_n439), .B2(new_n301), .ZN(new_n440));
  OR3_X1    g0240(.A1(new_n438), .A2(KEYINPUT13), .A3(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT13), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(G169), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(G179), .A3(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n443), .B2(G169), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n434), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n443), .A2(G200), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n433), .B(new_n450), .C1(new_n385), .C2(new_n443), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n420), .A2(new_n421), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n323), .A2(new_n397), .A3(new_n452), .ZN(new_n453));
  AND2_X1   g0253(.A1(KEYINPUT4), .A2(G244), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n282), .B(new_n454), .C1(new_n279), .C2(new_n280), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G33), .A2(G283), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n410), .B1(new_n285), .B2(new_n286), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n455), .B(new_n456), .C1(new_n457), .C2(KEYINPUT4), .ZN(new_n458));
  OAI21_X1  g0258(.A(G250), .B1(new_n279), .B2(new_n280), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n282), .B1(new_n459), .B2(KEYINPUT4), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n361), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(G41), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n265), .B(G45), .C1(new_n462), .C2(KEYINPUT5), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT5), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n464), .A2(G41), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n296), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n464), .A2(G41), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n265), .A4(G45), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G257), .A3(new_n278), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n461), .A2(new_n306), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n461), .A2(new_n472), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n359), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT79), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT6), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT78), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT78), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT6), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(G97), .B(G107), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n482), .A3(new_n484), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G20), .ZN(new_n491));
  AOI21_X1  g0291(.A(KEYINPUT77), .B1(new_n256), .B2(G77), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT77), .ZN(new_n493));
  AOI211_X1 g0293(.A(new_n493), .B(new_n205), .C1(new_n253), .C2(new_n255), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(G107), .B1(new_n336), .B2(new_n337), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n491), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n497), .A2(new_n260), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n272), .A2(new_n476), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n265), .A2(G33), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n270), .A2(new_n344), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n476), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n473), .B(new_n475), .C1(new_n498), .C2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n461), .A2(new_n385), .A3(new_n472), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n467), .A2(new_n471), .ZN(new_n505));
  INV_X1    g0305(.A(G250), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n506), .B1(new_n285), .B2(new_n286), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT4), .ZN(new_n508));
  OAI21_X1  g0308(.A(G1698), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n456), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n291), .B2(new_n454), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n508), .B1(new_n281), .B2(new_n410), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n505), .B1(new_n513), .B2(new_n361), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n504), .B1(new_n514), .B2(G200), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n502), .B1(new_n497), .B2(new_n260), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(KEYINPUT80), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT80), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n503), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G45), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n506), .B1(new_n520), .B2(G1), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n265), .A2(new_n294), .A3(G45), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n278), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G116), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n252), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G244), .A2(G1698), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n439), .B2(G1698), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n525), .B1(new_n287), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n306), .B(new_n523), .C1(new_n528), .C2(new_n278), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT81), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n439), .A2(G1698), .ZN(new_n532));
  AND2_X1   g0332(.A1(G244), .A2(G1698), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n532), .A2(new_n533), .B1(new_n279), .B2(new_n280), .ZN(new_n534));
  INV_X1    g0334(.A(new_n525), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n361), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n537), .A2(KEYINPUT81), .A3(new_n306), .A4(new_n523), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  XNOR2_X1  g0340(.A(KEYINPUT79), .B(G97), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n540), .B1(new_n541), .B2(new_n250), .ZN(new_n542));
  NOR2_X1   g0342(.A1(G87), .A2(G107), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n477), .A2(new_n479), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n216), .B1(new_n437), .B2(new_n540), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n287), .A2(new_n216), .A3(G68), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n260), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n272), .A2(new_n398), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n270), .A2(new_n344), .A3(new_n399), .A4(new_n500), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n523), .B1(new_n528), .B2(new_n278), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n359), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n539), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n548), .A2(new_n260), .B1(new_n272), .B2(new_n398), .ZN(new_n556));
  INV_X1    g0356(.A(G87), .ZN(new_n557));
  OR2_X1    g0357(.A1(new_n501), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n278), .A2(new_n521), .A3(new_n522), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n559), .B1(new_n536), .B2(new_n361), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n553), .A2(G190), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n556), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n555), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n555), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n519), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G257), .B(G1698), .C1(new_n279), .C2(new_n280), .ZN(new_n570));
  OAI211_X1 g0370(.A(G250), .B(new_n282), .C1(new_n279), .C2(new_n280), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n361), .ZN(new_n574));
  OAI211_X1 g0374(.A(G264), .B(new_n278), .C1(new_n463), .C2(new_n465), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n467), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G169), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT88), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n470), .A2(new_n579), .A3(G264), .A4(new_n278), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n573), .A2(new_n361), .B1(new_n296), .B2(new_n466), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(G179), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT24), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n216), .B(G87), .C1(new_n279), .C2(new_n280), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT22), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT22), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n287), .A2(new_n588), .A3(new_n216), .A4(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n216), .A2(G33), .A3(G116), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT23), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n486), .A3(G20), .ZN(new_n593));
  OAI21_X1  g0393(.A(KEYINPUT23), .B1(new_n216), .B2(G107), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT87), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n591), .B(new_n593), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n585), .B1(new_n590), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n590), .A2(new_n585), .A3(new_n598), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n344), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OR2_X1    g0402(.A1(new_n501), .A2(new_n486), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT25), .B1(new_n270), .B2(G107), .ZN(new_n604));
  OR3_X1    g0404(.A1(new_n270), .A2(KEYINPUT25), .A3(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n584), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n601), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n260), .B1(new_n608), .B2(new_n599), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n576), .A2(G190), .ZN(new_n611));
  AOI21_X1  g0411(.A(G200), .B1(new_n581), .B2(new_n582), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(G264), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G1698), .ZN(new_n616));
  OR2_X1    g0416(.A1(G257), .A2(G1698), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n616), .A2(new_n617), .B1(new_n285), .B2(new_n286), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n279), .A2(new_n280), .A3(G303), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT83), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT83), .ZN(new_n621));
  INV_X1    g0421(.A(G303), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n285), .A2(new_n622), .A3(new_n286), .ZN(new_n623));
  NOR2_X1   g0423(.A1(G257), .A2(G1698), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n615), .B2(G1698), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n621), .B(new_n623), .C1(new_n625), .C2(new_n281), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n620), .A2(new_n361), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n470), .A2(G270), .A3(new_n278), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n467), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n359), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n270), .A2(new_n344), .A3(G116), .A4(new_n500), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n272), .A2(new_n524), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n216), .B(new_n456), .C1(new_n541), .C2(G33), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n259), .A2(new_n215), .B1(G20), .B2(new_n524), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT20), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(G33), .B1(new_n477), .B2(new_n479), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n456), .A2(new_n216), .ZN(new_n637));
  OAI211_X1 g0437(.A(KEYINPUT20), .B(new_n634), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n631), .B(new_n632), .C1(new_n635), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT21), .B1(new_n641), .B2(KEYINPUT86), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT86), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n630), .A2(new_n643), .A3(new_n640), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n630), .A2(KEYINPUT21), .A3(new_n640), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n630), .A2(new_n640), .A3(KEYINPUT84), .A4(KEYINPUT21), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT85), .ZN(new_n651));
  INV_X1    g0451(.A(new_n640), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n627), .A2(G179), .A3(new_n629), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n627), .A2(G179), .A3(new_n629), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(KEYINPUT85), .A3(new_n640), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n627), .A2(new_n629), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n640), .B1(G200), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n385), .B2(new_n658), .ZN(new_n660));
  AND4_X1   g0460(.A1(new_n645), .A2(new_n650), .A3(new_n657), .A4(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n453), .A2(new_n569), .A3(new_n614), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT89), .Z(G372));
  OAI21_X1  g0463(.A(new_n348), .B1(new_n364), .B2(new_n358), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n451), .A2(new_n415), .A3(new_n416), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n449), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n665), .B1(new_n667), .B2(new_n396), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n321), .A2(new_n322), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n309), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT91), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(KEYINPUT91), .B(new_n309), .C1(new_n668), .C2(new_n669), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n475), .A2(new_n473), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n516), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n566), .A2(new_n567), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n552), .A2(new_n529), .A3(new_n554), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n563), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n680), .A2(new_n516), .A3(new_n674), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n677), .A2(KEYINPUT90), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n645), .A2(new_n650), .A3(new_n607), .A4(new_n657), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n515), .A2(new_n516), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT80), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n515), .A2(KEYINPUT80), .A3(new_n516), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n675), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n680), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(new_n613), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n685), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n684), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT90), .B1(new_n677), .B2(new_n683), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n672), .A2(new_n673), .B1(new_n453), .B2(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(new_n697), .B(KEYINPUT92), .Z(G369));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n265), .A2(new_n216), .A3(G13), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  XNOR2_X1  g0504(.A(KEYINPUT93), .B(G343), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n661), .B1(new_n652), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n648), .A2(new_n649), .B1(new_n654), .B2(new_n656), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n645), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n640), .A3(new_n706), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n699), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n706), .B1(new_n602), .B2(new_n606), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n614), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n607), .B2(new_n707), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n706), .B1(new_n709), .B2(new_n645), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n614), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n607), .B2(new_n706), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n716), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n209), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n265), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n541), .A2(new_n524), .A3(new_n543), .ZN(new_n726));
  INV_X1    g0526(.A(new_n723), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n725), .A2(new_n726), .B1(new_n213), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  AND4_X1   g0529(.A1(new_n560), .A2(new_n574), .A3(new_n578), .A4(new_n580), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n655), .A2(KEYINPUT30), .A3(new_n730), .A4(new_n514), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT94), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n560), .A2(new_n574), .A3(new_n578), .A4(new_n580), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n474), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT30), .A4(new_n655), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n730), .A2(new_n514), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n738), .B2(new_n653), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n581), .A2(new_n582), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n560), .A2(G179), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n740), .A2(new_n658), .A3(new_n474), .A4(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n732), .A2(new_n736), .A3(new_n739), .A4(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT31), .B1(new_n743), .B2(new_n706), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n569), .A2(new_n661), .A3(new_n614), .A4(new_n707), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n699), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n707), .B1(new_n694), .B2(new_n695), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT29), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT95), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n519), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(KEYINPUT95), .B(new_n503), .C1(new_n517), .C2(new_n518), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n753), .A2(new_n685), .A3(new_n692), .A4(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n566), .A2(new_n682), .A3(new_n567), .A4(new_n675), .ZN(new_n756));
  OAI21_X1  g0556(.A(KEYINPUT26), .B1(new_n503), .B2(new_n680), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n756), .A2(new_n678), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n706), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n748), .B1(new_n751), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n729), .B1(new_n761), .B2(G1), .ZN(G364));
  INV_X1    g0562(.A(new_n712), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n216), .A2(G13), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G45), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT96), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n725), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n708), .A2(new_n699), .A3(new_n711), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n763), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n708), .A2(new_n711), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n722), .A2(new_n281), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G355), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G116), .B2(new_n209), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n243), .A2(G45), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n722), .A2(new_n287), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n520), .B2(new_n214), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n777), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n215), .B1(G20), .B2(new_n359), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n773), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n767), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G179), .A2(G200), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n216), .B1(new_n787), .B2(G190), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n476), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT97), .B(G159), .Z(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n216), .A2(G190), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n787), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NAND3_X1  g0596(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n385), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n789), .B(new_n796), .C1(G50), .C2(new_n798), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n792), .A2(new_n306), .A3(G200), .ZN(new_n800));
  XOR2_X1   g0600(.A(new_n800), .B(KEYINPUT98), .Z(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n486), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n216), .A2(new_n385), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n306), .A2(G200), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n287), .B1(new_n806), .B2(new_n242), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n804), .A2(new_n306), .A3(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n792), .A2(new_n805), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n808), .A2(new_n557), .B1(new_n809), .B2(new_n205), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n803), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n797), .A2(G190), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(KEYINPUT99), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n799), .B(new_n811), .C1(new_n220), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n798), .ZN(new_n818));
  XOR2_X1   g0618(.A(KEYINPUT100), .B(G326), .Z(new_n819));
  INV_X1    g0619(.A(G294), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n818), .A2(new_n819), .B1(new_n820), .B2(new_n788), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT101), .Z(new_n822));
  NAND2_X1  g0622(.A1(new_n794), .A2(G329), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n823), .B1(new_n622), .B2(new_n808), .C1(new_n824), .C2(new_n809), .ZN(new_n825));
  INV_X1    g0625(.A(new_n806), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n287), .B(new_n825), .C1(G322), .C2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT33), .B(G317), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n815), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n801), .A2(G283), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n817), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n786), .B1(new_n832), .B2(new_n783), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n774), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n770), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G396));
  NOR2_X1   g0636(.A1(new_n418), .A2(new_n706), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n405), .A2(new_n706), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n414), .A2(new_n838), .B1(new_n416), .B2(new_n415), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n417), .A2(new_n706), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n696), .A2(new_n837), .B1(new_n749), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n767), .B1(new_n843), .B2(new_n748), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT103), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n748), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n845), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n842), .A2(new_n771), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n783), .A2(new_n771), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n767), .B1(G77), .B2(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT102), .Z(new_n854));
  OAI21_X1  g0654(.A(new_n281), .B1(new_n806), .B2(new_n820), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n789), .B(new_n855), .C1(G303), .C2(new_n798), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n801), .A2(G87), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n815), .A2(G283), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n809), .A2(new_n524), .B1(new_n793), .B2(new_n824), .ZN(new_n859));
  INV_X1    g0659(.A(new_n808), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(G107), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n856), .A2(new_n857), .A3(new_n858), .A4(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n809), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n863), .A2(new_n791), .B1(new_n826), .B2(G143), .ZN(new_n864));
  INV_X1    g0664(.A(G137), .ZN(new_n865));
  INV_X1    g0665(.A(G150), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n865), .B2(new_n818), .C1(new_n816), .C2(new_n866), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT34), .Z(new_n868));
  NAND2_X1  g0668(.A1(new_n801), .A2(G68), .ZN(new_n869));
  INV_X1    g0669(.A(G132), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n287), .B1(new_n793), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(G50), .B2(new_n860), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n869), .B(new_n872), .C1(new_n242), .C2(new_n788), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n862), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n854), .B1(new_n874), .B2(new_n783), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n848), .A2(new_n849), .B1(new_n850), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(G384));
  OR2_X1    g0677(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(G116), .A3(new_n217), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT36), .Z(new_n881));
  OAI211_X1 g0681(.A(new_n214), .B(G77), .C1(new_n242), .C2(new_n220), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n201), .A2(G68), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n265), .B(G13), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT104), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n434), .A2(new_n886), .A3(new_n706), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT104), .B1(new_n433), .B2(new_n707), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n449), .A2(new_n887), .A3(new_n451), .A4(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n434), .B(new_n706), .C1(new_n447), .C2(new_n448), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n837), .B1(new_n694), .B2(new_n695), .ZN(new_n893));
  INV_X1    g0693(.A(new_n840), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n393), .A2(new_n394), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT105), .B1(new_n348), .B2(new_n704), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT105), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n899), .B(new_n703), .C1(new_n341), .C2(new_n347), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n897), .A2(new_n664), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n348), .A2(new_n704), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n905));
  NOR3_X1   g0705(.A1(new_n381), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n902), .A2(KEYINPUT37), .B1(new_n897), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n901), .B1(new_n383), .B2(new_n396), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n896), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n898), .A2(new_n900), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n395), .A2(KEYINPUT17), .ZN(new_n911));
  INV_X1    g0711(.A(new_n388), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n374), .B(new_n378), .C1(new_n379), .C2(new_n380), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n379), .A2(new_n380), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT18), .B1(new_n915), .B2(new_n348), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n910), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n906), .A2(new_n897), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n393), .A2(new_n394), .A3(new_n664), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n910), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n918), .A2(KEYINPUT38), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n909), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n895), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n449), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n707), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n907), .A2(new_n908), .A3(new_n896), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT38), .B1(new_n918), .B2(new_n922), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT39), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n664), .B(new_n374), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n903), .B1(new_n396), .B2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n664), .B(new_n903), .C1(new_n348), .C2(new_n392), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n906), .A2(new_n897), .B1(new_n905), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n896), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n923), .A2(new_n931), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n927), .B1(new_n930), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n932), .A2(new_n704), .ZN(new_n939));
  OR3_X1    g0739(.A1(new_n925), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n453), .A2(new_n751), .A3(new_n760), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n672), .A2(new_n673), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n940), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n743), .A2(new_n706), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT31), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n555), .A2(KEYINPUT82), .A3(new_n563), .ZN(new_n950));
  AOI21_X1  g0750(.A(KEYINPUT82), .B1(new_n555), .B2(new_n563), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n690), .A2(new_n952), .A3(new_n707), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n614), .A2(new_n709), .A3(new_n645), .A4(new_n660), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n949), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n891), .A2(new_n841), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT40), .B1(new_n924), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n904), .B1(new_n913), .B2(new_n665), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n934), .A2(new_n905), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n919), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(KEYINPUT38), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT107), .B1(new_n928), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT107), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n923), .A2(new_n965), .A3(new_n936), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT40), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n956), .A2(new_n957), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n959), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n947), .B(new_n948), .C1(new_n954), .C2(new_n953), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n453), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(G330), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n970), .B1(new_n453), .B2(new_n971), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n944), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n265), .B2(new_n764), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n944), .A2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n885), .B1(new_n977), .B2(new_n978), .ZN(G367));
  NAND2_X1  g0779(.A1(new_n237), .A2(new_n779), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n785), .B1(new_n722), .B2(new_n399), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n768), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n773), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n707), .B1(new_n556), .B2(new_n558), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n679), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n680), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n808), .A2(new_n524), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n987), .A2(KEYINPUT46), .B1(new_n824), .B2(new_n818), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(KEYINPUT46), .B2(new_n987), .ZN(new_n989));
  INV_X1    g0789(.A(G283), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n809), .A2(new_n990), .B1(new_n788), .B2(new_n486), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT111), .Z(new_n992));
  INV_X1    g0792(.A(G317), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n800), .A2(new_n541), .B1(new_n793), .B2(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n287), .B(new_n994), .C1(G303), .C2(new_n826), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n815), .A2(G294), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n989), .A2(new_n992), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n788), .A2(new_n220), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G150), .B2(new_n826), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT112), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n287), .B1(new_n793), .B2(new_n865), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n808), .A2(new_n242), .B1(new_n800), .B2(new_n205), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(G143), .C2(new_n798), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n201), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n815), .A2(new_n791), .B1(new_n1004), .B2(new_n863), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT113), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1000), .B(new_n1003), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1005), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT113), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n997), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT47), .Z(new_n1011));
  INV_X1    g0811(.A(new_n783), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n982), .B1(new_n983), .B2(new_n986), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n766), .A2(new_n265), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n753), .B(new_n754), .C1(new_n516), .C2(new_n707), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n675), .A2(new_n706), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n719), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT44), .Z(new_n1021));
  NAND2_X1  g0821(.A1(new_n720), .A2(new_n1018), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT45), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1021), .A2(new_n1024), .A3(new_n716), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n716), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1020), .B(KEYINPUT44), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1026), .B1(new_n1027), .B2(new_n1023), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n718), .B1(new_n715), .B2(new_n717), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n712), .B(new_n1029), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1025), .A2(new_n761), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n761), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n723), .B(KEYINPUT41), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1015), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT108), .Z(new_n1036));
  NOR2_X1   g0836(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(KEYINPUT109), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1018), .A2(new_n614), .A3(new_n717), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT42), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n503), .B1(new_n1016), .B2(new_n607), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1041), .A2(new_n707), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1038), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n716), .A2(new_n1019), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT110), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1044), .B(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1048), .A2(new_n1049), .B1(KEYINPUT109), .B2(new_n1037), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1049), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1037), .A2(KEYINPUT109), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n1052), .A3(new_n1047), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1013), .B1(new_n1034), .B2(new_n1054), .ZN(G387));
  INV_X1    g0855(.A(new_n788), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n860), .A2(G294), .B1(new_n1056), .B2(G283), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n798), .A2(G322), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n809), .B2(new_n622), .C1(new_n993), .C2(new_n806), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G311), .B2(new_n815), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT114), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1057), .B1(new_n1062), .B2(KEYINPUT48), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT49), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n281), .B1(new_n800), .B2(new_n524), .C1(new_n819), .C2(new_n793), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n281), .B1(new_n863), .B2(G68), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n333), .B2(new_n818), .C1(new_n398), .C2(new_n788), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n860), .A2(G77), .B1(new_n794), .B2(G150), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n240), .B2(new_n806), .C1(new_n802), .C2(new_n476), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n249), .C2(new_n815), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n783), .B1(new_n1067), .B2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n715), .A2(new_n983), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n780), .B1(new_n234), .B2(G45), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n726), .B2(new_n775), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n249), .A2(new_n240), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT50), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n520), .B1(new_n220), .B2(new_n205), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1078), .A2(new_n726), .A3(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1076), .A2(new_n1080), .B1(G107), .B2(new_n209), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n768), .B(new_n1074), .C1(new_n784), .C2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1073), .A2(new_n1082), .B1(new_n1030), .B2(new_n1015), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n761), .A2(new_n1030), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n723), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n761), .A2(new_n1030), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(G393));
  NAND2_X1  g0887(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1084), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n723), .A3(new_n1031), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1025), .A2(new_n1028), .A3(new_n1015), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n784), .B1(new_n209), .B2(new_n541), .C1(new_n246), .C2(new_n780), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n767), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n287), .B1(new_n794), .B2(G322), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n990), .B2(new_n808), .C1(new_n820), .C2(new_n809), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1095), .B(new_n803), .C1(G116), .C2(new_n1056), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n818), .A2(new_n993), .B1(new_n806), .B2(new_n824), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(new_n622), .C2(new_n816), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT115), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n818), .A2(new_n866), .B1(new_n806), .B2(new_n333), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT51), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n815), .A2(new_n1004), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n808), .A2(new_n220), .B1(new_n809), .B2(new_n248), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n788), .A2(new_n205), .ZN(new_n1106));
  INV_X1    g0906(.A(G143), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n287), .B1(new_n793), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1105), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1103), .A2(new_n857), .A3(new_n1104), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1101), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1093), .B1(new_n1112), .B2(new_n783), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n1018), .B2(new_n983), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1091), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1090), .A2(new_n1115), .ZN(G390));
  NAND3_X1  g0916(.A1(new_n930), .A2(new_n771), .A3(new_n937), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n767), .B1(new_n249), .B2(new_n852), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  INV_X1    g0919(.A(G128), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n287), .B1(new_n793), .B2(new_n1119), .C1(new_n818), .C2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(G159), .B2(new_n1056), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n815), .A2(G137), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n808), .A2(new_n866), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(KEYINPUT54), .B(G143), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n806), .A2(new_n870), .B1(new_n809), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n800), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1004), .B2(new_n1128), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n281), .B1(new_n808), .B2(new_n557), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1106), .B(new_n1131), .C1(G283), .C2(new_n798), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n809), .A2(new_n541), .B1(new_n793), .B2(new_n820), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G116), .B2(new_n826), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n869), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n816), .A2(new_n486), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1130), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1118), .B1(new_n1137), .B2(new_n783), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1117), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n927), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n930), .B(new_n937), .C1(new_n895), .C2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n706), .B(new_n839), .C1(new_n755), .C2(new_n758), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n891), .B1(new_n1142), .B2(new_n840), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n923), .A2(new_n965), .A3(new_n936), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n965), .B1(new_n923), .B2(new_n936), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n927), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1141), .A2(new_n1146), .ZN(new_n1147));
  AND4_X1   g0947(.A1(G330), .A2(new_n971), .A3(new_n841), .A4(new_n891), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1148), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1141), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1139), .B1(new_n1152), .B2(new_n1014), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n893), .A2(new_n894), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n891), .B1(new_n748), .B2(new_n841), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n1148), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT116), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT116), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1158), .B(new_n1154), .C1(new_n1155), .C2(new_n1148), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1155), .A2(new_n1148), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1142), .A2(new_n840), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n453), .A2(new_n748), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n941), .A2(new_n942), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n727), .B1(new_n1152), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1149), .A2(new_n1151), .A3(new_n1166), .A4(new_n1163), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1153), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n321), .A2(new_n322), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n276), .A2(new_n704), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT55), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1175), .A2(new_n309), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1177), .B1(new_n1175), .B2(new_n309), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1174), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1180), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n1173), .A3(new_n1178), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n970), .B2(G330), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n969), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n924), .A2(new_n958), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n968), .ZN(new_n1188));
  AND4_X1   g0988(.A1(G330), .A2(new_n1184), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n940), .B1(new_n1185), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1186), .A2(new_n1188), .A3(G330), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(new_n1183), .A3(new_n1181), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n970), .A2(G330), .A3(new_n1184), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n925), .A2(new_n938), .A3(new_n939), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1190), .A2(new_n1195), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1141), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1150), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1165), .B1(new_n1199), .B2(new_n1163), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1172), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1169), .A2(new_n1166), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1202), .A2(KEYINPUT57), .A3(new_n1195), .A4(new_n1190), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n723), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1184), .A2(new_n771), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n281), .A2(new_n462), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1206), .B(new_n998), .C1(G77), .C2(new_n860), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n815), .A2(G97), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n806), .A2(new_n486), .B1(new_n809), .B2(new_n398), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n800), .A2(new_n242), .B1(new_n793), .B2(new_n990), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n798), .A2(G116), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1207), .A2(new_n1208), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT58), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1206), .B(new_n240), .C1(G33), .C2(G41), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n818), .A2(new_n1119), .B1(new_n866), .B2(new_n788), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT117), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n808), .A2(new_n1126), .B1(new_n806), .B2(new_n1120), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G137), .B2(new_n863), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n870), .C2(new_n816), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT118), .Z(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n794), .C2(G124), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n800), .B2(new_n790), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n1224), .B2(KEYINPUT59), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1215), .B(new_n1218), .C1(new_n1225), .C2(new_n1228), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1229), .A2(new_n1012), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n768), .B(new_n1230), .C1(new_n201), .C2(new_n851), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1205), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1196), .B2(new_n1014), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1204), .A2(new_n1234), .ZN(G375));
  NAND2_X1  g1035(.A1(new_n1163), .A2(new_n1015), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n768), .B1(new_n220), .B2(new_n851), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n798), .A2(G132), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT122), .Z(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n865), .B2(new_n806), .C1(new_n816), .C2(new_n1126), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT123), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n808), .A2(new_n333), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n809), .A2(new_n866), .B1(new_n793), .B2(new_n1120), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n287), .B1(new_n788), .B2(new_n240), .C1(new_n800), .C2(new_n242), .ZN(new_n1245));
  NOR4_X1   g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n818), .A2(new_n820), .B1(new_n809), .B2(new_n486), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n815), .B2(G116), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT121), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n788), .A2(new_n398), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G283), .A2(new_n826), .B1(new_n794), .B2(G303), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n281), .C1(new_n476), .C2(new_n808), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1251), .B(new_n1253), .C1(G77), .C2(new_n801), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1246), .A2(new_n1247), .B1(new_n1250), .B2(new_n1254), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1237), .B1(new_n1255), .B2(new_n1012), .C1(new_n891), .C2(new_n772), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1236), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1156), .A2(KEYINPUT116), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n1165), .A3(new_n1159), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1033), .B(KEYINPUT120), .Z(new_n1261));
  NAND3_X1  g1061(.A1(new_n1167), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1262), .ZN(G381));
  OR4_X1    g1063(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1204), .A2(new_n1170), .A3(new_n1234), .ZN(new_n1265));
  OR4_X1    g1065(.A1(G387), .A2(new_n1264), .A3(new_n1265), .A4(G381), .ZN(G407));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n705), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(new_n1265), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT127), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(G2897), .ZN(new_n1272));
  AND4_X1   g1072(.A1(new_n1165), .A2(new_n1157), .A3(new_n1159), .A4(new_n1162), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(KEYINPUT60), .B2(new_n1167), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n723), .B1(new_n1260), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(KEYINPUT124), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1165), .B1(new_n1259), .B2(new_n1159), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1260), .B1(new_n1278), .B2(new_n1275), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n727), .B1(new_n1273), .B2(KEYINPUT60), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT124), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1277), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1283), .B2(new_n1258), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n876), .B(new_n1257), .C1(new_n1277), .C2(new_n1282), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1272), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1274), .A2(new_n1276), .A3(KEYINPUT124), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1281), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1258), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n876), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1283), .A2(G384), .A3(new_n1258), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1272), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1290), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1204), .A2(G378), .A3(new_n1234), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1261), .ZN(new_n1295));
  NOR3_X1   g1095(.A1(new_n1196), .A2(new_n1200), .A3(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1170), .B1(new_n1296), .B2(new_n1233), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1286), .A2(new_n1293), .B1(new_n1298), .B2(new_n1269), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1271), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1303));
  AND4_X1   g1103(.A1(new_n1302), .A2(new_n1298), .A3(new_n1269), .A4(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1268), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1302), .B1(new_n1305), .B2(new_n1303), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1286), .A2(new_n1293), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1298), .A2(new_n1269), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1300), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(KEYINPUT127), .A3(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1301), .A2(new_n1307), .A3(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G390), .B(new_n1013), .C1(new_n1034), .C2(new_n1054), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(G393), .B(new_n835), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(G387), .A2(new_n1090), .A3(new_n1115), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1314), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1319), .A2(KEYINPUT125), .A3(new_n1314), .A4(new_n1317), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1313), .A2(new_n1323), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1299), .A2(new_n1323), .A3(KEYINPUT61), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1305), .A2(KEYINPUT63), .A3(new_n1303), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1303), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1327), .B1(new_n1309), .B2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1325), .A2(new_n1326), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1324), .A2(new_n1330), .ZN(G405));
  NAND2_X1  g1131(.A1(G375), .A2(new_n1170), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1323), .A2(new_n1294), .A3(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1294), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1321), .A2(new_n1334), .A3(new_n1322), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(new_n1336), .B(new_n1328), .ZN(G402));
endmodule


