//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT64), .B(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n231), .B(new_n234), .Z(G358));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G58), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G351));
  NAND2_X1  g0044(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT8), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G58), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(new_n212), .A3(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n251), .A2(new_n254), .B1(new_n252), .B2(new_n248), .ZN(new_n255));
  AND2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(KEYINPUT7), .B1(new_n258), .B2(new_n213), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  NOR4_X1   g0060(.A1(new_n256), .A2(new_n257), .A3(new_n260), .A4(G20), .ZN(new_n261));
  OAI21_X1  g0061(.A(G68), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G68), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n202), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G58), .A2(G68), .ZN(new_n265));
  OAI21_X1  g0065(.A(G20), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G159), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n262), .A2(KEYINPUT16), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  OR2_X1    g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(new_n213), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n260), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n269), .B1(new_n278), .B2(G68), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT16), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n253), .A2(new_n212), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n262), .A2(new_n270), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT16), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n255), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI211_X1 g0089(.A(G226), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(KEYINPUT71), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT71), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n292), .A2(new_n293), .A3(G226), .A4(G1698), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G87), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n292), .A2(G223), .A3(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n291), .A2(new_n294), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G41), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  AOI21_X1  g0102(.A(G1), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n305), .A3(G274), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n228), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(G169), .B1(new_n300), .B2(new_n310), .ZN(new_n311));
  AOI211_X1 g0111(.A(G179), .B(new_n309), .C1(new_n298), .C2(new_n299), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT72), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G179), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n300), .A2(new_n314), .A3(new_n310), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT72), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n309), .B1(new_n298), .B2(new_n299), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n315), .B(new_n316), .C1(G169), .C2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT73), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n313), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n319), .B1(new_n313), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n289), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT18), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g0124(.A(KEYINPUT18), .B(new_n289), .C1(new_n320), .C2(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n252), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n263), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT12), .ZN(new_n329));
  INV_X1    g0129(.A(G33), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(G20), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(G77), .B1(G20), .B2(new_n263), .ZN(new_n332));
  INV_X1    g0132(.A(new_n267), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n201), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n335));
  INV_X1    g0135(.A(new_n254), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(G68), .A3(new_n250), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n329), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT11), .B1(new_n334), .B2(new_n283), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT68), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n306), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G274), .ZN(new_n345));
  INV_X1    g0145(.A(new_n212), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n346), .B2(new_n304), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(KEYINPUT68), .A3(new_n303), .ZN(new_n348));
  INV_X1    g0148(.A(new_n308), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n344), .A2(new_n348), .B1(G238), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n292), .A2(G232), .A3(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  OAI211_X1 g0152(.A(G226), .B(new_n296), .C1(new_n256), .C2(new_n257), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n299), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT13), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n350), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n350), .B2(new_n355), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n342), .B(G169), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n358), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n350), .A2(new_n355), .A3(new_n356), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n359), .B1(new_n362), .B2(new_n314), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n342), .B1(new_n362), .B2(G169), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n341), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  INV_X1    g0166(.A(new_n331), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n366), .A2(new_n367), .B1(new_n213), .B2(new_n217), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT8), .B(G58), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n333), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n283), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT67), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n217), .B1(new_n249), .B2(G20), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n336), .A2(new_n373), .B1(new_n217), .B2(new_n327), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n292), .A2(G238), .A3(G1698), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n292), .A2(G232), .A3(new_n296), .ZN(new_n377));
  INV_X1    g0177(.A(G107), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n376), .B(new_n377), .C1(new_n378), .C2(new_n292), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n299), .ZN(new_n380));
  INV_X1    g0180(.A(new_n216), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n349), .A2(new_n381), .B1(new_n347), .B2(new_n303), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G169), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n375), .B(new_n385), .C1(G179), .C2(new_n383), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n383), .A2(G200), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n380), .A2(G190), .A3(new_n382), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n372), .A3(new_n388), .A4(new_n374), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n357), .A2(new_n358), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n341), .B1(new_n391), .B2(G190), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT69), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n362), .B2(G200), .ZN(new_n394));
  INV_X1    g0194(.A(G200), .ZN(new_n395));
  AOI211_X1 g0195(.A(KEYINPUT69), .B(new_n395), .C1(new_n360), .C2(new_n361), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n392), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n248), .A2(new_n331), .B1(G150), .B2(new_n267), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n284), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n250), .A2(G50), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n254), .A2(new_n401), .B1(G50), .B2(new_n252), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G226), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n306), .B1(new_n405), .B2(new_n308), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n292), .A2(G222), .A3(new_n296), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n292), .A2(G223), .A3(G1698), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(new_n217), .C2(new_n292), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n409), .B2(new_n299), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n404), .B1(new_n410), .B2(G169), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n410), .A2(new_n314), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n403), .A2(KEYINPUT9), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT9), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n400), .B2(new_n402), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT10), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n410), .A2(new_n395), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(G190), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n417), .A2(new_n418), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n421), .A2(new_n414), .A3(new_n416), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT10), .B1(new_n423), .B2(new_n419), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n413), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AND4_X1   g0225(.A1(new_n365), .A2(new_n390), .A3(new_n397), .A4(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n280), .B1(new_n279), .B2(KEYINPUT16), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n263), .B1(new_n276), .B2(new_n277), .ZN(new_n428));
  NOR4_X1   g0228(.A1(new_n428), .A2(KEYINPUT70), .A3(new_n269), .A4(new_n286), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n287), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G190), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n300), .A2(new_n431), .A3(new_n310), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(G200), .B2(new_n317), .ZN(new_n433));
  INV_X1    g0233(.A(new_n255), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT17), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n288), .A2(KEYINPUT17), .A3(new_n433), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT74), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT74), .B1(new_n437), .B2(new_n438), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n326), .A2(new_n426), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT75), .B1(new_n330), .B2(G1), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT75), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n445), .A2(new_n249), .A3(G33), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G97), .B1(new_n447), .B2(new_n254), .ZN(new_n448));
  INV_X1    g0248(.A(G97), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n252), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(KEYINPUT76), .A3(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G107), .B1(new_n259), .B2(new_n261), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT6), .ZN(new_n457));
  AND2_X1   g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  NOR2_X1   g0258(.A1(G97), .A2(G107), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n378), .A2(KEYINPUT6), .A3(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n462), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(new_n283), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n455), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  OAI211_X1 g0267(.A(G250), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n468));
  OAI211_X1 g0268(.A(G244), .B(new_n296), .C1(new_n256), .C2(new_n257), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT77), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(KEYINPUT4), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n469), .A2(new_n471), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n299), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n249), .A2(G45), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n299), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n477), .A2(new_n476), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n478), .A2(G257), .B1(new_n479), .B2(new_n347), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n384), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n474), .A2(new_n314), .A3(new_n480), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n466), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n453), .A2(new_n454), .B1(new_n464), .B2(new_n283), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(G200), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n474), .A2(G190), .A3(new_n480), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n252), .A2(G116), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n447), .A2(new_n254), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(G116), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n467), .B(new_n213), .C1(G33), .C2(new_n449), .ZN(new_n493));
  INV_X1    g0293(.A(G116), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G20), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n283), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT20), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n493), .A2(new_n283), .A3(KEYINPUT20), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n492), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G264), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n503));
  OAI211_X1 g0303(.A(G257), .B(new_n296), .C1(new_n256), .C2(new_n257), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n273), .A2(G303), .A3(new_n274), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n299), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n478), .A2(G270), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n479), .A2(new_n347), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n502), .A2(new_n314), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(KEYINPUT80), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n299), .A2(new_n506), .B1(new_n478), .B2(G270), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT80), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n509), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n384), .B1(new_n492), .B2(new_n500), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT21), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n512), .A2(new_n515), .A3(new_n519), .A4(new_n516), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n511), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n512), .A2(new_n515), .A3(G200), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n512), .A2(new_n515), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n502), .B(new_n522), .C1(new_n523), .C2(new_n431), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n475), .A2(G250), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT78), .B1(new_n299), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT78), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n305), .A2(new_n527), .A3(G250), .A4(new_n475), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n526), .A2(new_n528), .B1(new_n476), .B2(new_n347), .ZN(new_n529));
  OAI211_X1 g0329(.A(G238), .B(new_n296), .C1(new_n256), .C2(new_n257), .ZN(new_n530));
  OAI211_X1 g0330(.A(G244), .B(G1698), .C1(new_n256), .C2(new_n257), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G116), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n299), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G200), .ZN(new_n536));
  INV_X1    g0336(.A(new_n366), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n252), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n292), .A2(new_n213), .A3(G68), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n367), .B2(new_n449), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n449), .A3(new_n378), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT79), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT79), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(new_n542), .A3(new_n449), .A4(new_n378), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n352), .A2(new_n540), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(G20), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n539), .B(new_n541), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n538), .B1(new_n550), .B2(new_n283), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n529), .A2(new_n534), .A3(G190), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n491), .A2(G87), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n536), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n549), .B1(new_n544), .B2(new_n546), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n541), .A2(new_n539), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n283), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n538), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n491), .A2(new_n537), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n529), .A2(new_n534), .A3(G179), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n384), .B1(new_n529), .B2(new_n534), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n554), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n489), .A2(new_n521), .A3(new_n524), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT81), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT25), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n252), .B2(G107), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n327), .A2(KEYINPUT25), .A3(new_n378), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n491), .A2(G107), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n213), .B(G87), .C1(new_n256), .C2(new_n257), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT22), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT22), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n292), .A2(new_n574), .A3(new_n213), .A4(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n532), .A2(G20), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT23), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n213), .B2(G107), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n378), .A2(KEYINPUT23), .A3(G20), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n577), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT24), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT24), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(new_n584), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n571), .B1(new_n586), .B2(new_n283), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n478), .A2(G264), .B1(new_n479), .B2(new_n347), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n589));
  OAI211_X1 g0389(.A(G250), .B(new_n296), .C1(new_n256), .C2(new_n257), .ZN(new_n590));
  NAND2_X1  g0390(.A1(G33), .A2(G294), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n299), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n384), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G179), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n566), .B1(new_n587), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(G169), .B1(new_n588), .B2(new_n593), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n588), .A2(new_n593), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n598), .B1(new_n314), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n585), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n584), .B1(new_n576), .B2(new_n581), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n283), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n600), .B(KEYINPUT81), .C1(new_n604), .C2(new_n571), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n594), .A2(G200), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n588), .A2(new_n593), .A3(G190), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n603), .A2(new_n570), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n597), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT82), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n597), .A2(new_n605), .A3(KEYINPUT82), .A4(new_n608), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n565), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n443), .A2(new_n613), .ZN(G372));
  INV_X1    g0414(.A(new_n484), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n564), .A2(KEYINPUT26), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n560), .ZN(new_n617));
  OAI21_X1  g0417(.A(KEYINPUT83), .B1(new_n561), .B2(new_n562), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n535), .A2(G169), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n529), .A2(new_n534), .A3(G179), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n617), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n554), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n623), .A2(new_n624), .A3(new_n484), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n616), .B1(new_n625), .B2(KEYINPUT26), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n618), .A2(new_n622), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n560), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n518), .A2(new_n520), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n600), .B1(new_n604), .B2(new_n571), .ZN(new_n630));
  INV_X1    g0430(.A(new_n511), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n608), .A2(new_n484), .A3(new_n488), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n623), .A2(new_n624), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n626), .A2(new_n628), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n443), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n340), .B1(new_n362), .B2(new_n431), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n362), .A2(new_n393), .A3(G200), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT69), .B1(new_n391), .B2(new_n395), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n365), .B1(new_n642), .B2(new_n386), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT74), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT17), .B1(new_n288), .B2(new_n433), .ZN(new_n645));
  AND4_X1   g0445(.A1(KEYINPUT17), .A2(new_n430), .A3(new_n433), .A4(new_n434), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT74), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n643), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n283), .B1(new_n279), .B2(KEYINPUT16), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n281), .B2(new_n272), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n313), .B(new_n318), .C1(new_n651), .C2(new_n255), .ZN(new_n652));
  XNOR2_X1  g0452(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n652), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n422), .A2(new_n424), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n413), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n638), .A2(new_n658), .ZN(G369));
  INV_X1    g0459(.A(G330), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n521), .A2(new_n524), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT86), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n249), .A2(new_n213), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(G213), .ZN(new_n666));
  XOR2_X1   g0466(.A(new_n666), .B(KEYINPUT85), .Z(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n502), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n662), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n629), .A2(new_n631), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n672), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(KEYINPUT87), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT87), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n674), .A2(new_n679), .A3(new_n676), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n660), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n611), .A2(new_n612), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n670), .B1(new_n604), .B2(new_n571), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n630), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n670), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n675), .A2(new_n671), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT88), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n671), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n688), .A2(new_n691), .A3(new_n692), .ZN(G399));
  NAND2_X1  g0493(.A1(new_n547), .A2(new_n494), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n207), .A2(new_n301), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G1), .ZN(new_n696));
  OAI22_X1  g0496(.A1(new_n694), .A2(new_n696), .B1(new_n210), .B2(new_n695), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n455), .A2(new_n465), .B1(new_n481), .B2(new_n384), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n554), .A3(new_n563), .A4(new_n483), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n628), .B1(new_n701), .B2(KEYINPUT26), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n628), .A2(new_n615), .A3(new_n554), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(KEYINPUT26), .B2(new_n703), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n633), .A2(new_n624), .A3(new_n623), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n521), .A2(new_n597), .A3(new_n605), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI211_X1 g0507(.A(new_n699), .B(new_n670), .C1(new_n704), .C2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT29), .B1(new_n637), .B2(new_n671), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g0510(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n599), .A2(new_n561), .A3(new_n513), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n481), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n513), .A2(new_n593), .A3(new_n588), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n621), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n474), .A2(new_n480), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n512), .A2(new_n515), .A3(new_n314), .A4(new_n535), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT90), .B1(new_n718), .B2(new_n599), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT90), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n481), .A2(new_n723), .A3(new_n594), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n721), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n670), .B(new_n712), .C1(new_n720), .C2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT30), .B1(new_n717), .B2(new_n718), .ZN(new_n727));
  NOR4_X1   g0527(.A1(new_n716), .A2(new_n481), .A3(new_n621), .A4(new_n713), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n722), .A2(new_n724), .ZN(new_n730));
  INV_X1    g0530(.A(new_n721), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n671), .B1(new_n729), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n726), .B1(new_n733), .B2(KEYINPUT31), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n734), .B1(new_n613), .B2(new_n671), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n660), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n710), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n698), .B1(new_n737), .B2(G1), .ZN(G364));
  AND2_X1   g0538(.A1(new_n213), .A2(G13), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n249), .B1(new_n739), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n695), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n681), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n678), .A2(new_n660), .A3(new_n680), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n212), .B1(G20), .B2(new_n384), .ZN(new_n747));
  NAND2_X1  g0547(.A1(G20), .A2(G179), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT92), .Z(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n395), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G326), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n213), .B1(new_n754), .B2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n749), .A2(new_n431), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n752), .B1(new_n753), .B2(new_n755), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT94), .Z(new_n761));
  NOR4_X1   g0561(.A1(new_n213), .A2(new_n431), .A3(new_n395), .A4(G179), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n292), .B1(new_n762), .B2(G303), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT95), .Z(new_n764));
  NOR4_X1   g0564(.A1(new_n213), .A2(new_n395), .A3(G179), .A4(G190), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  INV_X1    g0567(.A(G329), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n754), .A2(G20), .A3(new_n431), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n750), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n771), .B2(G322), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n756), .A2(new_n395), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(G317), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n772), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n761), .A2(new_n764), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n751), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n201), .A2(new_n779), .B1(new_n774), .B2(new_n263), .ZN(new_n780));
  INV_X1    g0580(.A(new_n771), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n202), .A2(new_n781), .B1(new_n758), .B2(new_n217), .ZN(new_n782));
  INV_X1    g0582(.A(new_n769), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G159), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  INV_X1    g0585(.A(new_n755), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G97), .B1(new_n765), .B2(G107), .ZN(new_n787));
  INV_X1    g0587(.A(new_n762), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n787), .B(new_n292), .C1(new_n542), .C2(new_n788), .ZN(new_n789));
  NOR4_X1   g0589(.A1(new_n780), .A2(new_n782), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n747), .B1(new_n778), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n292), .A2(new_n207), .ZN(new_n793));
  INV_X1    g0593(.A(G355), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n793), .A2(new_n794), .B1(G116), .B2(new_n207), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n238), .A2(G45), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n258), .A2(new_n207), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n302), .B2(new_n211), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n795), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n747), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n743), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT91), .ZN(new_n806));
  INV_X1    g0606(.A(new_n802), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n792), .B(new_n806), .C1(new_n677), .C2(new_n807), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n746), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G396));
  INV_X1    g0610(.A(new_n743), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n747), .A2(new_n800), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(new_n217), .B2(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G116), .A2(new_n757), .B1(new_n751), .B2(G303), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n753), .B2(new_n781), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n774), .A2(new_n767), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n258), .B1(new_n769), .B2(new_n759), .C1(new_n449), .C2(new_n755), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n788), .A2(new_n378), .B1(new_n766), .B2(new_n542), .ZN(new_n818));
  NOR4_X1   g0618(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n771), .B1(new_n757), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n779), .C1(new_n822), .C2(new_n774), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n292), .B1(new_n769), .B2(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n788), .A2(new_n201), .B1(new_n766), .B2(new_n263), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G58), .C2(new_n786), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n819), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n747), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n670), .A2(new_n375), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n389), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n386), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n386), .A2(new_n670), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n813), .B1(new_n829), .B2(new_n830), .C1(new_n801), .C2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n623), .B1(new_n705), .B2(new_n632), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n670), .B1(new_n838), .B2(new_n626), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(new_n835), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n736), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n736), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n811), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n841), .B1(new_n843), .B2(KEYINPUT97), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n843), .A2(KEYINPUT97), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n837), .B1(new_n845), .B2(new_n846), .ZN(G384));
  INV_X1    g0647(.A(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n667), .B1(new_n651), .B2(new_n255), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n645), .A2(new_n646), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n655), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n652), .A2(new_n435), .A3(new_n849), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(KEYINPUT99), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n849), .A2(new_n435), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n322), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT99), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n852), .A2(new_n858), .A3(KEYINPUT37), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n854), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT100), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n854), .A2(new_n857), .A3(KEYINPUT100), .A4(new_n859), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n287), .A2(KEYINPUT98), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n865), .A2(new_n282), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n287), .A2(KEYINPUT98), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n255), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n313), .A2(new_n318), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n435), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(new_n668), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT37), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n857), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n647), .A2(new_n648), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n324), .B2(new_n325), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n867), .A2(new_n282), .A3(new_n865), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n434), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n667), .ZN(new_n878));
  OAI211_X1 g0678(.A(KEYINPUT38), .B(new_n873), .C1(new_n875), .C2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n848), .B1(new_n864), .B2(new_n880), .ZN(new_n881));
  OR2_X1    g0681(.A1(new_n365), .A2(new_n670), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n878), .B1(new_n326), .B2(new_n441), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n877), .A2(new_n313), .A3(new_n318), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(new_n435), .A3(new_n878), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .B1(new_n322), .B2(new_n856), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n879), .A3(KEYINPUT39), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n881), .A2(new_n883), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n879), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n365), .A2(new_n397), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n670), .A2(new_n341), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n893), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n637), .A2(new_n671), .A3(new_n836), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n896), .B2(new_n834), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n652), .B(new_n653), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n892), .A2(new_n897), .B1(new_n898), .B2(new_n668), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n898), .B1(new_n441), .B2(new_n643), .ZN(new_n901));
  INV_X1    g0701(.A(new_n657), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n412), .B2(new_n411), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n710), .B2(new_n443), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT101), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n900), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n613), .A2(new_n671), .ZN(new_n907));
  OAI211_X1 g0707(.A(KEYINPUT31), .B(new_n670), .C1(new_n720), .C2(new_n725), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n733), .B2(new_n712), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n894), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n893), .B(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n911), .A2(KEYINPUT40), .A3(new_n836), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n860), .A2(new_n861), .ZN(new_n915));
  INV_X1    g0715(.A(new_n851), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(new_n863), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n884), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n914), .B1(new_n918), .B2(new_n879), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n913), .A2(new_n836), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n909), .B1(new_n613), .B2(new_n671), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT40), .B1(new_n892), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n921), .A2(new_n442), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(G330), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n906), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n929), .A2(KEYINPUT102), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(KEYINPUT102), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n906), .A2(new_n928), .B1(new_n249), .B2(new_n739), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n462), .A2(KEYINPUT35), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n934), .A2(G116), .A3(new_n214), .A4(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT36), .Z(new_n937));
  OAI211_X1 g0737(.A(new_n211), .B(G77), .C1(new_n202), .C2(new_n263), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n201), .A2(G68), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n249), .B(G13), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n933), .A2(new_n937), .A3(new_n940), .ZN(G367));
  INV_X1    g0741(.A(new_n691), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n489), .B1(new_n485), .B2(new_n671), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n615), .A2(new_n670), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n943), .B1(new_n597), .B2(new_n605), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n671), .B1(new_n948), .B2(new_n615), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT43), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n551), .A2(new_n553), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n670), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n628), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n635), .B2(new_n954), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n950), .A2(new_n951), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n952), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n681), .A2(new_n687), .A3(new_n945), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n695), .B(KEYINPUT41), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT103), .B1(new_n687), .B2(new_n690), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n681), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n681), .A2(new_n964), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n966), .A2(new_n967), .A3(new_n691), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n681), .A2(new_n964), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n942), .B1(new_n969), .B2(new_n965), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n737), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n691), .A2(new_n692), .A3(new_n945), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT45), .Z(new_n975));
  AOI21_X1  g0775(.A(new_n945), .B1(new_n691), .B2(new_n692), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT44), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n975), .A2(new_n688), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n688), .B1(new_n975), .B2(new_n977), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n691), .B1(new_n966), .B2(new_n967), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n969), .A2(new_n942), .A3(new_n965), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(KEYINPUT104), .A3(new_n737), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n973), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n962), .B1(new_n985), .B2(new_n737), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n961), .B1(new_n986), .B2(new_n741), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n292), .B1(new_n769), .B2(new_n821), .C1(new_n263), .C2(new_n755), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n788), .A2(new_n202), .B1(new_n766), .B2(new_n217), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n988), .B(new_n989), .C1(new_n757), .C2(G50), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G143), .A2(new_n751), .B1(new_n771), .B2(G150), .ZN(new_n991));
  INV_X1    g0791(.A(G159), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n990), .B(new_n991), .C1(new_n992), .C2(new_n774), .ZN(new_n993));
  INV_X1    g0793(.A(G303), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n994), .A2(new_n781), .B1(new_n779), .B2(new_n759), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT105), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(KEYINPUT106), .B(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n258), .B1(new_n998), .B2(new_n769), .C1(new_n378), .C2(new_n755), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G97), .B2(new_n765), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n762), .A2(G116), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT46), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G283), .A2(new_n757), .B1(new_n773), .B2(G294), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n997), .A2(new_n1000), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n995), .A2(new_n996), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n993), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n747), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n956), .A2(new_n802), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n803), .B1(new_n207), .B2(new_n366), .C1(new_n234), .C2(new_n797), .ZN(new_n1010));
  NAND4_X1  g0810(.A1(new_n1008), .A2(new_n743), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n987), .A2(new_n1011), .ZN(G387));
  NAND2_X1  g0812(.A1(new_n973), .A2(new_n984), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n742), .C1(new_n737), .C2(new_n983), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n684), .A2(new_n686), .A3(new_n802), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n694), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1016), .A2(new_n793), .B1(G107), .B2(new_n207), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n694), .C1(G68), .C2(G77), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n1018), .A2(KEYINPUT107), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(KEYINPUT107), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n369), .A2(G50), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n797), .B1(new_n231), .B2(G45), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1017), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n743), .B1(new_n1025), .B2(new_n804), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G50), .A2(new_n771), .B1(new_n757), .B2(G68), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n773), .A2(new_n248), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n292), .B1(new_n822), .B2(new_n769), .C1(new_n766), .C2(new_n449), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n755), .A2(new_n366), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n788), .A2(new_n217), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n751), .A2(G159), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1027), .A2(new_n1028), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G303), .A2(new_n757), .B1(new_n751), .B2(G322), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n759), .B2(new_n774), .C1(new_n781), .C2(new_n998), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n788), .A2(new_n753), .B1(new_n767), .B2(new_n755), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n292), .B1(new_n783), .B2(G326), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(new_n494), .C2(new_n766), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT49), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1034), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1026), .B1(new_n1045), .B2(new_n747), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n983), .A2(new_n741), .B1(new_n1015), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1014), .A2(new_n1047), .ZN(G393));
  AND2_X1   g0848(.A1(new_n985), .A2(new_n742), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n980), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT110), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n984), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT104), .B1(new_n983), .B2(new_n737), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1050), .B(new_n1051), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1013), .B2(new_n1050), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1049), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n943), .A2(new_n802), .A3(new_n944), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n243), .A2(new_n797), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n803), .B1(new_n449), .B2(new_n207), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n743), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT108), .Z(new_n1062));
  AOI22_X1  g0862(.A1(G311), .A2(new_n771), .B1(new_n751), .B2(G317), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1063), .B(new_n1064), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n788), .A2(new_n767), .B1(new_n494), .B2(new_n755), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n292), .B1(new_n783), .B2(G322), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n378), .B2(new_n766), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1066), .B(new_n1068), .C1(new_n757), .C2(G294), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n994), .B2(new_n774), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G150), .A2(new_n751), .B1(new_n771), .B2(G159), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n788), .A2(new_n263), .B1(new_n217), .B2(new_n755), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n258), .B1(new_n783), .B2(G143), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n542), .B2(new_n766), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1073), .B(new_n1075), .C1(new_n773), .C2(G50), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n369), .B2(new_n758), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1065), .A2(new_n1070), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1062), .B1(new_n1078), .B2(new_n747), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n980), .A2(new_n741), .B1(new_n1058), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1057), .A2(new_n1080), .ZN(G390));
  NOR2_X1   g0881(.A1(new_n835), .A2(new_n660), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n921), .A2(new_n895), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT111), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n897), .B2(new_n883), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n834), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n839), .B2(new_n836), .ZN(new_n1088));
  OAI211_X1 g0888(.A(KEYINPUT111), .B(new_n882), .C1(new_n1088), .C2(new_n895), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(new_n881), .B2(new_n890), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n864), .A2(new_n880), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n707), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT26), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n564), .A2(new_n1094), .A3(new_n615), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n628), .C1(new_n625), .C2(new_n1094), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n671), .B(new_n833), .C1(new_n1093), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n834), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n882), .B1(new_n1099), .B2(new_n895), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1092), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1084), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1092), .A2(new_n1100), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n734), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n907), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1105), .A2(new_n913), .A3(new_n1082), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n890), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n918), .A2(new_n879), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1107), .B1(new_n1108), .B2(new_n848), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1103), .B(new_n1106), .C1(new_n1109), .C2(new_n1090), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1102), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n735), .A2(new_n1083), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1098), .B1(new_n1112), .B2(new_n913), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n895), .B1(new_n921), .B2(new_n1083), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n895), .B1(new_n735), .B2(new_n1083), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n670), .B(new_n565), .C1(new_n611), .C2(new_n612), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n913), .B(new_n1082), .C1(new_n1116), .C2(new_n909), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1088), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1113), .A2(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT112), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n925), .B2(G330), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n921), .A2(new_n442), .A3(KEYINPUT112), .A4(new_n660), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n904), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(KEYINPUT113), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(KEYINPUT29), .B(new_n671), .C1(new_n1093), .C2(new_n1096), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n839), .B2(KEYINPUT29), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n658), .B1(new_n1127), .B2(new_n442), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n925), .A2(G330), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(KEYINPUT112), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n925), .A2(new_n1121), .A3(G330), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1128), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1099), .A2(new_n1106), .A3(new_n1114), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT113), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1132), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1125), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1111), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1102), .A2(new_n1138), .A3(new_n1110), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n742), .A3(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1102), .A2(new_n1110), .A3(new_n741), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n811), .B1(new_n369), .B2(new_n812), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n449), .A2(new_n758), .B1(new_n774), .B2(new_n378), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G116), .B2(new_n771), .ZN(new_n1146));
  OAI221_X1 g0946(.A(new_n258), .B1(new_n217), .B2(new_n755), .C1(new_n788), .C2(new_n542), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n751), .B2(G283), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n766), .A2(new_n263), .B1(new_n753), .B2(new_n769), .ZN(new_n1149));
  XOR2_X1   g0949(.A(new_n1149), .B(KEYINPUT116), .Z(new_n1150));
  NAND3_X1  g0950(.A1(new_n1146), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n773), .A2(G137), .B1(G159), .B2(new_n786), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(KEYINPUT54), .B(G143), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n758), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT114), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n258), .B1(new_n783), .B2(G125), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n201), .B2(new_n766), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT115), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n771), .A2(G132), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n751), .A2(G128), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n762), .A2(G150), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT53), .Z(new_n1162));
  NAND4_X1  g0962(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1151), .B1(new_n1155), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT117), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n747), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1144), .B1(new_n1166), .B2(new_n1168), .C1(new_n1109), .C2(new_n801), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1143), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1142), .A2(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(new_n1153), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n771), .A2(G128), .B1(new_n762), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT118), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n773), .A2(G132), .B1(G150), .B2(new_n786), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G125), .A2(new_n751), .B1(new_n757), .B2(G137), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT59), .Z(new_n1178));
  AOI211_X1 g0978(.A(G33), .B(G41), .C1(new_n783), .C2(G124), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(new_n992), .C2(new_n766), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n378), .A2(new_n781), .B1(new_n758), .B2(new_n366), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n766), .A2(new_n202), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n755), .A2(new_n263), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n258), .B(new_n301), .C1(new_n769), .C2(new_n767), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1031), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n449), .B2(new_n774), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1181), .B(new_n1186), .C1(G116), .C2(new_n751), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1188));
  AOI21_X1  g0988(.A(G50), .B1(new_n330), .B2(new_n301), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n292), .B2(G41), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1187), .A2(KEYINPUT58), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1180), .A2(new_n1188), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1192), .A2(new_n747), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n811), .B(new_n1193), .C1(new_n201), .C2(new_n812), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n667), .A2(new_n404), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n425), .B(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n800), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1194), .A2(new_n1199), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n891), .A2(new_n899), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT40), .ZN(new_n1202));
  NOR3_X1   g1002(.A1(new_n920), .A2(new_n921), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1203), .B1(new_n864), .B2(new_n880), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n911), .A2(new_n836), .A3(new_n913), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(new_n879), .B2(new_n889), .ZN(new_n1206));
  OAI211_X1 g1006(.A(new_n1204), .B(G330), .C1(KEYINPUT40), .C2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1198), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n923), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1198), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1209), .A2(G330), .A3(new_n1204), .A4(new_n1210), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1201), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1208), .A2(new_n1211), .B1(new_n891), .B2(new_n899), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1200), .B1(new_n1214), .B2(new_n740), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1141), .A2(new_n1132), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1210), .B1(new_n924), .B2(G330), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n919), .A2(new_n923), .A3(new_n660), .A4(new_n1198), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n900), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1201), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT57), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1223), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n695), .B1(new_n1225), .B2(new_n1216), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1215), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(G375));
  NAND2_X1  g1028(.A1(new_n895), .A2(new_n800), .ZN(new_n1229));
  XNOR2_X1  g1029(.A(new_n1229), .B(KEYINPUT119), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n788), .A2(new_n992), .B1(new_n201), .B2(new_n755), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n258), .B1(new_n783), .B2(G128), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n202), .B2(new_n766), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(new_n771), .C2(G137), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n773), .A2(new_n1172), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n751), .A2(G132), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n757), .A2(G150), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n258), .B1(new_n994), .B2(new_n769), .C1(new_n766), .C2(new_n217), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1030), .B(new_n1239), .C1(G97), .C2(new_n762), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n494), .B2(new_n774), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G107), .A2(new_n757), .B1(new_n751), .B2(G294), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n767), .B2(new_n781), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1238), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT120), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n830), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1245), .B2(new_n1244), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n811), .B1(new_n263), .B2(new_n812), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1135), .A2(new_n741), .B1(new_n1230), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n962), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1250), .B1(new_n1138), .B2(new_n1253), .ZN(G381));
  AND4_X1   g1054(.A1(new_n987), .A2(new_n1057), .A3(new_n1011), .A4(new_n1080), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1014), .A2(new_n809), .A3(new_n1047), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1256), .A2(G384), .A3(G378), .A4(G381), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n1227), .A3(new_n1257), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT121), .ZN(G407));
  INV_X1    g1059(.A(G378), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1227), .A2(new_n669), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(G407), .A2(G213), .A3(new_n1261), .ZN(G409));
  NAND2_X1  g1062(.A1(G393), .A2(G396), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1256), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n987), .A2(new_n1011), .B1(new_n1057), .B2(new_n1080), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1265), .B1(new_n1255), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(G390), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n987), .A2(new_n1057), .A3(new_n1011), .A4(new_n1080), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1268), .A2(new_n1269), .A3(new_n1264), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1267), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n740), .B1(new_n1221), .B2(KEYINPUT123), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(KEYINPUT123), .B2(new_n1221), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1274), .B(new_n1200), .C1(new_n962), .C2(new_n1222), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1260), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1215), .ZN(new_n1278));
  AND4_X1   g1078(.A1(KEYINPUT122), .A2(new_n1277), .A3(G378), .A4(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT122), .B1(new_n1227), .B2(G378), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1276), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n669), .A2(G213), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n669), .A2(G213), .A3(G2897), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT60), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1251), .B1(new_n1138), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT124), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT124), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1288), .B(new_n1251), .C1(new_n1138), .C2(new_n1285), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n742), .B1(new_n1251), .B2(new_n1285), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(KEYINPUT125), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1290), .B1(new_n1286), .B2(KEYINPUT124), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT125), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1294), .A2(new_n1295), .A3(new_n1289), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(G384), .B1(new_n1297), .B2(new_n1250), .ZN(new_n1298));
  INV_X1    g1098(.A(G384), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1250), .ZN(new_n1300));
  AOI211_X1 g1100(.A(new_n1299), .B(new_n1300), .C1(new_n1293), .C2(new_n1296), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1284), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1296), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1295), .B1(new_n1294), .B2(new_n1289), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1250), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1299), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1297), .A2(G384), .A3(new_n1250), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1284), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1302), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT62), .B1(new_n1283), .B2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1281), .A2(new_n1312), .A3(new_n1282), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1272), .B1(new_n1311), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1313), .A2(KEYINPUT126), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1281), .A2(new_n1317), .A3(new_n1312), .A4(new_n1282), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT62), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1271), .B1(new_n1315), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT63), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1316), .A2(new_n1321), .A3(new_n1318), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1314), .A2(KEYINPUT63), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1271), .A2(KEYINPUT61), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1310), .A2(KEYINPUT127), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT127), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1302), .A2(new_n1309), .A3(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1325), .A2(new_n1283), .A3(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1320), .A2(new_n1329), .ZN(G405));
  INV_X1    g1130(.A(new_n1312), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G375), .A2(new_n1260), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1271), .A2(new_n1332), .A3(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1271), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1331), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1271), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1340), .A2(new_n1312), .A3(new_n1334), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1337), .A2(new_n1341), .ZN(G402));
endmodule


