//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n494, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XNOR2_X1  g016(.A(KEYINPUT66), .B(G57), .ZN(G237));
  XNOR2_X1  g017(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT69), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT68), .B(KEYINPUT2), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(new_n453), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT70), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT72), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT71), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(KEYINPUT3), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n473), .A2(KEYINPUT71), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT73), .B1(new_n480), .B2(G137), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n475), .B1(KEYINPUT72), .B2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT3), .B1(new_n469), .B2(KEYINPUT71), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n479), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AND4_X1   g059(.A1(KEYINPUT73), .A2(new_n484), .A3(G137), .A4(new_n464), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n472), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT74), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(G137), .A3(new_n464), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n484), .A2(KEYINPUT73), .A3(G137), .A4(new_n464), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(new_n493), .A3(new_n472), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n468), .B1(new_n487), .B2(new_n494), .ZN(G160));
  OAI21_X1  g070(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G112), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n480), .A2(G136), .ZN(new_n499));
  XOR2_X1   g074(.A(new_n499), .B(KEYINPUT75), .Z(new_n500));
  AOI21_X1  g075(.A(new_n464), .B1(new_n477), .B2(new_n479), .ZN(new_n501));
  AOI211_X1 g076(.A(new_n498), .B(new_n500), .C1(G124), .C2(new_n501), .ZN(G162));
  NAND2_X1  g077(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n478), .A2(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(new_n464), .A3(G138), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT76), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT76), .ZN(new_n509));
  INV_X1    g084(.A(G138), .ZN(new_n510));
  NOR3_X1   g085(.A1(new_n510), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n465), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n510), .A2(G2105), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n477), .B2(new_n479), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n508), .B(new_n512), .C1(new_n515), .C2(new_n506), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT77), .ZN(new_n517));
  OAI21_X1  g092(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n518));
  INV_X1    g093(.A(G114), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(G2105), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n501), .B2(G126), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n517), .B1(new_n516), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(G164));
  XNOR2_X1  g099(.A(KEYINPUT78), .B(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT6), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G50), .ZN(new_n532));
  OR2_X1    g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(KEYINPUT5), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n529), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G88), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n535), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n525), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n532), .A2(new_n538), .A3(new_n540), .ZN(G303));
  INV_X1    g116(.A(G303), .ZN(G166));
  NAND2_X1  g117(.A1(new_n531), .A2(G51), .ZN(new_n543));
  XNOR2_X1  g118(.A(KEYINPUT80), .B(G89), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n537), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT79), .B(KEYINPUT7), .ZN(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AND2_X1   g123(.A1(G63), .A2(G651), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n548), .B1(new_n535), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n543), .A2(new_n545), .A3(new_n550), .ZN(G286));
  INV_X1    g126(.A(G286), .ZN(G168));
  NAND2_X1  g127(.A1(new_n537), .A2(G90), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n531), .A2(G52), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n525), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  NAND2_X1  g133(.A1(new_n537), .A2(G81), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n531), .A2(G43), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n535), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n525), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g141(.A(KEYINPUT81), .B(KEYINPUT8), .Z(new_n567));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  OR2_X1    g145(.A1(new_n527), .A2(new_n528), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G543), .ZN(new_n572));
  NAND2_X1  g147(.A1(KEYINPUT82), .A2(G53), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT9), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n531), .A2(KEYINPUT82), .A3(new_n575), .A4(G53), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n537), .A2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G65), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n536), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n577), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n529), .A2(new_n585), .A3(new_n530), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT83), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n535), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n537), .A2(G87), .B1(G651), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  INV_X1    g165(.A(new_n525), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n535), .A2(G61), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT84), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI211_X1 g170(.A(G48), .B(G543), .C1(new_n527), .C2(new_n528), .ZN(new_n596));
  OAI211_X1 g171(.A(G86), .B(new_n535), .C1(new_n527), .C2(new_n528), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n537), .A2(G85), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n531), .A2(G47), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n525), .C2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n537), .A2(G92), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT10), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n536), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n531), .A2(G54), .B1(G651), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n603), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n564), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n465), .A2(new_n470), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n480), .A2(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n464), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n501), .A2(new_n632), .A3(G123), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n632), .B1(new_n501), .B2(G123), .ZN(new_n634));
  OAI221_X1 g209(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(G2096), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n628), .A2(new_n636), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT14), .ZN(new_n644));
  XOR2_X1   g219(.A(G1341), .B(G1348), .Z(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2451), .B(G2454), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(KEYINPUT87), .B(KEYINPUT18), .Z(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  INV_X1    g237(.A(new_n655), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n658), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(KEYINPUT88), .B(KEYINPUT19), .Z(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1956), .B(G2474), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1961), .B(G1966), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n673), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT20), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n670), .A2(new_n674), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(KEYINPUT89), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(KEYINPUT89), .ZN(new_n680));
  AOI211_X1 g255(.A(new_n675), .B(new_n677), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT90), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT91), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n683), .B(new_n688), .ZN(G229));
  NAND2_X1  g264(.A1(new_n480), .A2(G131), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n501), .A2(G119), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n464), .A2(G107), .ZN(new_n692));
  OAI21_X1  g267(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT35), .B(G1991), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  MUX2_X1   g272(.A(G24), .B(G290), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT92), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n701), .A2(G22), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G166), .B2(new_n701), .ZN(new_n709));
  INV_X1    g284(.A(G1971), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n704), .A2(new_n706), .ZN(new_n712));
  NOR2_X1   g287(.A1(G6), .A2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G305), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G16), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT32), .B(G1981), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND4_X1  g292(.A1(new_n707), .A2(new_n711), .A3(new_n712), .A4(new_n717), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n697), .B(new_n700), .C1(new_n718), .C2(KEYINPUT34), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(KEYINPUT34), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(KEYINPUT36), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n720), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(G4), .A2(G16), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n612), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT94), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1348), .ZN(new_n727));
  NAND2_X1  g302(.A1(G160), .A2(G29), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G34), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n728), .B1(G29), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  NOR3_X1   g309(.A1(new_n727), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n736), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G2090), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT101), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n701), .A2(G19), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(new_n564), .B2(new_n701), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1341), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT98), .B(KEYINPUT31), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G11), .ZN(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT99), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n701), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n701), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n751), .B1(new_n736), .B2(new_n635), .C1(new_n753), .C2(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n736), .A2(G32), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n480), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n501), .A2(G129), .ZN(new_n757));
  NAND3_X1  g332(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT26), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n760), .A2(new_n761), .B1(G105), .B2(new_n470), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n756), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n755), .B1(new_n764), .B2(new_n736), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT27), .B(G1996), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n736), .A2(G26), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT28), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n480), .A2(G140), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n501), .A2(G128), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n464), .A2(G116), .ZN(new_n772));
  OAI21_X1  g347(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n769), .B1(new_n774), .B2(G29), .ZN(new_n775));
  INV_X1    g350(.A(G2067), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n744), .A2(new_n754), .A3(new_n767), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n736), .A2(G27), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT100), .Z(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n736), .ZN(new_n781));
  INV_X1    g356(.A(G2078), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n778), .B(new_n783), .C1(new_n739), .C2(G2090), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n701), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT102), .ZN(new_n788));
  INV_X1    g363(.A(G1956), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  INV_X1    g366(.A(G127), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n505), .B2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n464), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n794), .B2(new_n793), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT25), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n480), .B2(G139), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT96), .Z(new_n801));
  NOR2_X1   g376(.A1(new_n801), .A2(new_n736), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n736), .B2(G33), .ZN(new_n803));
  INV_X1    g378(.A(G2072), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n753), .A2(G1961), .ZN(new_n807));
  NOR2_X1   g382(.A1(G168), .A2(new_n701), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n701), .B2(G21), .ZN(new_n809));
  INV_X1    g384(.A(G1966), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n810), .B2(new_n809), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n790), .A2(new_n805), .A3(new_n806), .A4(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n741), .A2(new_n784), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n723), .A2(new_n735), .A3(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NOR2_X1   g391(.A1(new_n611), .A2(new_n619), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n537), .A2(G93), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n531), .A2(G55), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n535), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n819), .B(new_n820), .C1(new_n525), .C2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(new_n563), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n563), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n818), .B(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(KEYINPUT39), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n827), .A2(new_n828), .A3(G860), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n822), .A2(G860), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT37), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n829), .A2(new_n831), .ZN(G145));
  NAND2_X1  g407(.A1(new_n516), .A2(new_n521), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n774), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n763), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n801), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n835), .A2(new_n800), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n837), .A2(KEYINPUT104), .A3(new_n801), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n694), .B(new_n626), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n480), .A2(G142), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT105), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n501), .A2(G130), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n464), .A2(G118), .ZN(new_n848));
  OAI21_X1  g423(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n844), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(G160), .B(new_n635), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(G162), .Z(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n843), .B2(new_n852), .ZN(new_n856));
  AOI21_X1  g431(.A(G37), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n852), .A2(KEYINPUT106), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n843), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n843), .A2(new_n858), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n860), .A3(new_n855), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n857), .A2(KEYINPUT40), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(KEYINPUT40), .B1(new_n857), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(G395));
  XNOR2_X1  g439(.A(G288), .B(new_n714), .ZN(new_n865));
  XNOR2_X1  g440(.A(G166), .B(G290), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(KEYINPUT42), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(KEYINPUT42), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n621), .B(new_n825), .Z(new_n874));
  NOR2_X1   g449(.A1(new_n612), .A2(new_n616), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n611), .A2(G299), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(KEYINPUT41), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n875), .B2(new_n876), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n878), .B1(new_n874), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n873), .B(new_n883), .ZN(new_n884));
  MUX2_X1   g459(.A(new_n822), .B(new_n884), .S(G868), .Z(G295));
  MUX2_X1   g460(.A(new_n822), .B(new_n884), .S(G868), .Z(G331));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n887));
  OR3_X1    g462(.A1(new_n867), .A2(new_n868), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n867), .B2(new_n868), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n823), .A2(G301), .A3(new_n824), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G301), .B1(new_n823), .B2(new_n824), .ZN(new_n893));
  OAI21_X1  g468(.A(G286), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(G168), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n877), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n879), .A2(new_n894), .A3(new_n881), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n898), .B1(new_n897), .B2(new_n877), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n890), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(new_n869), .A3(new_n900), .A4(new_n899), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n897), .A2(new_n877), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n900), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n890), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n908), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n912), .A2(new_n905), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT110), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT43), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n903), .A2(new_n905), .A3(new_n913), .A4(new_n906), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n915), .B1(new_n922), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g498(.A(G1384), .B1(new_n516), .B2(new_n521), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n924), .A2(KEYINPUT50), .ZN(new_n925));
  INV_X1    g500(.A(G1384), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n522), .B2(new_n523), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT50), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n468), .ZN(new_n930));
  XOR2_X1   g505(.A(KEYINPUT112), .B(G40), .Z(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n493), .B1(new_n492), .B2(new_n472), .ZN(new_n933));
  AOI211_X1 g508(.A(KEYINPUT74), .B(new_n471), .C1(new_n490), .C2(new_n491), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n930), .B(new_n932), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n789), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT122), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT57), .B1(new_n577), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G299), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n577), .B(new_n583), .C1(new_n937), .C2(KEYINPUT57), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n924), .A2(KEYINPUT45), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n927), .B2(new_n943), .ZN(new_n944));
  AOI211_X1 g519(.A(new_n468), .B(new_n931), .C1(new_n487), .C2(new_n494), .ZN(new_n945));
  XNOR2_X1  g520(.A(KEYINPUT56), .B(G2072), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n936), .A2(new_n941), .A3(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n939), .A2(new_n940), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n924), .A2(KEYINPUT45), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n506), .B1(new_n484), .B2(new_n513), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n508), .A2(new_n512), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n520), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n484), .A2(G2105), .ZN(new_n956));
  INV_X1    g531(.A(G126), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT77), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n951), .B1(new_n961), .B2(KEYINPUT45), .ZN(new_n962));
  INV_X1    g537(.A(new_n946), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n962), .A2(new_n935), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n924), .A2(KEYINPUT50), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n961), .B2(KEYINPUT50), .ZN(new_n966));
  AOI21_X1  g541(.A(G1956), .B1(new_n945), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n950), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT123), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT123), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n950), .B(new_n970), .C1(new_n967), .C2(new_n964), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n949), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT60), .ZN(new_n973));
  OAI211_X1 g548(.A(KEYINPUT50), .B(new_n926), .C1(new_n522), .C2(new_n523), .ZN(new_n974));
  INV_X1    g549(.A(new_n924), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n928), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G1348), .B1(new_n945), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n935), .A2(G2067), .A3(new_n975), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n973), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n945), .A2(new_n977), .ZN(new_n981));
  INV_X1    g556(.A(G1348), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n935), .A2(new_n975), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n981), .A2(new_n982), .B1(new_n983), .B2(new_n776), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n611), .B1(new_n984), .B2(KEYINPUT60), .ZN(new_n985));
  NOR4_X1   g560(.A1(new_n978), .A2(new_n979), .A3(new_n973), .A4(new_n612), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n980), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n968), .A2(new_n948), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT61), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n962), .A2(G1996), .A3(new_n935), .ZN(new_n991));
  XNOR2_X1  g566(.A(KEYINPUT58), .B(G1341), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n945), .B2(new_n924), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n564), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n995), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n564), .B(new_n997), .C1(new_n991), .C2(new_n993), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n972), .A2(new_n987), .A3(new_n990), .A4(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n969), .B(new_n971), .C1(new_n611), .C2(new_n984), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n948), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT119), .B(G2084), .Z(new_n1005));
  NAND3_X1  g580(.A1(new_n945), .A2(new_n977), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n975), .A2(new_n943), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n927), .B2(new_n943), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n810), .B1(new_n1010), .B2(new_n935), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n945), .A2(new_n977), .A3(KEYINPUT120), .A4(new_n1005), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1008), .A2(G168), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1013), .A2(new_n1014), .A3(G8), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n935), .B1(new_n976), .B2(new_n974), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT120), .B1(new_n1017), .B2(new_n1005), .ZN(new_n1018));
  OAI21_X1  g593(.A(G286), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(G8), .A3(new_n1013), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(KEYINPUT51), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n962), .B2(new_n935), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT114), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT53), .B1(new_n1025), .B2(new_n782), .ZN(new_n1026));
  INV_X1    g601(.A(G1961), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n981), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1010), .A2(new_n935), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(G171), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G40), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n942), .A2(new_n1033), .A3(new_n1030), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n924), .A2(KEYINPUT111), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n943), .B1(new_n924), .B2(KEYINPUT111), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1034), .B(G160), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1028), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(G2078), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1039), .B(G301), .C1(KEYINPUT53), .C2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT54), .B1(new_n1032), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1023), .A2(new_n1024), .A3(new_n710), .ZN(new_n1043));
  INV_X1    g618(.A(G2090), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1017), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G303), .A2(G8), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  NAND4_X1  g626(.A1(G303), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(G8), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n945), .A2(new_n924), .ZN(new_n1055));
  INV_X1    g630(.A(G1976), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(G288), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n587), .A2(G1976), .A3(new_n589), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1055), .A2(G8), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(G305), .A2(G1981), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1055), .A2(new_n1067), .A3(G8), .A4(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1058), .B(G8), .C1(new_n935), .C2(new_n975), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1059), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n929), .B2(new_n935), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n945), .A2(new_n966), .A3(KEYINPUT118), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1044), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1076), .B1(new_n1080), .B2(new_n1043), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1054), .B(new_n1075), .C1(new_n1081), .C2(new_n1053), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1021), .A2(new_n1042), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1026), .B2(new_n1038), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1039), .B(KEYINPUT126), .C1(KEYINPUT53), .C2(new_n1040), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(G171), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1087), .B(KEYINPUT54), .C1(G171), .C2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1000), .A2(new_n1090), .A3(new_n1002), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1004), .A2(new_n1083), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1071), .A2(new_n1056), .A3(new_n703), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n1065), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(KEYINPUT117), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1055), .A2(G8), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1095), .B2(KEYINPUT117), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1054), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1096), .A2(new_n1098), .B1(new_n1099), .B2(new_n1075), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1053), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1080), .A2(new_n1043), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n1076), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1076), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1074), .B1(new_n1104), .B2(new_n1053), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1106), .A2(new_n1076), .A3(G286), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT63), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G286), .A2(new_n1076), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT63), .B(new_n1111), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1104), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1101), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n1114), .A2(new_n1105), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1093), .B(new_n1100), .C1(new_n1110), .C2(new_n1115), .ZN(new_n1116));
  AOI22_X1  g691(.A1(new_n1108), .A2(new_n1109), .B1(new_n1105), .B2(new_n1114), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1099), .A2(new_n1075), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT121), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1021), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1082), .A2(new_n1032), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1021), .A2(new_n1122), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1092), .A2(new_n1116), .A3(new_n1121), .A4(new_n1126), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n935), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n694), .B(new_n696), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT113), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n774), .B(new_n776), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n763), .A2(G1996), .ZN(new_n1132));
  INV_X1    g707(.A(G1996), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n764), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1128), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G290), .B(G1986), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1128), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1127), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1128), .A2(new_n1135), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n696), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n694), .A2(new_n1143), .ZN(new_n1144));
  OAI22_X1  g719(.A1(new_n1142), .A2(new_n1144), .B1(G2067), .B2(new_n774), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1128), .B1(new_n1145), .B2(KEYINPUT127), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(KEYINPUT127), .B2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT46), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1128), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1131), .A2(new_n764), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT47), .Z(new_n1153));
  OR3_X1    g728(.A1(new_n1150), .A2(G1986), .A3(G290), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT48), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1137), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1147), .B(new_n1153), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1140), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g734(.A1(new_n857), .A2(new_n861), .ZN(new_n1161));
  NAND2_X1  g735(.A1(new_n908), .A2(new_n914), .ZN(new_n1162));
  NOR4_X1   g736(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1163));
  NAND3_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(G225));
  INV_X1    g738(.A(G225), .ZN(G308));
endmodule


