

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753;

  INV_X2 U374 ( .A(G953), .ZN(n748) );
  XNOR2_X2 U375 ( .A(G128), .B(G110), .ZN(n390) );
  NOR2_X1 U376 ( .A1(n637), .A2(G902), .ZN(n383) );
  XNOR2_X1 U377 ( .A(n369), .B(n397), .ZN(n617) );
  INV_X1 U378 ( .A(n468), .ZN(n386) );
  OR2_X1 U379 ( .A1(n697), .A2(n513), .ZN(n501) );
  OR2_X1 U380 ( .A1(n584), .A2(n565), .ZN(n567) );
  NOR2_X1 U381 ( .A1(n552), .A2(n355), .ZN(n368) );
  XNOR2_X1 U382 ( .A(n512), .B(n511), .ZN(n552) );
  XNOR2_X1 U383 ( .A(n473), .B(n472), .ZN(n517) );
  NAND2_X1 U384 ( .A1(n617), .A2(n471), .ZN(n405) );
  XNOR2_X2 U385 ( .A(n551), .B(n550), .ZN(n681) );
  AND2_X2 U386 ( .A1(n547), .A2(n546), .ZN(n657) );
  OR2_X1 U387 ( .A1(n577), .A2(n588), .ZN(n548) );
  XNOR2_X2 U388 ( .A(n475), .B(n374), .ZN(n739) );
  XNOR2_X2 U389 ( .A(n526), .B(KEYINPUT1), .ZN(n549) );
  INV_X1 U390 ( .A(n615), .ZN(n363) );
  OR2_X1 U391 ( .A1(n520), .A2(n685), .ZN(n431) );
  INV_X1 U392 ( .A(KEYINPUT101), .ZN(n458) );
  XNOR2_X1 U393 ( .A(n509), .B(n508), .ZN(n510) );
  INV_X1 U394 ( .A(KEYINPUT4), .ZN(n374) );
  XNOR2_X1 U395 ( .A(n595), .B(KEYINPUT45), .ZN(n659) );
  INV_X1 U396 ( .A(n507), .ZN(n508) );
  XNOR2_X1 U397 ( .A(n489), .B(KEYINPUT105), .ZN(n683) );
  XNOR2_X1 U398 ( .A(n426), .B(n425), .ZN(n520) );
  XNOR2_X1 U399 ( .A(KEYINPUT3), .B(G119), .ZN(n414) );
  XNOR2_X1 U400 ( .A(n368), .B(n360), .ZN(n584) );
  XNOR2_X1 U401 ( .A(n461), .B(n460), .ZN(n470) );
  XNOR2_X1 U402 ( .A(n609), .B(KEYINPUT86), .ZN(n648) );
  AND2_X1 U403 ( .A1(n546), .A2(n597), .ZN(n353) );
  AND2_X1 U404 ( .A1(n614), .A2(KEYINPUT44), .ZN(n354) );
  AND2_X1 U405 ( .A1(n556), .A2(n555), .ZN(n355) );
  XOR2_X1 U406 ( .A(n416), .B(n380), .Z(n356) );
  AND2_X1 U407 ( .A1(n536), .A2(n535), .ZN(n357) );
  AND2_X1 U408 ( .A1(n623), .A2(n354), .ZN(n358) );
  INV_X1 U409 ( .A(G902), .ZN(n471) );
  XOR2_X1 U410 ( .A(n454), .B(KEYINPUT39), .Z(n359) );
  XOR2_X1 U411 ( .A(KEYINPUT70), .B(KEYINPUT0), .Z(n360) );
  INV_X1 U412 ( .A(n721), .ZN(n370) );
  XOR2_X1 U413 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n361) );
  NAND2_X1 U414 ( .A1(n364), .A2(n362), .ZN(n594) );
  NAND2_X1 U415 ( .A1(n363), .A2(n358), .ZN(n362) );
  AND2_X1 U416 ( .A1(n367), .A2(n365), .ZN(n364) );
  NAND2_X1 U417 ( .A1(n366), .A2(n576), .ZN(n365) );
  NAND2_X1 U418 ( .A1(n623), .A2(n614), .ZN(n366) );
  NAND2_X1 U419 ( .A1(n615), .A2(n576), .ZN(n367) );
  XNOR2_X2 U420 ( .A(n563), .B(n562), .ZN(n623) );
  XNOR2_X2 U421 ( .A(n575), .B(n574), .ZN(n615) );
  AND2_X1 U422 ( .A1(n547), .A2(n353), .ZN(n596) );
  INV_X1 U423 ( .A(n657), .ZN(n652) );
  INV_X1 U424 ( .A(n742), .ZN(n369) );
  NAND2_X1 U425 ( .A1(n486), .A2(n370), .ZN(n541) );
  XNOR2_X2 U426 ( .A(n455), .B(n359), .ZN(n486) );
  OR2_X2 U427 ( .A1(n643), .A2(n597), .ZN(n509) );
  XNOR2_X2 U428 ( .A(n398), .B(G902), .ZN(n597) );
  XNOR2_X1 U429 ( .A(n411), .B(KEYINPUT72), .ZN(n577) );
  XNOR2_X2 U430 ( .A(n383), .B(n382), .ZN(n526) );
  XNOR2_X2 U431 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n392) );
  XNOR2_X2 U432 ( .A(G119), .B(KEYINPUT23), .ZN(n389) );
  XNOR2_X2 U433 ( .A(KEYINPUT92), .B(KEYINPUT93), .ZN(n391) );
  XNOR2_X2 U434 ( .A(n441), .B(KEYINPUT77), .ZN(n506) );
  BUF_X1 U435 ( .A(n577), .Z(n666) );
  XNOR2_X1 U436 ( .A(n450), .B(n449), .ZN(n643) );
  XNOR2_X1 U437 ( .A(n450), .B(n356), .ZN(n637) );
  AND2_X1 U438 ( .A1(n683), .A2(n490), .ZN(n371) );
  NOR2_X1 U439 ( .A1(n513), .A2(n552), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n742) );
  BUF_X1 U442 ( .A(n520), .Z(n581) );
  NAND2_X1 U443 ( .A1(n619), .A2(n648), .ZN(n620) );
  XNOR2_X2 U444 ( .A(G143), .B(KEYINPUT65), .ZN(n373) );
  XNOR2_X2 U445 ( .A(n373), .B(G128), .ZN(n475) );
  XNOR2_X1 U446 ( .A(KEYINPUT71), .B(G101), .ZN(n375) );
  XNOR2_X2 U447 ( .A(n739), .B(n375), .ZN(n423) );
  XNOR2_X1 U448 ( .A(G110), .B(G104), .ZN(n376) );
  XNOR2_X1 U449 ( .A(n376), .B(G107), .ZN(n726) );
  XNOR2_X1 U450 ( .A(n726), .B(KEYINPUT75), .ZN(n377) );
  XNOR2_X2 U451 ( .A(n423), .B(n377), .ZN(n450) );
  XNOR2_X2 U452 ( .A(G134), .B(G131), .ZN(n740) );
  XNOR2_X1 U453 ( .A(n740), .B(G146), .ZN(n416) );
  NAND2_X1 U454 ( .A1(G227), .A2(n748), .ZN(n378) );
  XNOR2_X1 U455 ( .A(n378), .B(KEYINPUT78), .ZN(n379) );
  XNOR2_X1 U456 ( .A(G140), .B(G137), .ZN(n385) );
  XNOR2_X1 U457 ( .A(n379), .B(n385), .ZN(n380) );
  INV_X1 U458 ( .A(KEYINPUT74), .ZN(n381) );
  XOR2_X1 U459 ( .A(n381), .B(G469), .Z(n382) );
  XNOR2_X2 U460 ( .A(G146), .B(G125), .ZN(n447) );
  INV_X1 U461 ( .A(KEYINPUT10), .ZN(n384) );
  XNOR2_X1 U462 ( .A(n447), .B(n384), .ZN(n468) );
  XNOR2_X1 U463 ( .A(KEYINPUT73), .B(KEYINPUT8), .ZN(n388) );
  NAND2_X1 U464 ( .A1(n748), .A2(G234), .ZN(n387) );
  XNOR2_X1 U465 ( .A(n388), .B(n387), .ZN(n474) );
  NAND2_X1 U466 ( .A1(n474), .A2(G221), .ZN(n396) );
  XNOR2_X1 U467 ( .A(n390), .B(n389), .ZN(n394) );
  XNOR2_X1 U468 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U469 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U470 ( .A(n396), .B(n395), .ZN(n397) );
  INV_X1 U471 ( .A(KEYINPUT15), .ZN(n398) );
  INV_X1 U472 ( .A(G234), .ZN(n399) );
  OR2_X2 U473 ( .A1(n597), .A2(n399), .ZN(n400) );
  XNOR2_X1 U474 ( .A(n400), .B(KEYINPUT20), .ZN(n406) );
  NAND2_X1 U475 ( .A1(n406), .A2(G217), .ZN(n403) );
  XNOR2_X1 U476 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n401) );
  XNOR2_X1 U477 ( .A(n401), .B(KEYINPUT25), .ZN(n402) );
  XNOR2_X1 U478 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X2 U479 ( .A(n405), .B(n404), .ZN(n494) );
  INV_X1 U480 ( .A(n406), .ZN(n408) );
  INV_X1 U481 ( .A(G221), .ZN(n407) );
  OR2_X2 U482 ( .A1(n408), .A2(n407), .ZN(n410) );
  XNOR2_X1 U483 ( .A(KEYINPUT96), .B(KEYINPUT21), .ZN(n409) );
  XNOR2_X2 U484 ( .A(n410), .B(n409), .ZN(n669) );
  XNOR2_X1 U485 ( .A(n669), .B(KEYINPUT97), .ZN(n564) );
  NAND2_X1 U486 ( .A1(n494), .A2(n564), .ZN(n411) );
  NOR2_X1 U487 ( .A1(n526), .A2(n577), .ZN(n413) );
  INV_X1 U488 ( .A(KEYINPUT98), .ZN(n412) );
  XNOR2_X1 U489 ( .A(n413), .B(n412), .ZN(n582) );
  XNOR2_X1 U490 ( .A(G113), .B(G116), .ZN(n415) );
  XNOR2_X1 U491 ( .A(n415), .B(n414), .ZN(n443) );
  XNOR2_X1 U492 ( .A(n416), .B(n443), .ZN(n422) );
  XOR2_X1 U493 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n418) );
  XNOR2_X1 U494 ( .A(G137), .B(KEYINPUT5), .ZN(n417) );
  XNOR2_X1 U495 ( .A(n418), .B(n417), .ZN(n420) );
  NOR2_X1 U496 ( .A1(G953), .A2(G237), .ZN(n464) );
  NAND2_X1 U497 ( .A1(G210), .A2(n464), .ZN(n419) );
  XNOR2_X1 U498 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U499 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U500 ( .A(n424), .B(n423), .ZN(n625) );
  NAND2_X1 U501 ( .A1(n625), .A2(n471), .ZN(n426) );
  INV_X1 U502 ( .A(G472), .ZN(n425) );
  INV_X1 U503 ( .A(G237), .ZN(n427) );
  NAND2_X1 U504 ( .A1(n471), .A2(n427), .ZN(n451) );
  NAND2_X1 U505 ( .A1(n451), .A2(G214), .ZN(n429) );
  INV_X1 U506 ( .A(KEYINPUT88), .ZN(n428) );
  XNOR2_X1 U507 ( .A(n429), .B(n428), .ZN(n685) );
  INV_X1 U508 ( .A(KEYINPUT30), .ZN(n430) );
  XNOR2_X1 U509 ( .A(n431), .B(n430), .ZN(n439) );
  XOR2_X1 U510 ( .A(KEYINPUT14), .B(KEYINPUT89), .Z(n433) );
  NAND2_X1 U511 ( .A1(G237), .A2(G234), .ZN(n432) );
  XNOR2_X1 U512 ( .A(n433), .B(n432), .ZN(n437) );
  NAND2_X1 U513 ( .A1(G902), .A2(n437), .ZN(n554) );
  NOR2_X1 U514 ( .A1(G900), .A2(n554), .ZN(n434) );
  NAND2_X1 U515 ( .A1(G953), .A2(n434), .ZN(n436) );
  INV_X1 U516 ( .A(KEYINPUT107), .ZN(n435) );
  XNOR2_X1 U517 ( .A(n436), .B(n435), .ZN(n438) );
  AND2_X1 U518 ( .A1(n437), .A2(G952), .ZN(n695) );
  NAND2_X1 U519 ( .A1(n695), .A2(n748), .ZN(n556) );
  NAND2_X1 U520 ( .A1(n438), .A2(n556), .ZN(n495) );
  NAND2_X1 U521 ( .A1(n439), .A2(n495), .ZN(n440) );
  OR2_X2 U522 ( .A1(n582), .A2(n440), .ZN(n441) );
  XNOR2_X1 U523 ( .A(KEYINPUT16), .B(G122), .ZN(n442) );
  XNOR2_X1 U524 ( .A(n443), .B(n442), .ZN(n728) );
  XNOR2_X1 U525 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n445) );
  NAND2_X1 U526 ( .A1(n748), .A2(G224), .ZN(n444) );
  XNOR2_X1 U527 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U528 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U529 ( .A(n728), .B(n448), .ZN(n449) );
  NAND2_X1 U530 ( .A1(n451), .A2(G210), .ZN(n453) );
  INV_X1 U531 ( .A(KEYINPUT87), .ZN(n452) );
  XNOR2_X1 U532 ( .A(n453), .B(n452), .ZN(n507) );
  XNOR2_X1 U533 ( .A(n509), .B(n507), .ZN(n503) );
  XNOR2_X1 U534 ( .A(n503), .B(KEYINPUT38), .ZN(n688) );
  NAND2_X1 U535 ( .A1(n506), .A2(n688), .ZN(n455) );
  INV_X1 U536 ( .A(KEYINPUT84), .ZN(n454) );
  XOR2_X1 U537 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n457) );
  XNOR2_X1 U538 ( .A(KEYINPUT103), .B(KEYINPUT11), .ZN(n456) );
  XNOR2_X1 U539 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U540 ( .A(G143), .B(G131), .ZN(n459) );
  XOR2_X1 U541 ( .A(G122), .B(G113), .Z(n463) );
  XNOR2_X1 U542 ( .A(G140), .B(G104), .ZN(n462) );
  XNOR2_X1 U543 ( .A(n463), .B(n462), .ZN(n466) );
  NAND2_X1 U544 ( .A1(G214), .A2(n464), .ZN(n465) );
  XNOR2_X1 U545 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U546 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U547 ( .A(n470), .B(n469), .ZN(n605) );
  NAND2_X1 U548 ( .A1(n605), .A2(n471), .ZN(n473) );
  XNOR2_X1 U549 ( .A(KEYINPUT13), .B(G475), .ZN(n472) );
  NAND2_X1 U550 ( .A1(n474), .A2(G217), .ZN(n476) );
  XNOR2_X1 U551 ( .A(n476), .B(n475), .ZN(n483) );
  XOR2_X1 U552 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n478) );
  XNOR2_X1 U553 ( .A(G122), .B(G134), .ZN(n477) );
  XNOR2_X1 U554 ( .A(n478), .B(n477), .ZN(n481) );
  XNOR2_X1 U555 ( .A(G107), .B(G116), .ZN(n479) );
  XNOR2_X1 U556 ( .A(n479), .B(KEYINPUT104), .ZN(n480) );
  XNOR2_X1 U557 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U558 ( .A(n483), .B(n482), .ZN(n630) );
  OR2_X1 U559 ( .A1(n630), .A2(G902), .ZN(n484) );
  XNOR2_X1 U560 ( .A(n484), .B(G478), .ZN(n516) );
  OR2_X1 U561 ( .A1(n517), .A2(n516), .ZN(n718) );
  INV_X1 U562 ( .A(n718), .ZN(n485) );
  NAND2_X2 U563 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X2 U564 ( .A(n487), .B(KEYINPUT40), .ZN(n622) );
  INV_X1 U565 ( .A(n517), .ZN(n488) );
  OR2_X1 U566 ( .A1(n488), .A2(n516), .ZN(n489) );
  INV_X1 U567 ( .A(n685), .ZN(n490) );
  NAND2_X1 U568 ( .A1(n688), .A2(n371), .ZN(n493) );
  INV_X1 U569 ( .A(KEYINPUT108), .ZN(n491) );
  XNOR2_X1 U570 ( .A(n491), .B(KEYINPUT41), .ZN(n492) );
  XNOR2_X1 U571 ( .A(n493), .B(n492), .ZN(n697) );
  INV_X1 U572 ( .A(n669), .ZN(n496) );
  NAND2_X1 U573 ( .A1(n496), .A2(n495), .ZN(n497) );
  OR2_X1 U574 ( .A1(n494), .A2(n497), .ZN(n521) );
  NOR2_X1 U575 ( .A1(n581), .A2(n521), .ZN(n499) );
  INV_X1 U576 ( .A(KEYINPUT28), .ZN(n498) );
  XNOR2_X1 U577 ( .A(n499), .B(n498), .ZN(n500) );
  OR2_X1 U578 ( .A1(n500), .A2(n526), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n501), .B(KEYINPUT42), .ZN(n616) );
  NAND2_X1 U580 ( .A1(n622), .A2(n616), .ZN(n502) );
  XNOR2_X1 U581 ( .A(n502), .B(n361), .ZN(n537) );
  INV_X1 U582 ( .A(n516), .ZN(n504) );
  OR2_X1 U583 ( .A1(n517), .A2(n504), .ZN(n559) );
  NOR2_X1 U584 ( .A1(n503), .A2(n559), .ZN(n505) );
  AND2_X1 U585 ( .A1(n506), .A2(n505), .ZN(n716) );
  XNOR2_X1 U586 ( .A(n716), .B(KEYINPUT81), .ZN(n536) );
  NAND2_X1 U587 ( .A1(n510), .A2(n490), .ZN(n512) );
  XNOR2_X1 U588 ( .A(KEYINPUT69), .B(KEYINPUT19), .ZN(n511) );
  INV_X1 U589 ( .A(KEYINPUT47), .ZN(n514) );
  NAND2_X1 U590 ( .A1(n372), .A2(n514), .ZN(n515) );
  NAND2_X1 U591 ( .A1(n515), .A2(KEYINPUT80), .ZN(n518) );
  NAND2_X1 U592 ( .A1(n517), .A2(n516), .ZN(n721) );
  AND2_X1 U593 ( .A1(n721), .A2(n718), .ZN(n686) );
  INV_X1 U594 ( .A(n686), .ZN(n585) );
  AND2_X1 U595 ( .A1(n518), .A2(n585), .ZN(n534) );
  INV_X1 U596 ( .A(KEYINPUT6), .ZN(n519) );
  XNOR2_X1 U597 ( .A(n520), .B(n519), .ZN(n588) );
  INV_X1 U598 ( .A(n521), .ZN(n523) );
  NOR2_X1 U599 ( .A1(n685), .A2(n718), .ZN(n522) );
  NAND2_X1 U600 ( .A1(n523), .A2(n522), .ZN(n524) );
  OR2_X1 U601 ( .A1(n588), .A2(n524), .ZN(n542) );
  NOR2_X1 U602 ( .A1(n542), .A2(n503), .ZN(n525) );
  XNOR2_X1 U603 ( .A(n525), .B(KEYINPUT36), .ZN(n527) );
  INV_X1 U604 ( .A(n549), .ZN(n572) );
  AND2_X1 U605 ( .A1(n527), .A2(n572), .ZN(n723) );
  NOR2_X1 U606 ( .A1(KEYINPUT80), .A2(KEYINPUT47), .ZN(n528) );
  NOR2_X1 U607 ( .A1(n723), .A2(n528), .ZN(n532) );
  NAND2_X1 U608 ( .A1(n686), .A2(KEYINPUT80), .ZN(n529) );
  NAND2_X1 U609 ( .A1(n372), .A2(n529), .ZN(n530) );
  NAND2_X1 U610 ( .A1(n530), .A2(KEYINPUT47), .ZN(n531) );
  NAND2_X1 U611 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U612 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U613 ( .A1(n537), .A2(n357), .ZN(n539) );
  INV_X1 U614 ( .A(KEYINPUT48), .ZN(n538) );
  XNOR2_X1 U615 ( .A(n539), .B(n538), .ZN(n547) );
  INV_X1 U616 ( .A(KEYINPUT109), .ZN(n540) );
  XNOR2_X1 U617 ( .A(n541), .B(n540), .ZN(n753) );
  INV_X1 U618 ( .A(n542), .ZN(n543) );
  NAND2_X1 U619 ( .A1(n549), .A2(n543), .ZN(n544) );
  XNOR2_X1 U620 ( .A(n544), .B(KEYINPUT43), .ZN(n545) );
  NAND2_X1 U621 ( .A1(n545), .A2(n503), .ZN(n612) );
  AND2_X1 U622 ( .A1(n753), .A2(n612), .ZN(n546) );
  OR2_X2 U623 ( .A1(n549), .A2(n548), .ZN(n551) );
  INV_X1 U624 ( .A(KEYINPUT33), .ZN(n550) );
  NOR2_X1 U625 ( .A1(G898), .A2(n748), .ZN(n553) );
  XOR2_X1 U626 ( .A(KEYINPUT90), .B(n553), .Z(n729) );
  OR2_X1 U627 ( .A1(n729), .A2(n554), .ZN(n555) );
  OR2_X2 U628 ( .A1(n681), .A2(n584), .ZN(n558) );
  INV_X1 U629 ( .A(KEYINPUT34), .ZN(n557) );
  XNOR2_X1 U630 ( .A(n558), .B(n557), .ZN(n561) );
  INV_X1 U631 ( .A(n559), .ZN(n560) );
  NAND2_X1 U632 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U633 ( .A(KEYINPUT79), .B(KEYINPUT35), .ZN(n562) );
  NAND2_X1 U634 ( .A1(n683), .A2(n564), .ZN(n565) );
  INV_X1 U635 ( .A(KEYINPUT22), .ZN(n566) );
  XNOR2_X2 U636 ( .A(n567), .B(n566), .ZN(n591) );
  INV_X1 U637 ( .A(n494), .ZN(n570) );
  AND2_X1 U638 ( .A1(n581), .A2(n570), .ZN(n568) );
  AND2_X1 U639 ( .A1(n549), .A2(n568), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n591), .A2(n569), .ZN(n614) );
  XNOR2_X1 U641 ( .A(n570), .B(KEYINPUT106), .ZN(n670) );
  AND2_X1 U642 ( .A1(n588), .A2(n670), .ZN(n571) );
  AND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n591), .A2(n573), .ZN(n575) );
  XNOR2_X1 U645 ( .A(KEYINPUT67), .B(KEYINPUT32), .ZN(n574) );
  INV_X1 U646 ( .A(KEYINPUT44), .ZN(n576) );
  OR2_X1 U647 ( .A1(n549), .A2(n666), .ZN(n578) );
  OR2_X1 U648 ( .A1(n578), .A2(n581), .ZN(n677) );
  OR2_X1 U649 ( .A1(n584), .A2(n677), .ZN(n580) );
  INV_X1 U650 ( .A(KEYINPUT31), .ZN(n579) );
  XNOR2_X1 U651 ( .A(n580), .B(n579), .ZN(n720) );
  INV_X1 U652 ( .A(n581), .ZN(n672) );
  OR2_X1 U653 ( .A1(n582), .A2(n672), .ZN(n583) );
  OR2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n707) );
  NAND2_X1 U655 ( .A1(n720), .A2(n707), .ZN(n586) );
  NAND2_X1 U656 ( .A1(n586), .A2(n585), .ZN(n592) );
  INV_X1 U657 ( .A(n670), .ZN(n587) );
  AND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  AND2_X1 U659 ( .A1(n549), .A2(n589), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n613) );
  AND2_X1 U661 ( .A1(n592), .A2(n613), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n596), .A2(n659), .ZN(n600) );
  NAND2_X1 U664 ( .A1(n597), .A2(KEYINPUT2), .ZN(n598) );
  XNOR2_X1 U665 ( .A(n598), .B(KEYINPUT68), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U667 ( .A(KEYINPUT66), .B(n601), .Z(n604) );
  INV_X1 U668 ( .A(n659), .ZN(n653) );
  NAND2_X1 U669 ( .A1(n657), .A2(KEYINPUT2), .ZN(n602) );
  NOR2_X2 U670 ( .A1(n653), .A2(n602), .ZN(n603) );
  XNOR2_X1 U671 ( .A(n603), .B(KEYINPUT76), .ZN(n664) );
  NOR2_X2 U672 ( .A1(n604), .A2(n664), .ZN(n642) );
  NAND2_X1 U673 ( .A1(n642), .A2(G475), .ZN(n607) );
  XOR2_X1 U674 ( .A(n605), .B(KEYINPUT59), .Z(n606) );
  XNOR2_X1 U675 ( .A(n607), .B(n606), .ZN(n610) );
  INV_X1 U676 ( .A(G952), .ZN(n608) );
  NAND2_X1 U677 ( .A1(n608), .A2(G953), .ZN(n609) );
  AND2_X2 U678 ( .A1(n610), .A2(n648), .ZN(n611) );
  XNOR2_X1 U679 ( .A(n611), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U680 ( .A(n612), .B(G140), .ZN(G42) );
  XNOR2_X1 U681 ( .A(n613), .B(G101), .ZN(G3) );
  XNOR2_X1 U682 ( .A(n614), .B(G110), .ZN(G12) );
  XOR2_X1 U683 ( .A(n615), .B(G119), .Z(G21) );
  XNOR2_X1 U684 ( .A(n616), .B(G137), .ZN(G39) );
  NAND2_X1 U685 ( .A1(n642), .A2(G217), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U687 ( .A(n620), .B(KEYINPUT121), .ZN(G66) );
  XOR2_X1 U688 ( .A(G131), .B(KEYINPUT127), .Z(n621) );
  XNOR2_X1 U689 ( .A(n622), .B(n621), .ZN(G33) );
  XNOR2_X1 U690 ( .A(G122), .B(KEYINPUT126), .ZN(n624) );
  XNOR2_X1 U691 ( .A(n623), .B(n624), .ZN(G24) );
  NAND2_X1 U692 ( .A1(n642), .A2(G472), .ZN(n627) );
  XNOR2_X1 U693 ( .A(n625), .B(KEYINPUT62), .ZN(n626) );
  XNOR2_X1 U694 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U695 ( .A1(n628), .A2(n648), .ZN(n629) );
  XNOR2_X1 U696 ( .A(n629), .B(KEYINPUT63), .ZN(G57) );
  BUF_X1 U697 ( .A(n642), .Z(n634) );
  NAND2_X1 U698 ( .A1(n634), .A2(G478), .ZN(n632) );
  XNOR2_X1 U699 ( .A(n630), .B(KEYINPUT120), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n632), .B(n631), .ZN(n633) );
  INV_X1 U701 ( .A(n648), .ZN(n640) );
  NOR2_X1 U702 ( .A1(n633), .A2(n640), .ZN(G63) );
  NAND2_X1 U703 ( .A1(n634), .A2(G469), .ZN(n639) );
  XNOR2_X1 U704 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n635) );
  XNOR2_X1 U705 ( .A(n635), .B(KEYINPUT58), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n641) );
  NOR2_X1 U708 ( .A1(n641), .A2(n640), .ZN(G54) );
  NAND2_X1 U709 ( .A1(n642), .A2(G210), .ZN(n647) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n644) );
  XOR2_X1 U711 ( .A(n644), .B(KEYINPUT55), .Z(n645) );
  XNOR2_X1 U712 ( .A(n643), .B(n645), .ZN(n646) );
  XNOR2_X1 U713 ( .A(n647), .B(n646), .ZN(n649) );
  NAND2_X1 U714 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U715 ( .A(KEYINPUT83), .B(KEYINPUT56), .ZN(n650) );
  XNOR2_X1 U716 ( .A(n651), .B(n650), .ZN(G51) );
  NOR2_X1 U717 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U718 ( .A1(n654), .A2(KEYINPUT2), .ZN(n656) );
  INV_X1 U719 ( .A(KEYINPUT82), .ZN(n655) );
  NOR2_X1 U720 ( .A1(n656), .A2(n655), .ZN(n663) );
  NOR2_X1 U721 ( .A1(KEYINPUT2), .A2(KEYINPUT82), .ZN(n658) );
  NAND2_X1 U722 ( .A1(n657), .A2(n658), .ZN(n661) );
  BUF_X1 U723 ( .A(n659), .Z(n660) );
  NOR2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n665) );
  NOR2_X1 U726 ( .A1(n665), .A2(n664), .ZN(n703) );
  NAND2_X1 U727 ( .A1(n549), .A2(n666), .ZN(n668) );
  XOR2_X1 U728 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n667) );
  XNOR2_X1 U729 ( .A(n668), .B(n667), .ZN(n676) );
  NAND2_X1 U730 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U731 ( .A(n671), .B(KEYINPUT49), .ZN(n673) );
  NOR2_X1 U732 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U733 ( .A(n674), .B(KEYINPUT116), .ZN(n675) );
  NAND2_X1 U734 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U735 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n679), .B(KEYINPUT51), .ZN(n680) );
  NOR2_X1 U737 ( .A1(n680), .A2(n697), .ZN(n693) );
  INV_X1 U738 ( .A(n688), .ZN(n682) );
  NAND2_X1 U739 ( .A1(n682), .A2(n685), .ZN(n684) );
  NAND2_X1 U740 ( .A1(n684), .A2(n683), .ZN(n690) );
  NOR2_X1 U741 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U742 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U743 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U744 ( .A1(n681), .A2(n691), .ZN(n692) );
  NOR2_X1 U745 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U746 ( .A(KEYINPUT52), .B(n694), .Z(n696) );
  NAND2_X1 U747 ( .A1(n696), .A2(n695), .ZN(n701) );
  NOR2_X1 U748 ( .A1(n681), .A2(n697), .ZN(n698) );
  XNOR2_X1 U749 ( .A(n698), .B(KEYINPUT118), .ZN(n699) );
  NOR2_X1 U750 ( .A1(n699), .A2(G953), .ZN(n700) );
  NAND2_X1 U751 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U752 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U753 ( .A(n704), .B(KEYINPUT53), .ZN(G75) );
  NOR2_X1 U754 ( .A1(n707), .A2(n718), .ZN(n705) );
  XOR2_X1 U755 ( .A(KEYINPUT110), .B(n705), .Z(n706) );
  XNOR2_X1 U756 ( .A(G104), .B(n706), .ZN(G6) );
  NOR2_X1 U757 ( .A1(n707), .A2(n721), .ZN(n712) );
  XOR2_X1 U758 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n709) );
  XNOR2_X1 U759 ( .A(G107), .B(KEYINPUT26), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U761 ( .A(KEYINPUT111), .B(n710), .ZN(n711) );
  XNOR2_X1 U762 ( .A(n712), .B(n711), .ZN(G9) );
  XOR2_X1 U763 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n714) );
  NAND2_X1 U764 ( .A1(n372), .A2(n370), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U766 ( .A(G128), .B(n715), .Z(G30) );
  XOR2_X1 U767 ( .A(G143), .B(n716), .Z(G45) );
  NAND2_X1 U768 ( .A1(n372), .A2(n485), .ZN(n717) );
  XNOR2_X1 U769 ( .A(n717), .B(G146), .ZN(G48) );
  NOR2_X1 U770 ( .A1(n718), .A2(n720), .ZN(n719) );
  XOR2_X1 U771 ( .A(G113), .B(n719), .Z(G15) );
  NOR2_X1 U772 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U773 ( .A(G116), .B(n722), .Z(G18) );
  XNOR2_X1 U774 ( .A(n723), .B(KEYINPUT114), .ZN(n724) );
  XNOR2_X1 U775 ( .A(n724), .B(KEYINPUT37), .ZN(n725) );
  XNOR2_X1 U776 ( .A(G125), .B(n725), .ZN(G27) );
  XOR2_X1 U777 ( .A(G101), .B(n726), .Z(n727) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n730), .A2(n729), .ZN(n737) );
  NAND2_X1 U780 ( .A1(n660), .A2(n748), .ZN(n731) );
  XNOR2_X1 U781 ( .A(n731), .B(KEYINPUT122), .ZN(n735) );
  NAND2_X1 U782 ( .A1(G953), .A2(G224), .ZN(n732) );
  XNOR2_X1 U783 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U784 ( .A1(n733), .A2(G898), .ZN(n734) );
  NAND2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(KEYINPUT123), .B(n738), .ZN(G69) );
  XNOR2_X1 U788 ( .A(n739), .B(n740), .ZN(n741) );
  XOR2_X1 U789 ( .A(n742), .B(n741), .Z(n746) );
  XNOR2_X1 U790 ( .A(G227), .B(n746), .ZN(n743) );
  NAND2_X1 U791 ( .A1(n743), .A2(G900), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(G953), .ZN(n745) );
  XOR2_X1 U793 ( .A(KEYINPUT125), .B(n745), .Z(n751) );
  XNOR2_X1 U794 ( .A(n746), .B(KEYINPUT124), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n652), .B(n747), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U797 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U798 ( .A(G134), .B(KEYINPUT115), .Z(n752) );
  XNOR2_X1 U799 ( .A(n753), .B(n752), .ZN(G36) );
endmodule

