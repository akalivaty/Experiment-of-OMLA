//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT2), .ZN(new_n207));
  OR2_X1    g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211));
  INV_X1    g010(.A(new_n206), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(KEYINPUT83), .A3(new_n206), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n206), .B1(new_n217), .B2(KEYINPUT2), .ZN(new_n220));
  INV_X1    g019(.A(new_n209), .ZN(new_n221));
  NOR2_X1   g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT84), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT84), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n224), .A3(new_n209), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n220), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT29), .ZN(new_n230));
  INV_X1    g029(.A(G218gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G211gat), .ZN(new_n232));
  INV_X1    g031(.A(G211gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G218gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n232), .B2(new_n234), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT22), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT80), .B(G211gat), .Z(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(new_n231), .ZN(new_n241));
  INV_X1    g040(.A(G197gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT79), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT79), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G197gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n245), .A3(G204gat), .ZN(new_n246));
  INV_X1    g045(.A(G204gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n244), .A2(G197gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n242), .A2(KEYINPUT79), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n238), .A2(new_n241), .A3(new_n246), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n246), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT80), .B(G211gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT22), .B1(new_n253), .B2(G218gat), .ZN(new_n254));
  OAI22_X1  g053(.A1(new_n252), .A2(new_n254), .B1(new_n237), .B2(new_n236), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n229), .A2(new_n230), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n219), .A2(new_n226), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g057(.A1(G228gat), .A2(G233gat), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n251), .A2(new_n255), .A3(new_n230), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n227), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G22gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT86), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n251), .A2(new_n255), .A3(KEYINPUT86), .A4(new_n230), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n228), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n256), .B1(new_n269), .B2(new_n257), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n264), .B(new_n265), .C1(new_n270), .C2(new_n260), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT3), .B1(new_n263), .B2(new_n266), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n227), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n259), .B1(new_n274), .B2(new_n256), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n265), .B1(new_n275), .B2(new_n264), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n272), .A2(new_n276), .A3(G78gat), .ZN(new_n277));
  INV_X1    g076(.A(G78gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n264), .B1(new_n270), .B2(new_n260), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G22gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n278), .B1(new_n280), .B2(new_n271), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n205), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(G78gat), .B1(new_n272), .B2(new_n276), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n278), .A3(new_n271), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n204), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G113gat), .B(G120gat), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT73), .B(G134gat), .C1(new_n287), .C2(KEYINPUT1), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n289));
  INV_X1    g088(.A(G134gat), .ZN(new_n290));
  INV_X1    g089(.A(G113gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(G120gat), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G113gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n289), .B(new_n290), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G127gat), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n288), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(new_n288), .B2(new_n295), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT74), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n299), .A2(KEYINPUT74), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT24), .ZN(new_n303));
  INV_X1    g102(.A(G183gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(G183gat), .A3(G190gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n302), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G183gat), .B(G190gat), .ZN(new_n312));
  OAI211_X1 g111(.A(KEYINPUT64), .B(new_n309), .C1(new_n312), .C2(new_n303), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT65), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G169gat), .ZN(new_n318));
  INV_X1    g117(.A(G176gat), .ZN(new_n319));
  AND4_X1   g118(.A1(KEYINPUT23), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT66), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NOR3_X1   g127(.A1(new_n320), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT25), .B1(new_n314), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n319), .A3(KEYINPUT23), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n327), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT25), .A4(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(new_n326), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n306), .A2(G183gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n304), .A2(G190gat), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT24), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT68), .B1(new_n339), .B2(new_n309), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n308), .A2(new_n341), .A3(new_n310), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n336), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT69), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n341), .B1(new_n308), .B2(new_n310), .ZN(new_n345));
  OAI211_X1 g144(.A(KEYINPUT68), .B(new_n309), .C1(new_n312), .C2(new_n303), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT69), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n336), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n330), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT26), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n327), .B1(new_n321), .B2(new_n351), .ZN(new_n352));
  NOR3_X1   g151(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n353));
  OAI22_X1  g152(.A1(new_n352), .A2(new_n353), .B1(new_n304), .B2(new_n306), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT72), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n304), .A2(KEYINPUT27), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(G183gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT28), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT70), .B1(new_n356), .B2(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n357), .A2(G183gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT70), .ZN(new_n365));
  AOI21_X1  g164(.A(G190gat), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT28), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT71), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n362), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n355), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n300), .B(new_n301), .C1(new_n350), .C2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n314), .A2(new_n329), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT25), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n347), .A2(new_n348), .A3(new_n336), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n348), .B1(new_n347), .B2(new_n336), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n354), .B(KEYINPUT72), .Z(new_n382));
  INV_X1    g181(.A(new_n371), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(new_n369), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n381), .A2(new_n384), .A3(KEYINPUT74), .A4(new_n299), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n373), .A2(new_n375), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(KEYINPUT32), .ZN(new_n389));
  XOR2_X1   g188(.A(G15gat), .B(G43gat), .Z(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT75), .ZN(new_n391));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(KEYINPUT33), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n386), .A2(KEYINPUT32), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(KEYINPUT76), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n373), .A2(new_n385), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT34), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n374), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT78), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n398), .A2(new_n402), .A3(new_n399), .A4(new_n374), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n374), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT34), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT76), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n388), .A2(new_n389), .A3(new_n407), .A4(new_n393), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n397), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n406), .B1(new_n397), .B2(new_n408), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n286), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT0), .ZN(new_n413));
  XNOR2_X1  g212(.A(G57gat), .B(G85gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  OAI21_X1  g214(.A(new_n227), .B1(new_n297), .B2(new_n298), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n299), .A2(new_n229), .A3(new_n258), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT4), .B(new_n227), .C1(new_n297), .C2(new_n298), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n288), .A2(new_n295), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G127gat), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n288), .A2(new_n295), .A3(new_n296), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n257), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n416), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n422), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n299), .A2(KEYINPUT85), .A3(new_n257), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n421), .A2(new_n422), .B1(new_n431), .B2(KEYINPUT5), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n418), .A2(new_n419), .A3(new_n422), .A4(new_n420), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n415), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n433), .ZN(new_n439));
  INV_X1    g238(.A(new_n415), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n421), .A2(KEYINPUT5), .A3(new_n422), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n441), .A4(new_n440), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n251), .A2(new_n255), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G226gat), .ZN(new_n448));
  INV_X1    g247(.A(G233gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n450), .A2(KEYINPUT29), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n350), .B2(new_n372), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n381), .A2(new_n384), .A3(KEYINPUT82), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n381), .A2(new_n384), .A3(new_n450), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n447), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n450), .A3(new_n455), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n451), .B1(new_n350), .B2(new_n372), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n446), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G8gat), .B(G36gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  AND3_X1   g264(.A1(new_n459), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n459), .B2(new_n462), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n459), .A2(new_n462), .A3(new_n468), .A4(new_n465), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n445), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT88), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT35), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n443), .A2(new_n444), .ZN(new_n475));
  INV_X1    g274(.A(new_n465), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n350), .A2(new_n372), .A3(new_n453), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT82), .B1(new_n381), .B2(new_n384), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n451), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n446), .B1(new_n479), .B2(new_n457), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n460), .A2(new_n446), .A3(new_n461), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n459), .A2(new_n462), .A3(new_n465), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(KEYINPUT30), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n475), .B1(new_n484), .B2(new_n470), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n411), .A2(new_n473), .A3(new_n474), .A4(new_n487), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n396), .A2(KEYINPUT76), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n408), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT77), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n492), .A3(new_n406), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n406), .A2(new_n492), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n397), .A3(new_n408), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n277), .A2(new_n281), .A3(new_n205), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n204), .B1(new_n283), .B2(new_n284), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n485), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n488), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n446), .B1(new_n456), .B2(new_n458), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n460), .A2(new_n447), .A3(new_n461), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT37), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT38), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n465), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n506), .C1(new_n467), .C2(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n443), .A2(new_n444), .A3(new_n483), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n507), .B1(new_n459), .B2(new_n462), .ZN(new_n511));
  INV_X1    g310(.A(new_n508), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n482), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n509), .B(new_n510), .C1(new_n513), .C2(new_n506), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n429), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n428), .A2(new_n430), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n422), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n518), .A3(KEYINPUT39), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(new_n415), .C1(KEYINPUT39), .C2(new_n516), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT40), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n442), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n519), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n415), .B1(new_n516), .B2(KEYINPUT39), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n520), .A2(new_n527), .A3(new_n521), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n529), .A2(new_n484), .A3(new_n470), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n530), .A3(new_n499), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n493), .A2(new_n495), .A3(KEYINPUT36), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n399), .B1(new_n398), .B2(new_n374), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(KEYINPUT78), .B2(new_n400), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n491), .A2(new_n403), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT36), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n397), .A2(new_n406), .A3(new_n408), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n472), .A2(new_n286), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n531), .A2(new_n532), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n502), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NAND3_X1  g344(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT14), .ZN(new_n549));
  INV_X1    g348(.A(G29gat), .ZN(new_n550));
  INV_X1    g349(.A(G36gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n548), .B1(KEYINPUT89), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(KEYINPUT89), .B2(new_n552), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n550), .B2(new_n551), .ZN(new_n555));
  XOR2_X1   g354(.A(G43gat), .B(G50gat), .Z(new_n556));
  INV_X1    g355(.A(KEYINPUT15), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n556), .A2(new_n557), .B1(new_n552), .B2(new_n547), .ZN(new_n560));
  OAI221_X1 g359(.A(new_n560), .B1(new_n557), .B2(new_n556), .C1(new_n550), .C2(new_n551), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT7), .ZN(new_n564));
  NAND2_X1  g363(.A1(G99gat), .A2(G106gat), .ZN(new_n565));
  INV_X1    g364(.A(G85gat), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G99gat), .B(G106gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n546), .B1(new_n562), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT96), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n571), .B(KEYINPUT95), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n577), .B1(new_n562), .B2(KEYINPUT90), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n561), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT90), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT17), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n576), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n544), .B(new_n545), .C1(new_n574), .C2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n572), .B(KEYINPUT96), .ZN(new_n584));
  INV_X1    g383(.A(new_n582), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(new_n585), .A3(new_n543), .A4(new_n542), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(KEYINPUT99), .A3(new_n591), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n583), .A2(new_n586), .A3(new_n590), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT98), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n583), .A2(new_n586), .A3(new_n598), .A4(new_n590), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n594), .A2(new_n595), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G57gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(G64gat), .ZN(new_n602));
  INV_X1    g401(.A(G64gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(G57gat), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n605));
  OAI22_X1  g404(.A1(new_n602), .A2(new_n604), .B1(new_n605), .B2(KEYINPUT9), .ZN(new_n606));
  NOR2_X1   g405(.A1(G71gat), .A2(G78gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n607), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n606), .B(new_n609), .C1(new_n605), .C2(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(KEYINPUT9), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n608), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT94), .B1(new_n601), .B2(G64gat), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(G57gat), .B2(new_n603), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n601), .A2(KEYINPUT94), .A3(G64gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(new_n296), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n622));
  XNOR2_X1  g421(.A(G15gat), .B(G22gat), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT16), .ZN(new_n624));
  OAI21_X1  g423(.A(KEYINPUT91), .B1(new_n624), .B2(G1gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n624), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n627));
  OAI221_X1 g426(.A(new_n622), .B1(G1gat), .B2(new_n623), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(G8gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(G8gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(KEYINPUT21), .B2(new_n617), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n621), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(new_n215), .ZN(new_n635));
  XOR2_X1   g434(.A(G183gat), .B(G211gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n633), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n600), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n562), .B(new_n631), .ZN(new_n640));
  NAND2_X1  g439(.A1(G229gat), .A2(G233gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(KEYINPUT13), .Z(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n631), .B1(new_n578), .B2(new_n581), .ZN(new_n645));
  INV_X1    g444(.A(new_n631), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n562), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n641), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT18), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(G197gat), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT11), .B(G169gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT12), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n651), .B(new_n657), .C1(new_n650), .C2(new_n649), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n649), .A2(new_n650), .ZN(new_n659));
  INV_X1    g458(.A(new_n641), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n645), .A2(new_n660), .A3(new_n647), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n661), .A2(KEYINPUT18), .B1(new_n640), .B2(new_n643), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n656), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n571), .B(new_n617), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n617), .ZN(new_n671));
  OR3_X1    g470(.A1(new_n671), .A2(new_n667), .A3(new_n571), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n666), .A2(KEYINPUT100), .A3(new_n667), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n666), .A2(new_n675), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G120gat), .B(G148gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  OR2_X1    g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n676), .A2(new_n677), .A3(new_n681), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n639), .A2(new_n665), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n541), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n475), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g487(.A1(new_n484), .A2(new_n470), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT16), .B(G8gat), .Z(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n686), .ZN(new_n693));
  OAI21_X1  g492(.A(G8gat), .B1(new_n693), .B2(new_n689), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n692), .ZN(new_n695));
  MUX2_X1   g494(.A(new_n692), .B(new_n695), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g495(.A1(new_n538), .A2(new_n532), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G15gat), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n535), .A2(new_n537), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n700), .A2(G15gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n693), .B2(new_n701), .ZN(G1326gat));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n286), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT43), .B(G22gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  NAND2_X1  g504(.A1(new_n597), .A2(new_n599), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT99), .B1(new_n587), .B2(new_n591), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n593), .B(new_n590), .C1(new_n583), .C2(new_n586), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n689), .A2(new_n486), .A3(new_n445), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n486), .B1(new_n689), .B2(new_n445), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n700), .A2(KEYINPUT35), .A3(new_n286), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n712), .A2(new_n713), .B1(KEYINPUT35), .B2(new_n500), .ZN(new_n714));
  AND4_X1   g513(.A1(new_n531), .A2(new_n532), .A3(new_n538), .A4(new_n539), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n709), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n665), .A2(new_n638), .A3(new_n684), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n550), .A3(new_n475), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT45), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n709), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n594), .A2(new_n595), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT102), .B1(new_n725), .B2(new_n706), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n502), .B2(new_n540), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n600), .B1(new_n502), .B2(new_n540), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT101), .B1(new_n731), .B2(new_n728), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT101), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n733), .A3(KEYINPUT44), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n730), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(new_n718), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n722), .B1(new_n736), .B2(new_n445), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G29gat), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n736), .A2(new_n722), .A3(new_n445), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n721), .B1(new_n738), .B2(new_n739), .ZN(G1328gat));
  OAI21_X1  g539(.A(G36gat), .B1(new_n736), .B2(new_n689), .ZN(new_n741));
  AOI21_X1  g540(.A(G36gat), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n719), .A2(new_n690), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(G1329gat));
  NOR3_X1   g545(.A1(new_n735), .A2(new_n698), .A3(new_n718), .ZN(new_n747));
  INV_X1    g546(.A(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT105), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n700), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n719), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n747), .B2(new_n748), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n749), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  OAI221_X1 g553(.A(new_n751), .B1(KEYINPUT105), .B2(KEYINPUT47), .C1(new_n747), .C2(new_n748), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1330gat));
  INV_X1    g555(.A(KEYINPUT106), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n735), .A2(new_n499), .A3(new_n718), .ZN(new_n758));
  INV_X1    g557(.A(G50gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n719), .A2(new_n759), .A3(new_n286), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n762), .A3(KEYINPUT48), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT48), .ZN(new_n764));
  OAI221_X1 g563(.A(new_n761), .B1(new_n757), .B2(new_n764), .C1(new_n758), .C2(new_n759), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(G1331gat));
  AND2_X1   g565(.A1(new_n682), .A2(new_n683), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n639), .A2(new_n664), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n541), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n475), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n690), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT49), .B(G64gat), .Z(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n772), .B2(new_n774), .ZN(G1333gat));
  AND2_X1   g574(.A1(new_n769), .A2(new_n750), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n776), .A2(KEYINPUT107), .ZN(new_n777));
  INV_X1    g576(.A(G71gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(KEYINPUT107), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n769), .A2(G71gat), .A3(new_n697), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT50), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT50), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n780), .A2(new_n784), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(G1334gat));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n286), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  INV_X1    g587(.A(new_n638), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n665), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n716), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n664), .A2(new_n638), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT108), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n731), .A2(new_n793), .B1(new_n794), .B2(KEYINPUT51), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT109), .Z(new_n797));
  NAND3_X1  g596(.A1(new_n684), .A2(new_n566), .A3(new_n475), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n793), .A2(new_n684), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n735), .A2(new_n445), .A3(new_n799), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n797), .A2(new_n798), .B1(new_n566), .B2(new_n800), .ZN(G1336gat));
  NAND3_X1  g600(.A1(new_n690), .A2(new_n684), .A3(new_n567), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(KEYINPUT110), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT111), .B1(new_n796), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n735), .A2(new_n689), .A3(new_n799), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n567), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g606(.A(G99gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n750), .A2(new_n808), .A3(new_n684), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT112), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n735), .A2(new_n698), .A3(new_n799), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n797), .A2(new_n810), .B1(new_n808), .B2(new_n811), .ZN(G1338gat));
  NOR3_X1   g611(.A1(new_n767), .A2(new_n499), .A3(G106gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n792), .B2(new_n795), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(KEYINPUT113), .B2(new_n815), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n735), .A2(new_n499), .A3(new_n799), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(G106gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(KEYINPUT113), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n819), .ZN(new_n821));
  AOI211_X1 g620(.A(new_n821), .B(new_n816), .C1(new_n817), .C2(G106gat), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(G1339gat));
  AND2_X1   g622(.A1(new_n674), .A2(new_n675), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n681), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n675), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n670), .A2(new_n827), .A3(new_n672), .A4(new_n673), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n676), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n683), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n648), .A2(KEYINPUT115), .A3(new_n641), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n640), .A2(new_n643), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT115), .B1(new_n648), .B2(new_n641), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n655), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n826), .A2(new_n829), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n831), .A2(new_n658), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n724), .A2(new_n726), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n709), .A2(new_n723), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n725), .A2(KEYINPUT102), .A3(new_n706), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n684), .A2(new_n658), .A3(new_n836), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n831), .A2(new_n664), .A3(new_n839), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n842), .A2(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n789), .B1(new_n841), .B2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n600), .A2(new_n665), .A3(new_n638), .A4(new_n767), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n690), .A2(new_n445), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n411), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n291), .A3(new_n665), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n286), .B1(new_n495), .B2(new_n493), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n845), .A2(new_n844), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n856), .B1(new_n724), .B2(new_n726), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n683), .A3(new_n830), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n836), .A2(new_n658), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n843), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n638), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n848), .B(KEYINPUT114), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n475), .B(new_n855), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n690), .B1(new_n864), .B2(KEYINPUT116), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n866), .A3(new_n475), .A4(new_n855), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n664), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n854), .B1(new_n868), .B2(new_n291), .ZN(G1340gat));
  NOR3_X1   g668(.A1(new_n853), .A2(new_n293), .A3(new_n767), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n865), .A2(new_n684), .A3(new_n867), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n293), .ZN(G1341gat));
  XOR2_X1   g671(.A(KEYINPUT73), .B(G127gat), .Z(new_n873));
  NOR3_X1   g672(.A1(new_n853), .A2(new_n789), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n865), .A2(new_n638), .A3(new_n867), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n875), .B2(new_n873), .ZN(G1342gat));
  NOR2_X1   g675(.A1(new_n600), .A2(G134gat), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n865), .A2(new_n867), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n880), .A3(new_n867), .A4(new_n877), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n853), .B2(new_n600), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n879), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT117), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n879), .A2(new_n885), .A3(new_n881), .A4(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1343gat));
  AOI21_X1  g686(.A(new_n499), .B1(new_n847), .B2(new_n850), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n698), .A2(new_n852), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G141gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n664), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT118), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n837), .A2(new_n896), .A3(new_n838), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n895), .A2(new_n831), .A3(new_n664), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n709), .B1(new_n898), .B2(new_n844), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n861), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT119), .B(new_n709), .C1(new_n898), .C2(new_n844), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n789), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n850), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n894), .B1(new_n904), .B2(new_n286), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n851), .A2(new_n894), .A3(new_n286), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n890), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n907), .A3(new_n665), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n893), .B1(new_n908), .B2(new_n892), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT58), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n893), .B(new_n911), .C1(new_n908), .C2(new_n892), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n684), .ZN(new_n914));
  AOI21_X1  g713(.A(G148gat), .B1(new_n914), .B2(KEYINPUT59), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n905), .A2(new_n907), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n767), .A2(KEYINPUT59), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT57), .B(new_n286), .C1(new_n862), .C2(new_n863), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921));
  INV_X1    g720(.A(new_n848), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n860), .A2(new_n709), .ZN(new_n923));
  INV_X1    g722(.A(new_n844), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n896), .B1(new_n837), .B2(new_n838), .ZN(new_n925));
  AOI211_X1 g724(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n826), .C2(new_n829), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n830), .A2(new_n683), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n924), .B1(new_n928), .B2(new_n664), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n923), .B1(new_n929), .B2(new_n709), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n922), .B1(new_n930), .B2(new_n789), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n921), .B(new_n894), .C1(new_n931), .C2(new_n499), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n851), .A2(new_n933), .A3(KEYINPUT57), .A4(new_n286), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n840), .A2(new_n600), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n789), .B1(new_n899), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n499), .B1(new_n936), .B2(new_n848), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT121), .B1(new_n937), .B2(KEYINPUT57), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n920), .A2(new_n932), .A3(new_n934), .A4(new_n938), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(new_n684), .A3(new_n890), .ZN(new_n940));
  NAND2_X1  g739(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n918), .B1(new_n940), .B2(new_n941), .ZN(G1345gat));
  NAND3_X1  g741(.A1(new_n891), .A2(new_n215), .A3(new_n638), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n905), .A2(new_n907), .A3(new_n789), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n215), .ZN(G1346gat));
  AOI21_X1  g744(.A(G162gat), .B1(new_n891), .B2(new_n709), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n724), .A2(new_n726), .A3(new_n216), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n916), .B2(new_n947), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n689), .A2(new_n475), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n411), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n851), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n665), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n851), .A2(new_n855), .A3(new_n949), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT122), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n664), .A2(new_n316), .A3(new_n318), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(G1348gat));
  NAND3_X1  g758(.A1(new_n951), .A2(G176gat), .A3(new_n684), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT123), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n955), .A2(new_n684), .A3(new_n956), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n319), .ZN(G1349gat));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n638), .A2(new_n359), .ZN(new_n965));
  OR3_X1    g764(.A1(new_n954), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n954), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(G183gat), .B1(new_n952), .B2(new_n789), .ZN(new_n969));
  XNOR2_X1  g768(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(G1350gat));
  AOI21_X1  g772(.A(new_n306), .B1(new_n951), .B2(new_n709), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT61), .Z(new_n975));
  NAND2_X1  g774(.A1(new_n727), .A2(new_n306), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n957), .B2(new_n976), .ZN(G1351gat));
  NAND2_X1  g776(.A1(new_n698), .A2(new_n949), .ZN(new_n978));
  INV_X1    g777(.A(new_n978), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n888), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(G197gat), .B1(new_n980), .B2(new_n664), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n939), .A2(new_n979), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n665), .A2(new_n242), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(G1352gat));
  NAND3_X1  g783(.A1(new_n939), .A2(new_n684), .A3(new_n979), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(G204gat), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n888), .A2(new_n979), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n684), .A2(new_n247), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT62), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OR3_X1    g788(.A1(new_n987), .A2(KEYINPUT62), .A3(new_n988), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n939), .A2(new_n638), .A3(new_n979), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G211gat), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(KEYINPUT63), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT63), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n992), .A2(new_n995), .A3(G211gat), .ZN(new_n996));
  AND4_X1   g795(.A1(new_n240), .A2(new_n888), .A3(new_n638), .A4(new_n979), .ZN(new_n997));
  XOR2_X1   g796(.A(new_n997), .B(KEYINPUT126), .Z(new_n998));
  NAND3_X1  g797(.A1(new_n994), .A2(new_n996), .A3(new_n998), .ZN(G1354gat));
  AOI21_X1  g798(.A(G218gat), .B1(new_n980), .B2(new_n727), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n1000), .B(KEYINPUT127), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n982), .A2(G218gat), .A3(new_n709), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1355gat));
endmodule


