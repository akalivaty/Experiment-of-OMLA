//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g030(.A1(G113), .A2(G2104), .ZN(new_n456));
  XNOR2_X1  g031(.A(KEYINPUT3), .B(G2104), .ZN(new_n457));
  AOI21_X1  g032(.A(KEYINPUT65), .B1(new_n457), .B2(G125), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  AND4_X1   g037(.A1(KEYINPUT65), .A2(new_n460), .A3(new_n462), .A4(G125), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n456), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n459), .A2(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(new_n461), .A3(G2104), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(new_n460), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n470), .A2(KEYINPUT67), .A3(new_n471), .A4(new_n473), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n471), .A2(new_n469), .A3(new_n460), .A4(new_n473), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n467), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g053(.A1(new_n465), .A2(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n471), .A2(new_n469), .A3(G2105), .A4(new_n460), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT68), .ZN(new_n486));
  INV_X1    g061(.A(G2105), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n470), .A2(new_n487), .A3(new_n471), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g064(.A(new_n482), .B(new_n486), .C1(G136), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n490), .B(KEYINPUT69), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n471), .A2(new_n469), .A3(new_n460), .A4(new_n494), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n495), .A2(KEYINPUT4), .B1(new_n457), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(G114), .B2(new_n487), .ZN(new_n500));
  INV_X1    g075(.A(G126), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n480), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(G164));
  OR2_X1    g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n509), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT6), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(new_n508), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n525), .C1(new_n526), .C2(new_n511), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n504), .A2(new_n528), .A3(new_n505), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT70), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n532), .A3(G651), .ZN(new_n533));
  INV_X1    g108(.A(G63), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n527), .A2(new_n535), .ZN(G168));
  NAND3_X1  g111(.A1(new_n529), .A2(new_n532), .A3(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n508), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  INV_X1    g115(.A(G52), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n511), .A2(new_n540), .B1(new_n513), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  NAND3_X1  g118(.A1(new_n529), .A2(new_n532), .A3(G56), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n508), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n511), .A2(new_n547), .B1(new_n513), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  AOI22_X1  g130(.A1(new_n504), .A2(new_n505), .B1(new_n520), .B2(new_n521), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n504), .A2(new_n561), .A3(new_n505), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT73), .B1(new_n530), .B2(new_n531), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n560), .B1(new_n564), .B2(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n557), .B1(new_n565), .B2(new_n508), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n522), .A2(KEYINPUT71), .A3(G53), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  OR2_X1    g146(.A1(new_n539), .A2(new_n542), .ZN(G301));
  INV_X1    g147(.A(G168), .ZN(G286));
  AOI22_X1  g148(.A1(new_n556), .A2(G87), .B1(new_n522), .B2(G49), .ZN(new_n574));
  NAND2_X1  g149(.A1(G74), .A2(G651), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n533), .A2(KEYINPUT74), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT74), .B1(new_n533), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(G288));
  OAI21_X1  g153(.A(G61), .B1(new_n530), .B2(new_n531), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n556), .B2(G86), .ZN(new_n582));
  AND2_X1   g157(.A1(KEYINPUT6), .A2(G651), .ZN(new_n583));
  NOR2_X1   g158(.A1(KEYINPUT6), .A2(G651), .ZN(new_n584));
  OAI211_X1 g159(.A(G48), .B(G543), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT75), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n510), .A2(new_n587), .A3(G48), .A4(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n582), .A2(new_n589), .ZN(G305));
  NAND3_X1  g165(.A1(new_n529), .A2(new_n532), .A3(G60), .ZN(new_n591));
  INV_X1    g166(.A(G72), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n592), .B2(new_n518), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n508), .B1(new_n593), .B2(KEYINPUT76), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(KEYINPUT76), .B2(new_n593), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n556), .A2(G85), .B1(new_n522), .B2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n556), .A2(G92), .ZN(new_n599));
  XOR2_X1   g174(.A(new_n599), .B(KEYINPUT10), .Z(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT77), .B(G66), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n564), .A2(new_n601), .B1(G79), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n602), .A2(new_n508), .B1(new_n603), .B2(new_n513), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT78), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI221_X1 g181(.A(KEYINPUT78), .B1(new_n603), .B2(new_n513), .C1(new_n602), .C2(new_n508), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n598), .B1(new_n608), .B2(G868), .ZN(G284));
  OAI21_X1  g184(.A(new_n598), .B1(new_n608), .B2(G868), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n570), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n570), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n608), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n608), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  INV_X1    g195(.A(G111), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n620), .A2(KEYINPUT80), .B1(new_n621), .B2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(KEYINPUT80), .B2(new_n620), .ZN(new_n623));
  INV_X1    g198(.A(G123), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI221_X1 g200(.A(new_n623), .B1(new_n624), .B2(new_n480), .C1(new_n488), .C2(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n457), .A2(new_n466), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n626), .A2(G2096), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n627), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT81), .ZN(G156));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n639), .B2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT82), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n655), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n652), .B(new_n656), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n652), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n654), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n655), .A2(new_n652), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n658), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n660), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2100), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT83), .B(G2096), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n676), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n677), .A2(KEYINPUT20), .A3(new_n676), .ZN(new_n682));
  OAI221_X1 g257(.A(new_n678), .B1(new_n676), .B2(new_n674), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1981), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  NOR2_X1   g267(.A1(G16), .A2(G23), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT87), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(G288), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n696), .B(new_n697), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(G22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT88), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G303), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1971), .ZN(new_n702));
  MUX2_X1   g277(.A(G6), .B(G305), .S(G16), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT32), .B(G1981), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n698), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT34), .ZN(new_n707));
  INV_X1    g282(.A(G119), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n480), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT85), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n489), .A2(G131), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n487), .A2(G107), .ZN(new_n712));
  OAI21_X1  g287(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n710), .B(new_n711), .C1(new_n712), .C2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G25), .B(new_n714), .S(G29), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G290), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G24), .ZN(new_n719));
  OR3_X1    g294(.A1(new_n719), .A2(KEYINPUT86), .A3(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT86), .B1(new_n719), .B2(G16), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G1986), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n707), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n726), .A2(KEYINPUT89), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G35), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G162), .B2(new_n729), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n608), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G4), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1348), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n695), .A2(G19), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n550), .B2(new_n695), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1341), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT24), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n743), .B2(new_n744), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G160), .B2(new_n729), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n742), .B1(G2084), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n737), .A2(new_n738), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n747), .A2(G2084), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n739), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n695), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n695), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1966), .ZN(new_n755));
  NOR2_X1   g330(.A1(G164), .A2(new_n729), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G27), .B2(new_n729), .ZN(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n755), .B1(G2078), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n695), .A2(G5), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G171), .B2(new_n695), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(G1961), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(G1961), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n626), .A2(new_n729), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT30), .B(G28), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n765), .A2(new_n729), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n763), .B1(new_n770), .B2(KEYINPUT95), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n772));
  INV_X1    g347(.A(G2078), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n769), .A2(new_n772), .B1(new_n757), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n759), .A2(new_n762), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n729), .A2(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n487), .A2(G103), .A3(G2104), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  AOI22_X1  g353(.A1(new_n457), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  INV_X1    g354(.A(G139), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n778), .B1(new_n779), .B2(new_n487), .C1(new_n488), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT93), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n782), .B2(new_n729), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2072), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n729), .A2(G32), .ZN(new_n785));
  NAND3_X1  g360(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT26), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(G105), .B2(new_n466), .ZN(new_n790));
  INV_X1    g365(.A(G129), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n480), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n489), .B2(G141), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n785), .B1(new_n793), .B2(new_n729), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT94), .Z(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT27), .B(G1996), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n775), .A2(new_n784), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n695), .A2(G20), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT23), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n570), .B2(new_n695), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1956), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n796), .B2(new_n795), .ZN(new_n803));
  INV_X1    g378(.A(G104), .ZN(new_n804));
  AND3_X1   g379(.A1(new_n804), .A2(new_n487), .A3(KEYINPUT90), .ZN(new_n805));
  AOI21_X1  g380(.A(KEYINPUT90), .B1(new_n804), .B2(new_n487), .ZN(new_n806));
  OAI221_X1 g381(.A(G2104), .B1(G116), .B2(new_n487), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(G128), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(new_n480), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G140), .B2(new_n489), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n729), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT91), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n729), .A2(G26), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT28), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT92), .B(G2067), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  AND3_X1   g392(.A1(new_n798), .A2(new_n803), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n728), .A2(new_n735), .A3(new_n752), .A4(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  NAND3_X1  g395(.A1(new_n529), .A2(new_n532), .A3(G67), .ZN(new_n821));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n508), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n511), .A2(new_n824), .B1(new_n513), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n829));
  INV_X1    g404(.A(new_n550), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT97), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n550), .A2(new_n827), .A3(new_n831), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n608), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n828), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n782), .B(new_n793), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n714), .B(new_n629), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n457), .A2(new_n496), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n497), .A2(KEYINPUT98), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n502), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n810), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n489), .A2(G142), .ZN(new_n858));
  INV_X1    g433(.A(G130), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n487), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n858), .B1(new_n859), .B2(new_n480), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n857), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n849), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(G160), .B(new_n626), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n491), .B(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n847), .A2(new_n848), .A3(new_n863), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G37), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n865), .A2(new_n868), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n872), .B(KEYINPUT40), .C1(new_n867), .C2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n867), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n876), .B2(new_n871), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n874), .A2(new_n877), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n616), .B(new_n835), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n606), .A2(new_n607), .ZN(new_n881));
  INV_X1    g456(.A(new_n600), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n570), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n608), .A2(G299), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n879), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n888), .B1(new_n608), .B2(G299), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n883), .A2(KEYINPUT99), .A3(new_n570), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n608), .B2(G299), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n891), .A2(new_n892), .B1(new_n893), .B2(new_n884), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n887), .B1(new_n894), .B2(new_n880), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT101), .ZN(new_n896));
  NAND2_X1  g471(.A1(G290), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n595), .A2(KEYINPUT101), .A3(new_n596), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(G288), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(G288), .A3(new_n898), .ZN(new_n902));
  XNOR2_X1  g477(.A(G303), .B(G305), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT42), .ZN(new_n908));
  OR3_X1    g483(.A1(new_n894), .A2(KEYINPUT100), .A3(new_n880), .ZN(new_n909));
  OR3_X1    g484(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT42), .ZN(new_n910));
  AND4_X1   g485(.A1(new_n895), .A2(new_n908), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n908), .A2(new_n910), .B1(new_n909), .B2(new_n895), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g489(.A(new_n913), .B1(G868), .B2(new_n827), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n916));
  NAND2_X1  g491(.A1(G301), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G171), .A2(KEYINPUT102), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(G168), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(G286), .A2(G301), .A3(new_n916), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g496(.A1(new_n835), .A2(new_n921), .A3(KEYINPUT104), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n835), .A2(new_n921), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n833), .A2(new_n919), .A3(new_n834), .A4(new_n920), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(KEYINPUT104), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n889), .A2(new_n893), .A3(new_n890), .ZN(new_n927));
  INV_X1    g502(.A(new_n886), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n927), .B1(new_n928), .B2(KEYINPUT41), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n923), .A2(new_n930), .A3(new_n924), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n835), .A2(KEYINPUT103), .A3(new_n921), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n926), .A2(new_n929), .B1(new_n886), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n870), .B1(new_n934), .B2(new_n907), .ZN(new_n935));
  OAI22_X1  g510(.A1(new_n926), .A2(new_n928), .B1(new_n894), .B2(new_n933), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(new_n906), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n936), .B2(new_n906), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n894), .A2(new_n933), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n941), .B(new_n907), .C1(new_n928), .C2(new_n926), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT43), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT44), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n935), .A2(new_n937), .A3(KEYINPUT43), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n938), .B1(new_n940), .B2(new_n942), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(G397));
  INV_X1    g524(.A(new_n502), .ZN(new_n950));
  AOI221_X4 g525(.A(new_n853), .B1(new_n457), .B2(new_n496), .C1(new_n495), .C2(KEYINPUT4), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT98), .B1(new_n850), .B2(new_n851), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT45), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n465), .A2(new_n478), .A3(G40), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n810), .B(G2067), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n793), .B(G1996), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT105), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n714), .B(new_n716), .Z(new_n962));
  OAI21_X1  g537(.A(new_n961), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n957), .ZN(new_n964));
  XNOR2_X1  g539(.A(G290), .B(G1986), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G2067), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n854), .A2(new_n855), .ZN(new_n968));
  AOI21_X1  g543(.A(G1384), .B1(new_n968), .B2(new_n950), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT116), .B1(new_n969), .B2(new_n956), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n953), .A2(new_n954), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n465), .A2(new_n478), .A3(G40), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n967), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n953), .A2(new_n976), .A3(new_n954), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n954), .B1(new_n497), .B2(new_n502), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT50), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n956), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n738), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT60), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT120), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n608), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n975), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n608), .A2(new_n983), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n986), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n975), .A2(new_n988), .A3(new_n981), .A4(new_n984), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n975), .A2(new_n981), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n982), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT110), .B(G1956), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT50), .B1(new_n856), .B2(G1384), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n976), .B(new_n954), .C1(new_n497), .C2(new_n502), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n973), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n993), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n999), .A2(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n953), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n978), .A2(new_n999), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT114), .B(KEYINPUT56), .Z(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(G2072), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1001), .A2(new_n956), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n973), .B1(new_n999), .B2(new_n978), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1008), .A2(KEYINPUT115), .A3(new_n1001), .A4(new_n1004), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n998), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n565), .A2(new_n508), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n567), .B(KEYINPUT9), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(KEYINPUT57), .A3(new_n1012), .A4(new_n557), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT113), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n566), .A2(KEYINPUT111), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(new_n557), .C1(new_n565), .C2(new_n508), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1015), .A2(new_n1012), .A3(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n1018), .A2(KEYINPUT112), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT112), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1014), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT61), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1010), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1010), .B2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1010), .A2(new_n1022), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT59), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT118), .ZN(new_n1029));
  XOR2_X1   g604(.A(new_n1029), .B(KEYINPUT119), .Z(new_n1030));
  OAI21_X1  g605(.A(new_n972), .B1(new_n971), .B2(new_n973), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n956), .A2(KEYINPUT116), .A3(new_n954), .A4(new_n953), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT58), .B(G1341), .Z(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1996), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1008), .A2(new_n1035), .A3(new_n1001), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n550), .B1(KEYINPUT118), .B2(new_n1028), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1030), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1030), .ZN(new_n1041));
  AOI211_X1 g616(.A(new_n1041), .B(new_n1038), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n992), .A2(new_n1024), .A3(new_n1027), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1010), .B1(new_n1045), .B2(new_n1022), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1022), .A2(new_n1045), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n883), .B1(new_n975), .B2(new_n981), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1046), .A2(new_n1047), .B1(new_n1026), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g625(.A(KEYINPUT123), .B(G1961), .Z(new_n1051));
  OAI21_X1  g626(.A(new_n1000), .B1(new_n497), .B2(new_n502), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1052), .A2(new_n465), .A3(G40), .A4(new_n478), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n971), .B2(new_n999), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(G2078), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n980), .A2(new_n1051), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1001), .A2(new_n773), .A3(new_n956), .A4(new_n1002), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1058), .A2(KEYINPUT124), .A3(new_n1055), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT124), .B1(new_n1058), .B2(new_n1055), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1057), .B(G301), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n953), .A2(new_n976), .A3(new_n954), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n956), .A2(new_n979), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1051), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n971), .A2(new_n999), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n478), .A2(G40), .A3(new_n1056), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT126), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n464), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n487), .B1(new_n464), .B2(new_n1067), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1066), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1001), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1058), .A2(new_n1055), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1058), .A2(KEYINPUT124), .A3(new_n1055), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1061), .B(KEYINPUT54), .C1(new_n1077), .C2(G301), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n955), .B2(new_n1053), .ZN(new_n1081));
  INV_X1    g656(.A(G2084), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n977), .A2(new_n1082), .A3(new_n956), .A4(new_n979), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G8), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT121), .B1(new_n1085), .B2(G168), .ZN(new_n1086));
  INV_X1    g661(.A(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1087), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(G286), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G168), .A2(new_n1087), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT51), .B1(new_n1092), .B2(KEYINPUT122), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1085), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1093), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1086), .A2(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(G1976), .B(new_n574), .C1(new_n576), .C2(new_n577), .ZN(new_n1098));
  OAI211_X1 g673(.A(G8), .B(new_n1098), .C1(new_n971), .C2(new_n973), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT52), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT108), .ZN(new_n1101));
  INV_X1    g676(.A(G1981), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n556), .A2(G86), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n581), .A2(G651), .ZN(new_n1104));
  AND4_X1   g679(.A1(new_n1102), .A2(new_n589), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1102), .B1(new_n582), .B2(new_n589), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1101), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT49), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n956), .A2(new_n954), .A3(new_n953), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT49), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1101), .B(new_n1110), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1108), .A2(new_n1109), .A3(G8), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1100), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(G1976), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT52), .B1(G288), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1109), .A2(G8), .A3(new_n1098), .A4(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT107), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1087), .B1(new_n969), .B2(new_n956), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT107), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1098), .A4(new_n1115), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1113), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1971), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n956), .A2(new_n1002), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1000), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n968), .B2(new_n950), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1122), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n994), .A2(new_n732), .A3(new_n997), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1087), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G303), .A2(G8), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT55), .Z(new_n1130));
  OR2_X1    g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n977), .A2(new_n732), .A3(new_n956), .A4(new_n979), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1087), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1133), .A2(KEYINPUT106), .A3(new_n1130), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT106), .B1(new_n1133), .B2(new_n1130), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1121), .B(new_n1131), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1079), .A2(new_n1097), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(G171), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT125), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1141), .A3(G171), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1077), .A2(G301), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1050), .A2(new_n1137), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT63), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1088), .A2(G168), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1136), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1133), .A2(new_n1130), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1151), .A2(new_n1149), .A3(new_n1148), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1152), .B(new_n1121), .C1(new_n1135), .C2(new_n1134), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1150), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1093), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1088), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1156));
  AND4_X1   g731(.A1(new_n1089), .A2(new_n1084), .A3(G8), .A4(G286), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1089), .B1(new_n1088), .B2(G286), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1155), .A2(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT62), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1113), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1163), .B(new_n1164), .C1(new_n1130), .C2(new_n1128), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1160), .A2(new_n1161), .A3(new_n1166), .A4(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1112), .A2(new_n1114), .A3(new_n900), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(G1981), .B2(G305), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1118), .B(KEYINPUT109), .Z(new_n1174));
  AOI22_X1  g749(.A1(new_n1162), .A2(new_n1121), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1154), .A2(new_n1171), .A3(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n966), .B1(new_n1147), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n957), .B1(new_n958), .B2(new_n793), .ZN(new_n1178));
  OR3_X1    g753(.A1(new_n957), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT46), .B1(new_n957), .B2(G1996), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT47), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n714), .A2(new_n716), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n961), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n810), .A2(new_n967), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n957), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n957), .A2(G1986), .A3(G290), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT127), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1188), .A2(KEYINPUT48), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n963), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1188), .A2(KEYINPUT48), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1182), .B(new_n1186), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1177), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g768(.A1(new_n946), .A2(new_n947), .ZN(new_n1195));
  OAI21_X1  g769(.A(G319), .B1(new_n649), .B2(new_n650), .ZN(new_n1196));
  OR2_X1    g770(.A1(G227), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n690), .B2(new_n691), .ZN(new_n1198));
  OAI21_X1  g772(.A(new_n1198), .B1(new_n876), .B2(new_n871), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1195), .A2(new_n1199), .ZN(G308));
  OAI221_X1 g774(.A(new_n1198), .B1(new_n876), .B2(new_n871), .C1(new_n946), .C2(new_n947), .ZN(G225));
endmodule


