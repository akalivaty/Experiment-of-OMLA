//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1205, new_n1206, new_n1207;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT65), .B(G452), .ZN(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G101), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n467), .A2(new_n473), .ZN(G160));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n472), .B2(G112), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT69), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n469), .B2(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n475), .A2(KEYINPUT68), .A3(new_n472), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  OAI221_X1 g061(.A(new_n478), .B1(new_n479), .B2(new_n481), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NOR2_X1   g063(.A1(new_n462), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G102), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(new_n462), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n475), .B2(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n490), .B1(new_n493), .B2(new_n472), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n472), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n475), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n494), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(new_n506), .A3(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n502), .A2(new_n504), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT70), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(G50), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n512), .A2(G651), .B1(new_n513), .B2(new_n516), .ZN(G166));
  NAND3_X1  g092(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n519), .A2(G543), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n513), .A2(new_n502), .A3(new_n504), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n528), .A2(new_n529), .B1(G89), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  NAND2_X1  g111(.A1(new_n531), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n509), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n537), .B(new_n541), .C1(new_n542), .C2(new_n524), .ZN(G301));
  INV_X1    g118(.A(G301), .ZN(G171));
  AND3_X1   g119(.A1(new_n519), .A2(G543), .A3(new_n523), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n509), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n531), .A2(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND3_X1  g134(.A1(new_n545), .A2(KEYINPUT9), .A3(G53), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT73), .B(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n509), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n531), .A2(G91), .B1(new_n563), .B2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n524), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n560), .A2(new_n564), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND4_X1  g144(.A1(new_n519), .A2(G49), .A3(G543), .A4(new_n523), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n505), .A2(G87), .A3(new_n513), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  NAND3_X1  g148(.A1(new_n505), .A2(G86), .A3(new_n513), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n505), .A2(KEYINPUT74), .A3(G86), .A4(new_n513), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n513), .A2(G48), .A3(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  INV_X1    g156(.A(G73), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n509), .A2(new_n581), .B1(new_n582), .B2(new_n501), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n580), .B1(G651), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n578), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n545), .A2(G47), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT75), .B(G85), .Z(new_n587));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n509), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n531), .A2(new_n587), .B1(new_n590), .B2(G651), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n586), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n530), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n509), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n598), .B(new_n602), .C1(new_n603), .C2(new_n524), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT76), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n593), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n552), .A2(new_n608), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n605), .A2(new_n612), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT77), .Z(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g193(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT79), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n475), .A2(new_n489), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n620), .B(new_n621), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n477), .A2(G123), .ZN(new_n625));
  NOR2_X1   g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(new_n472), .B2(G111), .ZN(new_n627));
  INV_X1    g202(.A(G135), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n625), .B1(new_n626), .B2(new_n627), .C1(new_n485), .C2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT80), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n624), .A2(new_n631), .ZN(G156));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  OAI21_X1  g210(.A(KEYINPUT14), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT81), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n639), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(G14), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2067), .B(G2678), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n650), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n652), .B2(new_n653), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n655), .B1(new_n654), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n658), .B(new_n661), .Z(G227));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n674), .C1(new_n672), .C2(new_n671), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G1981), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G22), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G166), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G1971), .ZN(new_n687));
  INV_X1    g262(.A(G1971), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n688), .B(new_n685), .C1(G166), .C2(new_n684), .ZN(new_n689));
  NAND4_X1  g264(.A1(new_n570), .A2(G16), .A3(new_n571), .A4(new_n572), .ZN(new_n690));
  OR2_X1    g265(.A1(G16), .A2(G23), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT33), .B(G1976), .Z(new_n692));
  AND3_X1   g267(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n690), .B2(new_n691), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n687), .A2(new_n689), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(G305), .A2(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n684), .A2(G6), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n699), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n684), .B1(new_n578), .B2(new_n584), .ZN(new_n702));
  INV_X1    g277(.A(new_n698), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n683), .B1(new_n696), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n696), .A2(new_n705), .A3(new_n683), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(KEYINPUT34), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n707), .B2(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n684), .A2(G24), .ZN(new_n713));
  INV_X1    g288(.A(G290), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n684), .ZN(new_n715));
  INV_X1    g290(.A(G1986), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G131), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n485), .A2(KEYINPUT85), .A3(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(G95), .A2(G2105), .ZN(new_n720));
  INV_X1    g295(.A(G107), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n462), .B1(new_n721), .B2(G2105), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n477), .A2(G119), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(KEYINPUT85), .B1(new_n485), .B2(new_n718), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT84), .B(G29), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n726), .A2(G25), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n717), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(KEYINPUT87), .B1(new_n712), .B2(new_n734), .ZN(new_n735));
  AND3_X1   g310(.A1(new_n687), .A2(new_n689), .A3(new_n695), .ZN(new_n736));
  INV_X1    g311(.A(new_n705), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT86), .ZN(new_n738));
  AOI21_X1  g313(.A(KEYINPUT34), .B1(new_n738), .B2(new_n706), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT87), .ZN(new_n740));
  NOR3_X1   g315(.A1(new_n739), .A2(new_n740), .A3(new_n733), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n710), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(KEYINPUT88), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n712), .A2(KEYINPUT87), .A3(new_n734), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n740), .B1(new_n739), .B2(new_n733), .ZN(new_n745));
  AOI22_X1  g320(.A1(new_n744), .A2(new_n745), .B1(new_n709), .B2(KEYINPUT34), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n743), .A2(new_n748), .A3(KEYINPUT36), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n750));
  AOI21_X1  g325(.A(KEYINPUT89), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n743), .A2(new_n748), .A3(KEYINPUT89), .A4(KEYINPUT36), .ZN(new_n753));
  NAND2_X1  g328(.A1(G160), .A2(G29), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT24), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n726), .B1(new_n755), .B2(G34), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n755), .A2(G34), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n756), .A2(new_n757), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT98), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n726), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n726), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT29), .ZN(new_n768));
  INV_X1    g343(.A(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(KEYINPUT29), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n684), .A2(G19), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n553), .B2(new_n684), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT92), .B(G1341), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n765), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(G29), .A2(G32), .ZN(new_n777));
  INV_X1    g352(.A(new_n485), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G141), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n489), .A2(G105), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n477), .A2(G129), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n782));
  NAND3_X1  g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n779), .A2(new_n780), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n777), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n762), .A2(new_n763), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT30), .B(G28), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n790), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT31), .B(G11), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n789), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(G299), .A2(G16), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n684), .A2(KEYINPUT23), .A3(G20), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT23), .ZN(new_n797));
  INV_X1    g372(.A(G20), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G16), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n795), .A2(new_n796), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1956), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n776), .A2(new_n794), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n726), .A2(G27), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n726), .ZN(new_n804));
  INV_X1    g379(.A(G2078), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n684), .A2(G21), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G168), .B2(new_n684), .ZN(new_n808));
  INV_X1    g383(.A(G1966), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n812));
  NAND2_X1  g387(.A1(G171), .A2(G16), .ZN(new_n813));
  OR2_X1    g388(.A1(G5), .A2(G16), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n812), .B1(new_n816), .B2(G1961), .ZN(new_n817));
  INV_X1    g392(.A(G1961), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n815), .A2(KEYINPUT97), .A3(new_n818), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n811), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n802), .A2(new_n806), .A3(new_n810), .A4(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n629), .A2(new_n726), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n489), .A2(G103), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT25), .Z(new_n824));
  AOI22_X1  g399(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n825));
  INV_X1    g400(.A(G139), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n824), .B1(new_n472), .B2(new_n825), .C1(new_n485), .C2(new_n826), .ZN(new_n827));
  MUX2_X1   g402(.A(G33), .B(new_n827), .S(G29), .Z(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(G2072), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(G2072), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n829), .B(new_n830), .C1(G1961), .C2(new_n816), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n821), .A2(new_n822), .A3(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n605), .A2(G16), .ZN(new_n833));
  NOR2_X1   g408(.A1(G4), .A2(G16), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT90), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(KEYINPUT90), .B2(new_n834), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT91), .B(G1348), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n836), .B(new_n837), .Z(new_n838));
  NAND2_X1  g413(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n726), .A2(KEYINPUT28), .A3(G26), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n778), .A2(G140), .ZN(new_n842));
  OR2_X1    g417(.A1(G104), .A2(G2105), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n843), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n844));
  INV_X1    g419(.A(G128), .ZN(new_n845));
  OAI21_X1  g420(.A(KEYINPUT93), .B1(new_n476), .B2(new_n845), .ZN(new_n846));
  OR3_X1    g421(.A1(new_n476), .A2(KEYINPUT93), .A3(new_n845), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n842), .A2(new_n844), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n841), .B1(new_n849), .B2(new_n786), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT28), .B1(new_n726), .B2(G26), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT94), .B(G2067), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n752), .A2(new_n753), .A3(new_n840), .A4(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(G311));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n839), .B1(new_n749), .B2(new_n751), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n859), .A2(KEYINPUT99), .A3(new_n753), .A4(new_n854), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(G150));
  NAND2_X1  g436(.A1(new_n605), .A2(G559), .ZN(new_n862));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n509), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G651), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT101), .B(G55), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n545), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n531), .A2(G93), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(new_n874), .A3(new_n552), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n552), .A2(new_n874), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n867), .A2(new_n868), .B1(G93), .B2(new_n531), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n546), .A2(KEYINPUT102), .A3(new_n550), .A4(new_n551), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n871), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n862), .B(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n883), .A2(KEYINPUT104), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(G860), .B1(new_n883), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT104), .B1(new_n883), .B2(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n873), .A2(G860), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT37), .Z(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(G145));
  XNOR2_X1  g466(.A(new_n629), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  INV_X1    g468(.A(G126), .ZN(new_n894));
  OAI22_X1  g469(.A1(new_n469), .A2(new_n894), .B1(new_n491), .B2(new_n462), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n895), .A2(G2105), .B1(G102), .B2(new_n489), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n497), .A2(new_n498), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n497), .B2(new_n498), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n848), .B(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(new_n827), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n827), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n785), .ZN(new_n905));
  INV_X1    g480(.A(new_n785), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n778), .A2(G142), .B1(G130), .B2(new_n477), .ZN(new_n909));
  NOR2_X1   g484(.A1(G106), .A2(G2105), .ZN(new_n910));
  OAI21_X1  g485(.A(G2104), .B1(new_n472), .B2(G118), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(new_n725), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n622), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n905), .A2(new_n914), .A3(new_n907), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n893), .B1(new_n918), .B2(KEYINPUT106), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G37), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n893), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g500(.A1(new_n873), .A2(new_n608), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n616), .B(new_n880), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n602), .B1(new_n524), .B2(new_n603), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n597), .B2(new_n594), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n929), .A2(G299), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(G299), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT41), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n930), .A2(new_n931), .A3(KEYINPUT107), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n929), .A2(G299), .A3(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n934), .B1(new_n937), .B2(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n927), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n927), .B2(new_n933), .ZN(new_n940));
  XNOR2_X1  g515(.A(G290), .B(G288), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  OR2_X1    g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  XNOR2_X1  g519(.A(G305), .B(G166), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n945), .A2(new_n941), .A3(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n946), .A2(KEYINPUT109), .A3(new_n947), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT109), .B1(new_n946), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n953), .B2(KEYINPUT42), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n940), .B(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n926), .B1(new_n955), .B2(new_n608), .ZN(G295));
  OAI21_X1  g531(.A(new_n926), .B1(new_n955), .B2(new_n608), .ZN(G331));
  NAND2_X1  g532(.A1(G301), .A2(KEYINPUT110), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT111), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n880), .ZN(new_n961));
  NOR2_X1   g536(.A1(G301), .A2(KEYINPUT110), .ZN(new_n962));
  NOR2_X1   g537(.A1(G286), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n875), .A3(new_n879), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n961), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n932), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n963), .ZN(new_n969));
  INV_X1    g544(.A(new_n964), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n959), .B1(new_n875), .B2(new_n879), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n938), .A3(new_n965), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n952), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G37), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n952), .B1(new_n968), .B2(new_n973), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n976), .A2(KEYINPUT43), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n937), .A2(KEYINPUT41), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT41), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n932), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(KEYINPUT112), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n937), .A2(new_n983), .A3(KEYINPUT41), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n982), .A2(new_n972), .A3(new_n965), .A4(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n985), .A2(KEYINPUT113), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n968), .B1(new_n985), .B2(KEYINPUT113), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n953), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n974), .A2(new_n975), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n978), .B(KEYINPUT44), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n991), .A3(new_n989), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT43), .B1(new_n976), .B2(new_n977), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  AOI211_X1 g573(.A(KEYINPUT114), .B(KEYINPUT44), .C1(new_n994), .C2(new_n995), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(G397));
  NAND2_X1  g575(.A1(new_n499), .A2(KEYINPUT105), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n497), .A2(new_n498), .A3(new_n897), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(G1384), .B1(new_n1003), .B2(new_n896), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(KEYINPUT45), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n467), .A2(new_n473), .A3(G40), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(G1996), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT116), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n848), .A2(G2067), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(G1996), .B2(new_n785), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n848), .A2(G2067), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g590(.A1(new_n1011), .A2(new_n785), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1016), .A2(new_n729), .A3(new_n725), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1009), .B1(new_n1017), .B2(new_n1012), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n725), .B(new_n729), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1016), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G290), .A2(G1986), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT115), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(new_n1008), .ZN(new_n1023));
  XOR2_X1   g598(.A(new_n1023), .B(KEYINPUT48), .Z(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1011), .B(KEYINPUT46), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1012), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n906), .A3(new_n1014), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1026), .B1(new_n1008), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1030), .A2(KEYINPUT47), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(KEYINPUT47), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1018), .B(new_n1025), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1384), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n900), .A2(KEYINPUT45), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n494), .B2(new_n499), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1006), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT56), .B(G2072), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1041), .A2(KEYINPUT124), .ZN(new_n1042));
  INV_X1    g617(.A(G1956), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1004), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1007), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g622(.A(G299), .B(KEYINPUT57), .Z(new_n1048));
  NAND2_X1  g623(.A1(new_n1041), .A2(KEYINPUT124), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1042), .A2(new_n1047), .A3(new_n1048), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT61), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n900), .A2(new_n1007), .A3(new_n1035), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT58), .B(G1341), .Z(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1055), .B1(new_n1056), .B2(G1996), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n553), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT59), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n900), .A2(new_n1044), .A3(new_n1035), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1037), .A2(KEYINPUT50), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1007), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n837), .ZN(new_n1063));
  INV_X1    g638(.A(G2067), .ZN(new_n1064));
  AND4_X1   g639(.A1(new_n1035), .A2(new_n900), .A3(new_n1064), .A4(new_n1007), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT60), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1067), .A2(KEYINPUT125), .A3(new_n1068), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1068), .B(new_n1065), .C1(new_n837), .C2(new_n1062), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n929), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI211_X1 g647(.A(KEYINPUT125), .B(new_n604), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT60), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1052), .B(new_n1059), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1050), .A2(new_n929), .A3(new_n1067), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1042), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1048), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(new_n1077), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1056), .A2(G2078), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(KEYINPUT53), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n818), .B2(new_n1062), .ZN(new_n1084));
  XNOR2_X1  g659(.A(G301), .B(KEYINPUT54), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1036), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n900), .A2(new_n1035), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1006), .B1(new_n1088), .B2(new_n1038), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(KEYINPUT53), .A3(new_n805), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1084), .B(new_n1086), .C1(new_n1087), .C2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT119), .B(G8), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1093), .B1(new_n532), .B2(new_n534), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1966), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1060), .A2(new_n763), .A3(new_n1007), .A4(new_n1061), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G8), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1095), .B(new_n1007), .C1(new_n1004), .C2(KEYINPUT45), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n809), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1102), .B2(new_n1097), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT51), .B(new_n1099), .C1(new_n1103), .C2(new_n1094), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1094), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1105), .B(new_n1106), .C1(new_n1107), .C2(new_n1093), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1091), .A2(new_n1104), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1095), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1084), .B1(new_n1110), .B2(new_n1090), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1085), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G1976), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1053), .B(new_n1092), .C1(new_n1113), .C2(G288), .ZN(new_n1114));
  AND2_X1   g689(.A1(G288), .A2(new_n1113), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1114), .A2(KEYINPUT52), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1114), .A2(KEYINPUT52), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT120), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1114), .A2(new_n1119), .A3(KEYINPUT52), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1116), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n582), .A2(new_n501), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n505), .B2(G61), .ZN(new_n1123));
  INV_X1    g698(.A(G651), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n579), .B(new_n574), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G1981), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT121), .ZN(new_n1127));
  INV_X1    g702(.A(G1981), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n578), .A2(new_n584), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(new_n1130), .A3(G1981), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT49), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1127), .A2(KEYINPUT49), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1093), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT122), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1134), .A2(new_n1139), .A3(new_n1136), .A4(new_n1135), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1121), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(G303), .A2(G8), .ZN(new_n1143));
  XOR2_X1   g718(.A(new_n1143), .B(KEYINPUT55), .Z(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1046), .B1(KEYINPUT50), .B2(new_n1088), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  AOI21_X1  g722(.A(G2090), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT123), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1149));
  AOI22_X1  g724(.A1(new_n1148), .A2(new_n1149), .B1(new_n688), .B2(new_n1056), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1145), .B1(new_n1150), .B2(new_n1093), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1152), .B1(new_n1056), .B2(new_n688), .ZN(new_n1153));
  AOI211_X1 g728(.A(KEYINPUT117), .B(G1971), .C1(new_n1036), .C2(new_n1039), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1060), .A2(new_n769), .A3(new_n1007), .A4(new_n1061), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1100), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT118), .B1(new_n1157), .B2(new_n1144), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1056), .A2(new_n688), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT117), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1056), .A2(new_n1152), .A3(new_n688), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n1156), .A3(new_n1161), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1162), .A2(KEYINPUT118), .A3(G8), .A4(new_n1144), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1142), .B(new_n1151), .C1(new_n1158), .C2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(KEYINPUT126), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1121), .A2(new_n1141), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1162), .A2(G8), .A3(new_n1144), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT118), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1168), .B1(new_n1171), .B2(new_n1163), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1167), .B1(new_n1172), .B2(new_n1151), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1081), .B(new_n1112), .C1(new_n1166), .C2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g749(.A(G1976), .B(G288), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1129), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1136), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1157), .A2(new_n1144), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1107), .A2(new_n1093), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(G168), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n1178), .A2(new_n1168), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1177), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1151), .A2(new_n1182), .A3(G168), .A4(new_n1179), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1171), .A2(new_n1163), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1168), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1174), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1165), .A2(KEYINPUT126), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1172), .A2(new_n1167), .A3(new_n1151), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1104), .A2(new_n1192), .A3(new_n1108), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1194));
  OAI211_X1 g769(.A(G171), .B(new_n1111), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1191), .A2(KEYINPUT127), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT127), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1188), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1022), .B1(new_n716), .B2(new_n714), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n1009), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1020), .A2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1034), .B1(new_n1199), .B2(new_n1202), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g778(.A(G227), .ZN(new_n1205));
  OAI21_X1  g779(.A(new_n1205), .B1(new_n647), .B2(new_n648), .ZN(new_n1206));
  AOI21_X1  g780(.A(new_n1206), .B1(new_n922), .B2(new_n923), .ZN(new_n1207));
  NAND4_X1  g781(.A1(new_n1207), .A2(G319), .A3(new_n681), .A4(new_n996), .ZN(G225));
  INV_X1    g782(.A(G225), .ZN(G308));
endmodule


