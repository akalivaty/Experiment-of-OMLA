//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n454), .B(new_n455), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n465), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  AOI211_X1 g049(.A(KEYINPUT68), .B(new_n474), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n476), .B1(new_n468), .B2(KEYINPUT3), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n466), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n477), .A2(new_n478), .A3(new_n474), .A4(new_n469), .ZN(new_n479));
  INV_X1    g054(.A(G137), .ZN(new_n480));
  INV_X1    g055(.A(G101), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n474), .A2(G2104), .ZN(new_n482));
  OAI22_X1  g057(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR3_X1   g058(.A1(new_n473), .A2(new_n475), .A3(new_n483), .ZN(G160));
  AND4_X1   g059(.A1(new_n474), .A2(new_n477), .A3(new_n478), .A4(new_n469), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n474), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n477), .A2(new_n478), .A3(G2105), .A4(new_n469), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(KEYINPUT70), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n493), .B2(G124), .ZN(new_n494));
  XNOR2_X1  g069(.A(new_n494), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n477), .A2(new_n478), .A3(new_n497), .A4(new_n469), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT3), .B(G2104), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n498), .A2(KEYINPUT4), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(G114), .B2(new_n474), .ZN(new_n504));
  INV_X1    g079(.A(G126), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n490), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n501), .A2(new_n506), .ZN(G164));
  AND2_X1   g082(.A1(KEYINPUT72), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT72), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n514), .A2(new_n515), .B1(G75), .B2(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(KEYINPUT73), .A3(G62), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n510), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  OR2_X1    g095(.A1(KEYINPUT72), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT72), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(G543), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n513), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n519), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n518), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT6), .B1(new_n508), .B2(new_n509), .ZN(new_n533));
  INV_X1    g108(.A(new_n524), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G89), .ZN(new_n536));
  INV_X1    g111(.A(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n533), .B2(new_n534), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(KEYINPUT7), .ZN(new_n542));
  AND2_X1   g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n513), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n536), .A2(new_n539), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n536), .A2(new_n539), .A3(new_n547), .A4(new_n544), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(G168));
  NAND2_X1  g124(.A1(new_n535), .A2(G90), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n538), .A2(G52), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G64), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n532), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n510), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  NAND2_X1  g133(.A1(new_n535), .A2(G81), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n538), .A2(G43), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n532), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(new_n555), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n559), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  OAI211_X1 g146(.A(G53), .B(G543), .C1(new_n523), .C2(new_n524), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n538), .A2(new_n574), .A3(G53), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n532), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n535), .A2(G91), .B1(new_n579), .B2(G651), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI211_X1 g158(.A(G87), .B(new_n513), .C1(new_n523), .C2(new_n524), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n538), .A2(G49), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G288));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n511), .B2(new_n512), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT75), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n590), .B2(KEYINPUT75), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n555), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT76), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n597));
  OAI211_X1 g172(.A(new_n597), .B(new_n555), .C1(new_n592), .C2(new_n594), .ZN(new_n598));
  AOI22_X1  g173(.A1(G48), .A2(new_n538), .B1(new_n535), .B2(G86), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(G305));
  NAND2_X1  g175(.A1(new_n535), .A2(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n538), .A2(G47), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  OAI211_X1 g178(.A(new_n601), .B(new_n602), .C1(new_n510), .C2(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G54), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G651), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n525), .A2(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n535), .A2(G92), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n605), .B1(new_n616), .B2(G868), .ZN(G284));
  XOR2_X1   g192(.A(G284), .B(KEYINPUT78), .Z(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G286), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(G299), .B(KEYINPUT79), .Z(new_n621));
  AOI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G297));
  AOI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n619), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(new_n624), .B2(G860), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT80), .Z(G148));
  NAND2_X1  g201(.A1(new_n616), .A2(new_n624), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OR3_X1    g203(.A1(new_n628), .A2(KEYINPUT81), .A3(new_n619), .ZN(new_n629));
  OAI21_X1  g204(.A(KEYINPUT81), .B1(new_n628), .B2(new_n619), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n629), .B(new_n630), .C1(G868), .C2(new_n566), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n493), .A2(G123), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G111), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G2105), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n636), .B1(new_n485), .B2(G135), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n474), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT12), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT13), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n649), .B2(new_n648), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(G401));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n661), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2100), .ZN(new_n668));
  XOR2_X1   g243(.A(G2072), .B(G2078), .Z(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(KEYINPUT18), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  AND2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  MUX2_X1   g257(.A(new_n682), .B(new_n681), .S(new_n674), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1991), .B(G1996), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NOR2_X1   g268(.A1(G286), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT94), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g271(.A(KEYINPUT94), .B1(G16), .B2(G21), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT96), .B(G1966), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT95), .Z(new_n700));
  XOR2_X1   g275(.A(new_n698), .B(new_n700), .Z(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G26), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n493), .A2(G128), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT87), .ZN(new_n706));
  NOR2_X1   g281(.A1(G104), .A2(G2105), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  INV_X1    g283(.A(G116), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n468), .B1(new_n709), .B2(G2105), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n485), .A2(G140), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n704), .B1(new_n712), .B2(new_n702), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G2067), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n702), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n702), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT29), .B(G2090), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n701), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT31), .B(G11), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT30), .B(G28), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n702), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n638), .B2(new_n702), .ZN(new_n723));
  NAND2_X1  g298(.A1(G171), .A2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G5), .B2(G16), .ZN(new_n725));
  INV_X1    g300(.A(G1961), .ZN(new_n726));
  INV_X1    g301(.A(G1341), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n693), .A2(G19), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n565), .B2(G16), .ZN(new_n729));
  OAI22_X1  g304(.A1(new_n725), .A2(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n723), .B(new_n730), .C1(new_n727), .C2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n702), .A2(G33), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n733));
  NAND3_X1  g308(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n485), .A2(G139), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n735), .B(new_n736), .C1(new_n474), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT90), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n702), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n731), .B1(G2072), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n693), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT98), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n702), .B1(KEYINPUT24), .B2(G34), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(KEYINPUT24), .B2(G34), .ZN(new_n748));
  INV_X1    g323(.A(G160), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT97), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  NAND2_X1  g329(.A1(G164), .A2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G27), .B2(G29), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n725), .A2(new_n726), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n757), .B1(new_n754), .B2(new_n756), .C1(new_n751), .C2(new_n750), .ZN(new_n758));
  NOR4_X1   g333(.A1(new_n741), .A2(new_n746), .A3(new_n753), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n474), .A2(G105), .A3(G2104), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n762), .B(new_n763), .Z(new_n764));
  AOI211_X1 g339(.A(new_n761), .B(new_n764), .C1(G141), .C2(new_n485), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n493), .A2(G129), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n702), .A2(G32), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(KEYINPUT27), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(KEYINPUT27), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G1996), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n740), .A2(G2072), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT91), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n693), .A2(G4), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n616), .B2(new_n693), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1348), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n719), .A2(new_n759), .A3(new_n775), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n693), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n693), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT85), .ZN(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(G305), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G16), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G6), .B2(G16), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  AOI22_X1  g366(.A1(new_n785), .A2(new_n786), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n693), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n693), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT33), .B(G1976), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n790), .A2(new_n791), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n787), .A2(new_n792), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n799), .A2(new_n801), .ZN(new_n803));
  MUX2_X1   g378(.A(G24), .B(G290), .S(G16), .Z(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1986), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n485), .A2(G131), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n474), .A2(G107), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n491), .A2(new_n492), .ZN(new_n809));
  INV_X1    g384(.A(G119), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n806), .B1(new_n807), .B2(new_n808), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  MUX2_X1   g386(.A(G25), .B(new_n811), .S(G29), .Z(new_n812));
  XOR2_X1   g387(.A(KEYINPUT35), .B(G1991), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT82), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT83), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n805), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT86), .B(KEYINPUT36), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n802), .A2(new_n803), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n802), .A2(new_n803), .A3(new_n818), .ZN(new_n821));
  INV_X1    g396(.A(new_n819), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n782), .B1(new_n820), .B2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n820), .ZN(new_n825));
  INV_X1    g400(.A(new_n782), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n825), .B2(new_n826), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(G150));
  NAND2_X1  g405(.A1(G80), .A2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G67), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n532), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n555), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n837), .A2(new_n525), .B1(new_n526), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT102), .B(G860), .Z(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n565), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n566), .A2(KEYINPUT101), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n840), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n844), .B(new_n565), .C1(new_n836), .C2(new_n839), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n616), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT39), .Z(new_n853));
  AND3_X1   g428(.A1(new_n853), .A2(KEYINPUT103), .A3(new_n841), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT103), .B1(new_n853), .B2(new_n841), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n843), .B1(new_n854), .B2(new_n855), .ZN(G145));
  XOR2_X1   g431(.A(KEYINPUT104), .B(G37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n485), .A2(G142), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n474), .A2(G118), .ZN(new_n859));
  OAI21_X1  g434(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(new_n493), .B2(G130), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(new_n642), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n811), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n706), .A2(new_n711), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G164), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(G164), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n767), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n865), .A2(G164), .ZN(new_n870));
  INV_X1    g445(.A(new_n767), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n866), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n869), .A2(new_n738), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n739), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n869), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n864), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(new_n638), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G160), .ZN(new_n878));
  NOR3_X1   g453(.A1(new_n867), .A2(new_n767), .A3(new_n868), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n871), .B1(new_n870), .B2(new_n866), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n739), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n864), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n869), .A2(new_n738), .A3(new_n872), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n876), .A2(new_n878), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n878), .B1(new_n876), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n857), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(G395));
  NAND2_X1  g464(.A1(new_n788), .A2(G166), .ZN(new_n890));
  NAND2_X1  g465(.A1(G303), .A2(G305), .ZN(new_n891));
  XOR2_X1   g466(.A(G288), .B(G290), .Z(new_n892));
  OAI211_X1 g467(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(KEYINPUT108), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(KEYINPUT108), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n893), .B(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT109), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT42), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n616), .A2(G299), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n615), .A2(new_n576), .A3(new_n580), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT106), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n902), .B1(new_n616), .B2(G299), .ZN(new_n903));
  OAI21_X1  g478(.A(KEYINPUT41), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n849), .B(new_n627), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n899), .A2(new_n900), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n905), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n901), .A2(new_n903), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT107), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(new_n908), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n898), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n898), .B1(new_n910), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n619), .B1(new_n836), .B2(new_n839), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(G295));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n918), .ZN(G331));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  XNOR2_X1  g496(.A(G168), .B(G301), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n849), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n849), .A2(new_n922), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n849), .A2(KEYINPUT110), .A3(new_n922), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n904), .A3(new_n907), .A4(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n912), .A2(new_n925), .A3(new_n923), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n929), .A3(new_n895), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n923), .A2(new_n925), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n906), .A2(KEYINPUT41), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n927), .A3(new_n926), .ZN(new_n934));
  AOI22_X1  g509(.A1(new_n923), .A2(new_n925), .B1(new_n906), .B2(KEYINPUT41), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n934), .A2(new_n912), .B1(KEYINPUT41), .B2(new_n935), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n857), .B(new_n930), .C1(new_n936), .C2(new_n895), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(new_n929), .ZN(new_n939));
  AOI21_X1  g514(.A(G37), .B1(new_n939), .B2(new_n896), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(new_n930), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n921), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n926), .A2(new_n927), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n912), .B1(new_n944), .B2(new_n935), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n935), .A2(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n895), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n930), .A2(new_n941), .ZN(new_n948));
  INV_X1    g523(.A(new_n857), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n941), .B1(new_n940), .B2(new_n930), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT44), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n943), .A2(new_n952), .ZN(G397));
  XOR2_X1   g528(.A(KEYINPUT111), .B(G1384), .Z(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n501), .B2(new_n506), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n482), .A2(new_n481), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n485), .B2(G137), .ZN(new_n959));
  INV_X1    g534(.A(new_n471), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n499), .B2(G125), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT68), .B1(new_n961), .B2(new_n474), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n472), .A2(new_n465), .A3(G2105), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n959), .A2(new_n962), .A3(new_n963), .A4(G40), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n957), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n774), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT46), .Z(new_n967));
  INV_X1    g542(.A(G2067), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n865), .B(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n871), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n967), .B1(new_n970), .B2(new_n965), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n971), .B(KEYINPUT47), .Z(new_n972));
  XNOR2_X1  g547(.A(new_n767), .B(new_n774), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n811), .A2(new_n814), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n974), .A2(new_n975), .B1(new_n968), .B2(new_n712), .ZN(new_n976));
  INV_X1    g551(.A(new_n965), .ZN(new_n977));
  OR3_X1    g552(.A1(new_n976), .A2(KEYINPUT126), .A3(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n811), .B(new_n814), .Z(new_n979));
  NAND2_X1  g554(.A1(new_n974), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n965), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n977), .A2(G1986), .A3(G290), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n982), .B(KEYINPUT48), .Z(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT126), .B1(new_n976), .B2(new_n977), .ZN(new_n985));
  AND4_X1   g560(.A1(new_n972), .A2(new_n978), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n987), .A2(new_n596), .A3(new_n598), .A4(new_n599), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n598), .A2(new_n599), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n987), .B1(new_n990), .B2(new_n596), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n991), .B2(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(G1981), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(new_n987), .A3(new_n596), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT49), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n501), .B2(new_n506), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n964), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n992), .A2(new_n995), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G288), .A2(G1976), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n988), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND4_X1   g577(.A1(G40), .A2(new_n959), .A3(new_n962), .A4(new_n963), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n997), .A2(new_n956), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n954), .C1(new_n501), .C2(new_n506), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n786), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n786), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n964), .B1(KEYINPUT50), .B2(new_n997), .ZN(new_n1011));
  INV_X1    g586(.A(G2090), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n996), .C1(new_n501), .C2(new_n506), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n1010), .A3(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(KEYINPUT55), .B(G8), .C1(new_n518), .C2(new_n528), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1017), .A2(KEYINPUT113), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(KEYINPUT113), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1020), .B1(G166), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1016), .A2(G8), .A3(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n586), .A2(KEYINPUT114), .A3(G1976), .A4(new_n587), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n587), .A2(G1976), .A3(new_n584), .A4(new_n585), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1976), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(G288), .B2(new_n1029), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n999), .A2(new_n1025), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT52), .B1(new_n1032), .B2(new_n998), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1000), .A2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1002), .A2(new_n998), .B1(new_n1024), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G114), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n502), .B1(new_n1037), .B2(G2105), .ZN(new_n1038));
  INV_X1    g613(.A(new_n490), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(G126), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n499), .A2(new_n500), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1384), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  NAND4_X1  g620(.A1(G160), .A2(new_n1044), .A3(new_n1045), .A4(G40), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT117), .B1(new_n964), .B2(new_n997), .ZN(new_n1047));
  XOR2_X1   g622(.A(KEYINPUT58), .B(G1341), .Z(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1003), .A2(new_n1004), .A3(new_n774), .A4(new_n1005), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n566), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n566), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1052), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1956), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT56), .B(G2072), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .A4(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n576), .B2(new_n580), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n574), .B1(new_n538), .B2(G53), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1061), .B(new_n580), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI22_X1  g641(.A1(new_n1057), .A2(new_n1060), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1003), .A2(new_n1068), .A3(new_n1014), .ZN(new_n1069));
  INV_X1    g644(.A(G1956), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1066), .A2(new_n1062), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1059), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n1075));
  AOI22_X1  g650(.A1(new_n1053), .A2(new_n1056), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(KEYINPUT120), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1071), .A2(new_n1072), .A3(new_n1078), .A4(new_n1059), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1077), .A2(KEYINPUT61), .A3(new_n1079), .A4(new_n1067), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT121), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1072), .B1(new_n1071), .B2(new_n1059), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1079), .A4(new_n1077), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1087), .A2(new_n968), .B1(new_n1088), .B2(new_n1069), .ZN(new_n1089));
  OR2_X1    g664(.A1(new_n1089), .A2(KEYINPUT60), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n968), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1069), .A2(new_n1088), .ZN(new_n1092));
  AND4_X1   g667(.A1(KEYINPUT60), .A2(new_n1091), .A3(new_n615), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n615), .B1(new_n1089), .B2(KEYINPUT60), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1090), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1076), .A2(new_n1081), .A3(new_n1086), .A4(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1089), .A2(new_n615), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1082), .B1(new_n1097), .B2(new_n1073), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1003), .A2(new_n1004), .A3(new_n754), .A4(new_n1005), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1069), .A2(new_n726), .ZN(new_n1103));
  OAI211_X1 g678(.A(KEYINPUT45), .B(new_n996), .C1(new_n501), .C2(new_n506), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1101), .A2(G2078), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1003), .A2(new_n1004), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(new_n1103), .A3(G301), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(G40), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n961), .A2(new_n474), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1108), .B(new_n1109), .C1(new_n1110), .C2(new_n483), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n957), .A3(new_n1005), .A4(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1102), .A2(new_n1103), .A3(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT54), .B(new_n1107), .C1(new_n1114), .C2(G301), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1021), .B1(new_n1015), .B2(new_n1007), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1023), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n993), .A2(new_n994), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n998), .B1(new_n1120), .B2(new_n989), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1119), .B1(new_n1121), .B2(new_n995), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1115), .A2(new_n1118), .A3(new_n1024), .A4(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1102), .A2(new_n1103), .A3(new_n1113), .A4(G301), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1102), .A2(new_n1106), .A3(new_n1103), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1124), .A2(KEYINPUT123), .B1(new_n1125), .B2(G171), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1124), .A2(KEYINPUT123), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT54), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1003), .A2(new_n1004), .A3(new_n1104), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n699), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1003), .A2(new_n1068), .A3(new_n751), .A4(new_n1014), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1130), .A2(G168), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1132), .A2(new_n1133), .A3(G8), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(G286), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(G8), .A3(new_n1132), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1134), .B1(new_n1137), .B2(KEYINPUT51), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1123), .A2(new_n1128), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1036), .B1(new_n1099), .B2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(new_n1021), .B(G286), .C1(new_n1130), .C2(new_n1131), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1118), .A2(new_n1024), .A3(new_n1122), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT115), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1035), .A2(new_n1117), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT115), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1144), .A2(new_n1145), .A3(new_n1024), .A4(new_n1141), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1016), .A2(G8), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1023), .A2(KEYINPUT116), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1141), .A2(KEYINPUT63), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1151), .A2(new_n1122), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1148), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1138), .A2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1125), .A2(G171), .ZN(new_n1158));
  AND4_X1   g733(.A1(new_n1024), .A2(new_n1118), .A3(new_n1122), .A4(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1132), .A2(G8), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1133), .B1(new_n1160), .B2(new_n1136), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT62), .B1(new_n1161), .B2(new_n1134), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1157), .A2(new_n1159), .A3(new_n1162), .A4(KEYINPUT124), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1140), .A2(new_n1155), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(G290), .B(G1986), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n965), .B1(new_n980), .B2(new_n1168), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1167), .A2(KEYINPUT125), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT125), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n986), .B1(new_n1170), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g747(.A1(G401), .A2(new_n463), .A3(G227), .ZN(new_n1174));
  OAI21_X1  g748(.A(new_n1174), .B1(new_n690), .B2(new_n691), .ZN(new_n1175));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1176));
  XNOR2_X1  g750(.A(new_n1175), .B(new_n1176), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n887), .B(new_n1177), .C1(new_n951), .C2(new_n950), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


