//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  AND3_X1   g001(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n188));
  AOI21_X1  g002(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G131), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G125), .B(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(KEYINPUT16), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  OR2_X1    g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(new_n193), .B(KEYINPUT19), .Z(new_n200));
  OAI211_X1 g014(.A(new_n192), .B(new_n199), .C1(G146), .C2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n190), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(KEYINPUT18), .A3(G131), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT18), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n190), .B1(new_n204), .B2(new_n191), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n193), .B(new_n198), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n203), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n201), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n208), .A2(KEYINPUT88), .ZN(new_n209));
  XNOR2_X1  g023(.A(G113), .B(G122), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n210), .B(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(new_n208), .B2(KEYINPUT88), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n197), .B(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(KEYINPUT17), .A3(G131), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n214), .B(new_n215), .C1(KEYINPUT17), .C2(new_n192), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n209), .A2(new_n213), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  INV_X1    g033(.A(G475), .ZN(new_n220));
  INV_X1    g034(.A(G902), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OR3_X1    g036(.A1(new_n219), .A2(KEYINPUT20), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT20), .B1(new_n219), .B2(new_n222), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n212), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT89), .ZN(new_n227));
  OR2_X1    g041(.A1(new_n217), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n227), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n221), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G475), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n234), .A2(G143), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT65), .A2(G134), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT65), .A2(G134), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n238), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT14), .A3(G122), .ZN(new_n244));
  XOR2_X1   g058(.A(G116), .B(G122), .Z(new_n245));
  OAI211_X1 g059(.A(G107), .B(new_n244), .C1(new_n245), .C2(KEYINPUT14), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n246), .A2(KEYINPUT92), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(G107), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n242), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n249), .B1(KEYINPUT92), .B2(new_n246), .ZN(new_n250));
  OR3_X1    g064(.A1(new_n238), .A2(new_n240), .A3(new_n239), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n245), .A2(G107), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n237), .B1(new_n253), .B2(new_n235), .ZN(new_n254));
  AOI211_X1 g068(.A(KEYINPUT91), .B(new_n254), .C1(new_n237), .C2(new_n253), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(KEYINPUT91), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G134), .ZN(new_n257));
  OAI221_X1 g071(.A(new_n251), .B1(new_n252), .B2(new_n248), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT9), .B(G234), .ZN(new_n260));
  INV_X1    g074(.A(G217), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n260), .A2(new_n261), .A3(G953), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n259), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n221), .ZN(new_n265));
  INV_X1    g079(.A(G478), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(KEYINPUT15), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n265), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n233), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n221), .B(new_n272), .C1(G234), .C2(G237), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT21), .B(G898), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g089(.A1(KEYINPUT93), .A2(G952), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT93), .A2(G952), .ZN(new_n277));
  AOI21_X1  g091(.A(G953), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G234), .ZN(new_n279));
  INV_X1    g093(.A(G237), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n271), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G214), .B1(G237), .B2(G902), .ZN(new_n284));
  INV_X1    g098(.A(G101), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT3), .B1(new_n211), .B2(G107), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n287));
  INV_X1    g101(.A(G107), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n288), .A3(G104), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n211), .A2(G107), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n286), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n285), .B1(new_n291), .B2(KEYINPUT82), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(KEYINPUT82), .B2(new_n291), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT4), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n291), .A2(G101), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n297), .B2(new_n294), .ZN(new_n298));
  XNOR2_X1  g112(.A(G116), .B(G119), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT2), .B(G113), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n299), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n304), .A2(new_n302), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n288), .A2(G104), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n285), .B1(new_n307), .B2(new_n290), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n308), .B(new_n309), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n310), .A2(new_n296), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT5), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n301), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n314), .A3(G116), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G113), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n305), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n298), .A2(new_n306), .B1(new_n311), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G122), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n320), .B(KEYINPUT85), .Z(new_n321));
  OR2_X1    g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n320), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT6), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT86), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n198), .A2(G143), .ZN(new_n327));
  INV_X1    g141(.A(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G146), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT64), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT0), .A2(G128), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT0), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(new_n234), .ZN(new_n336));
  INV_X1    g150(.A(new_n333), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(KEYINPUT64), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n334), .A2(new_n338), .B1(new_n336), .B2(new_n331), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G125), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n234), .B1(new_n327), .B2(KEYINPUT1), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n331), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n340), .B1(G125), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G224), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G953), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT87), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n344), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n322), .A2(KEYINPUT6), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n322), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n323), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n326), .A2(new_n349), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(G210), .B1(G237), .B2(G902), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT7), .B1(new_n345), .B2(G953), .ZN(new_n354));
  XOR2_X1   g168(.A(new_n344), .B(new_n354), .Z(new_n355));
  NAND2_X1  g169(.A1(new_n310), .A2(new_n296), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n318), .A2(new_n356), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n320), .B(KEYINPUT8), .Z(new_n358));
  NOR2_X1   g172(.A1(new_n304), .A2(new_n312), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n305), .B1(new_n359), .B2(new_n316), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n311), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n355), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(G902), .B1(new_n362), .B2(new_n323), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n352), .A2(new_n353), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n353), .B1(new_n352), .B2(new_n363), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n284), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G469), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n356), .B(new_n342), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT12), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT11), .ZN(new_n371));
  INV_X1    g185(.A(G134), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n371), .A2(new_n372), .A3(G137), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT65), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT65), .A2(G134), .ZN(new_n376));
  AOI21_X1  g190(.A(G137), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT66), .B1(new_n377), .B2(KEYINPUT11), .ZN(new_n378));
  INV_X1    g192(.A(G137), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n379), .B1(new_n239), .B2(new_n240), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n371), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n373), .B1(new_n378), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n375), .A2(G137), .A3(new_n376), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n191), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n191), .ZN(new_n386));
  AOI211_X1 g200(.A(new_n373), .B(new_n386), .C1(new_n378), .C2(new_n382), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OR3_X1    g202(.A1(new_n369), .A2(new_n370), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n370), .B1(new_n369), .B2(new_n388), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(KEYINPUT84), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n393), .B1(new_n389), .B2(new_n390), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n311), .A2(new_n342), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT10), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n298), .A2(new_n339), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n388), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n272), .A2(G227), .ZN(new_n400));
  XOR2_X1   g214(.A(new_n399), .B(new_n400), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n392), .A2(new_n394), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n388), .B1(new_n396), .B2(new_n397), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n402), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n368), .B(new_n221), .C1(new_n404), .C2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n402), .B1(new_n391), .B2(new_n398), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n398), .A3(new_n402), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(G469), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n368), .A2(new_n221), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G221), .B1(new_n260), .B2(G902), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT80), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n417), .B(KEYINPUT81), .Z(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n283), .A2(new_n367), .A3(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(G472), .A2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT32), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n306), .B(KEYINPUT70), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n339), .B1(new_n385), .B2(new_n387), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n379), .A2(G134), .ZN(new_n428));
  OAI21_X1  g242(.A(G131), .B1(new_n377), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n428), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n380), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT67), .A3(G131), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n373), .ZN(new_n436));
  INV_X1    g250(.A(new_n386), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n380), .A2(new_n381), .A3(new_n371), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n381), .B1(new_n380), .B2(new_n371), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n435), .A2(new_n440), .A3(new_n342), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n427), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n426), .B1(new_n442), .B2(KEYINPUT73), .ZN(new_n443));
  INV_X1    g257(.A(new_n339), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n436), .B1(new_n438), .B2(new_n439), .ZN(new_n445));
  INV_X1    g259(.A(new_n384), .ZN(new_n446));
  OAI21_X1  g260(.A(G131), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n444), .B1(new_n447), .B2(new_n440), .ZN(new_n448));
  INV_X1    g262(.A(new_n441), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT73), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT28), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT72), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n435), .A2(new_n440), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n343), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n435), .A2(new_n440), .A3(KEYINPUT68), .ZN(new_n456));
  AOI211_X1 g270(.A(new_n373), .B(new_n446), .C1(new_n378), .C2(new_n382), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n440), .B1(new_n457), .B2(new_n191), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n455), .A2(new_n456), .B1(new_n458), .B2(new_n339), .ZN(new_n459));
  INV_X1    g273(.A(new_n306), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n452), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n426), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n427), .A3(new_n441), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n435), .A2(new_n440), .A3(KEYINPUT68), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT68), .B1(new_n435), .B2(new_n440), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n464), .A2(new_n465), .A3(new_n343), .ZN(new_n466));
  OAI211_X1 g280(.A(KEYINPUT72), .B(new_n306), .C1(new_n466), .C2(new_n448), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n463), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n451), .B1(new_n468), .B2(KEYINPUT28), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n187), .A2(G210), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT27), .Z(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT26), .B(G101), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n471), .B(new_n472), .Z(new_n473));
  OAI21_X1  g287(.A(KEYINPUT74), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT74), .ZN(new_n475));
  INV_X1    g289(.A(new_n473), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n442), .A2(new_n426), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT67), .B1(new_n433), .B2(G131), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n430), .B(new_n191), .C1(new_n380), .C2(new_n432), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n454), .B1(new_n387), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n342), .A3(new_n456), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n460), .B1(new_n483), .B2(new_n427), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n478), .B1(KEYINPUT72), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n477), .B1(new_n485), .B2(new_n461), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n475), .B(new_n476), .C1(new_n486), .C2(new_n451), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n474), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n483), .A2(new_n490), .A3(new_n427), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT30), .B1(new_n448), .B2(new_n449), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n478), .B1(new_n493), .B2(new_n306), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n489), .B1(new_n494), .B2(new_n473), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n460), .B1(new_n491), .B2(new_n492), .ZN(new_n496));
  NOR4_X1   g310(.A1(new_n496), .A2(KEYINPUT71), .A3(new_n478), .A4(new_n476), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT31), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n490), .B1(new_n427), .B2(new_n441), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n459), .B2(new_n490), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n463), .B(new_n473), .C1(new_n500), .C2(new_n460), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT31), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n488), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n505), .B1(new_n488), .B2(new_n504), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n425), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n494), .A2(new_n473), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(KEYINPUT29), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n467), .A2(new_n463), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n484), .A2(KEYINPUT72), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT28), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n451), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n510), .B1(new_n476), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g330(.A1(new_n514), .A2(KEYINPUT76), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n462), .B(new_n442), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT76), .B1(new_n518), .B2(new_n477), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n519), .B2(new_n451), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n473), .A2(KEYINPUT29), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n516), .A2(new_n221), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G472), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n475), .B1(new_n515), .B2(new_n476), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n469), .A2(KEYINPUT74), .A3(new_n473), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n501), .A2(KEYINPUT71), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n494), .A2(new_n489), .A3(new_n473), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n502), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n503), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n526), .A2(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n488), .A2(new_n504), .A3(new_n505), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n423), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n508), .B(new_n525), .C1(new_n535), .C2(KEYINPUT32), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n234), .A2(G119), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT23), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n314), .A2(G128), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n234), .A2(KEYINPUT23), .A3(G119), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT24), .B(G110), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AND2_X1   g358(.A1(new_n540), .A2(new_n537), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n542), .A2(G110), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n193), .A2(new_n198), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n199), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n542), .A2(G110), .ZN(new_n549));
  INV_X1    g363(.A(new_n545), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n543), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n548), .B1(new_n214), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT22), .B(G137), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n552), .B(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(G902), .B1(new_n279), .B2(G217), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT78), .Z(new_n559));
  OAI21_X1  g373(.A(G217), .B1(new_n279), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT25), .ZN(new_n561));
  AOI21_X1  g375(.A(G902), .B1(new_n561), .B2(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(KEYINPUT77), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n564), .B2(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n536), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT79), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT79), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n536), .A2(new_n571), .A3(new_n568), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n421), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(new_n285), .ZN(G3));
  OAI21_X1  g388(.A(new_n221), .B1(new_n506), .B2(new_n507), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n535), .B1(G472), .B2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n415), .A2(new_n418), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n576), .A2(new_n568), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n262), .B1(new_n250), .B2(new_n258), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT33), .B1(new_n579), .B2(KEYINPUT94), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n264), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n266), .A2(new_n221), .ZN(new_n583));
  INV_X1    g397(.A(new_n265), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n583), .B1(new_n584), .B2(new_n266), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n232), .ZN(new_n588));
  INV_X1    g402(.A(new_n284), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n352), .A2(new_n363), .ZN(new_n590));
  INV_X1    g404(.A(new_n353), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n589), .B1(new_n592), .B2(new_n364), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n282), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n578), .A2(new_n588), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT34), .B(G104), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(G6));
  OR2_X1    g411(.A1(new_n223), .A2(KEYINPUT95), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n223), .A2(KEYINPUT95), .A3(new_n224), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n268), .A2(new_n598), .A3(new_n231), .A4(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n578), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G107), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  INV_X1    g417(.A(new_n555), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(KEYINPUT36), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n552), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n557), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n566), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n283), .A2(new_n367), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n576), .A2(new_n577), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT37), .B(G110), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  INV_X1    g427(.A(new_n281), .ZN(new_n614));
  INV_X1    g428(.A(G900), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n615), .B2(new_n273), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n230), .B2(G475), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n268), .A2(new_n598), .A3(new_n599), .A4(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n577), .A2(new_n593), .A3(new_n608), .A4(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n533), .A2(new_n534), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n621), .A2(new_n425), .B1(G472), .B2(new_n524), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n422), .B1(new_n506), .B2(new_n507), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n424), .ZN(new_n624));
  AOI211_X1 g438(.A(KEYINPUT96), .B(new_n620), .C1(new_n622), .C2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n626));
  INV_X1    g440(.A(new_n620), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n536), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(new_n234), .ZN(G30));
  XOR2_X1   g444(.A(new_n616), .B(KEYINPUT39), .Z(new_n631));
  NAND2_X1  g445(.A1(new_n577), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(new_n632), .B(KEYINPUT40), .Z(new_n633));
  NAND2_X1  g447(.A1(new_n592), .A2(new_n364), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT38), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n233), .A2(new_n269), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n608), .A2(new_n589), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n633), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G472), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n528), .B(new_n529), .C1(new_n473), .C2(new_n518), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n639), .B1(new_n640), .B2(new_n221), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n621), .B2(new_n425), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(new_n624), .A3(KEYINPUT97), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT97), .B1(new_n642), .B2(new_n624), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n638), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n328), .ZN(G45));
  NOR3_X1   g462(.A1(new_n588), .A2(new_n609), .A3(new_n616), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n536), .A2(new_n577), .A3(new_n593), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G146), .ZN(G48));
  NOR2_X1   g465(.A1(new_n594), .A2(new_n588), .ZN(new_n652));
  INV_X1    g466(.A(new_n407), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n403), .A2(new_n394), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n653), .B1(new_n392), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n221), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(G469), .ZN(new_n657));
  INV_X1    g471(.A(new_n417), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n408), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n536), .A2(new_n568), .A3(new_n652), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT41), .B(G113), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G15));
  NOR2_X1   g477(.A1(new_n594), .A2(new_n600), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n536), .A2(new_n568), .A3(new_n664), .A4(new_n660), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  NOR4_X1   g480(.A1(new_n283), .A2(new_n659), .A3(new_n367), .A4(new_n609), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n536), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G119), .ZN(G21));
  NAND2_X1  g483(.A1(new_n593), .A2(new_n636), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n275), .A2(new_n281), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n670), .A2(new_n671), .A3(new_n659), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n520), .A2(new_n473), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n423), .B1(new_n673), .B2(new_n504), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n575), .B2(G472), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n672), .A2(new_n675), .A3(new_n568), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT98), .B(G122), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G24));
  NOR2_X1   g492(.A1(new_n659), .A2(new_n367), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n675), .A2(new_n649), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G125), .ZN(G27));
  NAND2_X1  g495(.A1(new_n569), .A2(KEYINPUT102), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n536), .A2(new_n683), .A3(new_n568), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n412), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n410), .A2(KEYINPUT99), .A3(G469), .A4(new_n411), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n408), .A2(new_n686), .A3(new_n414), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n658), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n689), .A2(KEYINPUT100), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n688), .B2(new_n658), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n592), .A2(new_n284), .A3(new_n364), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n588), .A2(new_n616), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n694), .A2(KEYINPUT42), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n682), .A2(new_n684), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n536), .A2(new_n694), .A3(new_n568), .A4(new_n695), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT103), .B(G131), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G33));
  NAND4_X1  g519(.A1(new_n536), .A2(new_n694), .A3(new_n568), .A4(new_n619), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G134), .ZN(G36));
  NOR2_X1   g521(.A1(new_n586), .A2(new_n232), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT43), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n608), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n576), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(KEYINPUT105), .Z(new_n713));
  NOR2_X1   g527(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT106), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(KEYINPUT106), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n410), .A2(KEYINPUT45), .A3(new_n411), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n403), .A2(new_n405), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n718), .B1(new_n719), .B2(new_n409), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n720), .A3(G469), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT104), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n717), .A2(new_n720), .A3(KEYINPUT104), .A4(G469), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n413), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n408), .A3(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n658), .A3(new_n631), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n693), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n713), .A2(new_n715), .A3(new_n716), .A4(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT107), .B(G137), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(G39));
  NAND2_X1  g547(.A1(new_n728), .A2(new_n658), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT47), .ZN(new_n735));
  INV_X1    g549(.A(new_n693), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n695), .A2(new_n736), .A3(new_n567), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n735), .A2(new_n536), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n195), .ZN(G42));
  AND2_X1   g553(.A1(new_n657), .A2(new_n408), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n741), .A2(KEYINPUT49), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(KEYINPUT49), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n708), .A2(new_n568), .A3(new_n418), .A4(new_n284), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n742), .A2(new_n743), .A3(new_n635), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n646), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n709), .A2(new_n614), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n660), .A3(new_n736), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT112), .ZN(new_n749));
  AND2_X1   g563(.A1(new_n682), .A2(new_n684), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n751), .B(KEYINPUT48), .Z(new_n752));
  AOI211_X1 g566(.A(new_n567), .B(new_n674), .C1(new_n575), .C2(G472), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n679), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n659), .A2(new_n693), .A3(new_n567), .A4(new_n281), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n646), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n278), .B(new_n755), .C1(new_n757), .C2(new_n588), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n757), .A2(new_n232), .A3(new_n587), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n749), .A2(new_n608), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n675), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n735), .B1(new_n418), .B2(new_n741), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n754), .A2(KEYINPUT111), .A3(new_n736), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n765));
  INV_X1    g579(.A(new_n754), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n765), .B1(new_n766), .B2(new_n693), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n635), .A2(new_n284), .A3(new_n659), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n754), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT50), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n762), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n759), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n650), .B(new_n680), .C1(new_n625), .C2(new_n628), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n616), .B(KEYINPUT110), .Z(new_n779));
  NOR4_X1   g593(.A1(new_n670), .A2(new_n608), .A3(new_n689), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n645), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(new_n643), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT52), .B1(new_n778), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n680), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT32), .B1(new_n621), .B2(new_n422), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n508), .A2(new_n525), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n627), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT96), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n536), .A2(new_n626), .A3(new_n627), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n780), .B1(new_n644), .B2(new_n645), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n650), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n598), .A2(new_n599), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n269), .A2(new_n608), .A3(new_n617), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n419), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n536), .A2(new_n736), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n694), .A2(new_n675), .A3(new_n649), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n706), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n703), .A2(new_n784), .A3(new_n794), .A4(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n661), .A2(new_n665), .A3(new_n668), .A4(new_n676), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT108), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n753), .A2(new_n672), .B1(new_n667), .B2(new_n536), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT108), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n805), .A3(new_n661), .A4(new_n665), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n270), .B1(new_n587), .B2(new_n233), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n594), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n576), .A2(new_n810), .A3(new_n568), .A4(new_n577), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n611), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n808), .B1(new_n573), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n572), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n571), .B1(new_n536), .B2(new_n568), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n420), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(KEYINPUT109), .A3(new_n611), .A4(new_n811), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n807), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n801), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n813), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n791), .A2(new_n792), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n804), .A2(KEYINPUT53), .A3(new_n661), .A4(new_n665), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n784), .A2(new_n794), .A3(new_n703), .A4(new_n800), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n820), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n819), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n801), .B(new_n818), .C1(KEYINPUT53), .C2(new_n822), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  INV_X1    g644(.A(new_n807), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n821), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n832), .B2(new_n826), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n828), .B1(KEYINPUT54), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n777), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(G952), .A2(G953), .ZN(new_n837));
  OAI211_X1 g651(.A(KEYINPUT113), .B(new_n746), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT113), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n777), .B2(new_n835), .ZN(new_n840));
  INV_X1    g654(.A(new_n746), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(G75));
  NOR2_X1   g657(.A1(new_n272), .A2(G952), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n844), .B(KEYINPUT116), .Z(new_n845));
  AND2_X1   g659(.A1(new_n784), .A2(new_n794), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n703), .A2(new_n800), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n821), .A4(new_n824), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(G902), .ZN(new_n850));
  INV_X1    g664(.A(G210), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n326), .A2(new_n350), .A3(new_n351), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT114), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n348), .B(KEYINPUT55), .Z(new_n855));
  XNOR2_X1  g669(.A(new_n854), .B(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n845), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  OR3_X1    g672(.A1(new_n850), .A2(KEYINPUT115), .A3(new_n851), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n850), .B2(new_n851), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n862), .B2(new_n856), .ZN(G51));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n819), .B2(new_n827), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n825), .A2(new_n826), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n819), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n833), .A2(KEYINPUT117), .A3(new_n820), .A4(new_n848), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n413), .B(KEYINPUT57), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n870), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n655), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n850), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n723), .A3(new_n724), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n844), .B1(new_n875), .B2(new_n877), .ZN(G54));
  NAND3_X1  g692(.A1(new_n876), .A2(KEYINPUT58), .A3(G475), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n879), .A2(new_n219), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n219), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n880), .A2(new_n881), .A3(new_n844), .ZN(G60));
  XNOR2_X1  g696(.A(new_n583), .B(KEYINPUT59), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n581), .B1(new_n835), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n845), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n581), .A2(new_n883), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n869), .B2(new_n886), .ZN(G63));
  NAND2_X1  g701(.A1(G217), .A2(G902), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT120), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n889), .B(new_n890), .Z(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n833), .B2(new_n848), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n556), .B(KEYINPUT121), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n606), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n845), .A3(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT61), .Z(G66));
  NOR2_X1   g712(.A1(new_n818), .A2(G953), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT122), .ZN(new_n900));
  OAI21_X1  g714(.A(G953), .B1(new_n274), .B2(new_n345), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(G898), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n854), .B1(new_n904), .B2(G953), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n903), .B(new_n905), .Z(G69));
  INV_X1    g720(.A(new_n778), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n729), .A2(new_n670), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n750), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n706), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n738), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n731), .A2(new_n907), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n703), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT125), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n911), .A2(new_n909), .A3(new_n907), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n703), .A4(new_n731), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n917), .A3(new_n272), .ZN(new_n918));
  NAND2_X1  g732(.A1(G900), .A2(G953), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n500), .B(new_n200), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(G227), .A2(G900), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(G953), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n570), .A2(new_n572), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n632), .A2(new_n693), .A3(new_n809), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n738), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR3_X1    g741(.A1(new_n647), .A2(new_n778), .A3(KEYINPUT62), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT62), .B1(new_n647), .B2(new_n778), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n927), .A2(new_n731), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(KEYINPUT124), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(KEYINPUT124), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n921), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(new_n272), .A3(new_n934), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n922), .A2(new_n924), .A3(new_n935), .ZN(new_n936));
  AND4_X1   g750(.A1(G953), .A2(new_n920), .A3(new_n923), .A4(new_n921), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(G72));
  INV_X1    g752(.A(new_n844), .ZN(new_n939));
  NAND2_X1  g753(.A1(G472), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT63), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n528), .A2(new_n529), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n834), .B(new_n941), .C1(new_n942), .C2(new_n509), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n914), .A2(new_n917), .A3(new_n818), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n944), .A2(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n494), .A2(new_n476), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT127), .Z(new_n947));
  OAI211_X1 g761(.A(new_n939), .B(new_n943), .C1(new_n945), .C2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n931), .A2(new_n932), .A3(new_n818), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n941), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n949), .A2(new_n952), .A3(new_n941), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n494), .A2(new_n476), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(G57));
endmodule


