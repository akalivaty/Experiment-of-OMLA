

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U554 ( .A(n700), .ZN(n732) );
  NOR2_X1 U555 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U556 ( .A1(n799), .A2(n798), .ZN(n520) );
  INV_X1 U557 ( .A(KEYINPUT96), .ZN(n706) );
  NOR2_X1 U558 ( .A1(n746), .A2(n993), .ZN(n751) );
  NAND2_X1 U559 ( .A1(n520), .A2(n804), .ZN(n805) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  NOR2_X1 U561 ( .A1(G651), .A2(n646), .ZN(n653) );
  NOR2_X1 U562 ( .A1(G543), .A2(G651), .ZN(n649) );
  NAND2_X1 U563 ( .A1(n896), .A2(G137), .ZN(n538) );
  NOR2_X1 U564 ( .A1(n545), .A2(n544), .ZN(G160) );
  XNOR2_X1 U565 ( .A(KEYINPUT7), .B(KEYINPUT80), .ZN(n535) );
  XOR2_X1 U566 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  NAND2_X1 U567 ( .A1(G51), .A2(n653), .ZN(n523) );
  INV_X1 U568 ( .A(G651), .ZN(n527) );
  NOR2_X1 U569 ( .A1(G543), .A2(n527), .ZN(n521) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n521), .Z(n654) );
  NAND2_X1 U571 ( .A1(G63), .A2(n654), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U573 ( .A(n524), .B(KEYINPUT79), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n525), .B(KEYINPUT6), .ZN(n533) );
  XNOR2_X1 U575 ( .A(KEYINPUT5), .B(KEYINPUT78), .ZN(n531) );
  NAND2_X1 U576 ( .A1(n649), .A2(G89), .ZN(n526) );
  XNOR2_X1 U577 ( .A(n526), .B(KEYINPUT4), .ZN(n529) );
  NOR2_X1 U578 ( .A1(n646), .A2(n527), .ZN(n650) );
  NAND2_X1 U579 ( .A1(G76), .A2(n650), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U581 ( .A(n531), .B(n530), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U583 ( .A(n535), .B(n534), .ZN(G168) );
  XOR2_X1 U584 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  AND2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n900) );
  NAND2_X1 U586 ( .A1(G113), .A2(n900), .ZN(n539) );
  XOR2_X1 U587 ( .A(KEYINPUT66), .B(n536), .Z(n537) );
  XNOR2_X2 U588 ( .A(n537), .B(KEYINPUT17), .ZN(n896) );
  NAND2_X1 U589 ( .A1(n539), .A2(n538), .ZN(n545) );
  XNOR2_X1 U590 ( .A(KEYINPUT65), .B(G2104), .ZN(n558) );
  NOR2_X1 U591 ( .A1(G2105), .A2(n558), .ZN(n610) );
  NAND2_X1 U592 ( .A1(G101), .A2(n610), .ZN(n541) );
  INV_X1 U593 ( .A(KEYINPUT23), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n541), .B(n540), .ZN(n543) );
  AND2_X1 U595 ( .A1(n558), .A2(G2105), .ZN(n903) );
  NAND2_X1 U596 ( .A1(n903), .A2(G125), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n544) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  INV_X1 U601 ( .A(G120), .ZN(G236) );
  INV_X1 U602 ( .A(G69), .ZN(G235) );
  INV_X1 U603 ( .A(G108), .ZN(G238) );
  NAND2_X1 U604 ( .A1(G90), .A2(n649), .ZN(n547) );
  NAND2_X1 U605 ( .A1(G77), .A2(n650), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT70), .B(KEYINPUT9), .Z(n548) );
  XNOR2_X1 U608 ( .A(n549), .B(n548), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G52), .A2(n653), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G64), .A2(n654), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U612 ( .A(KEYINPUT69), .B(n552), .Z(n553) );
  NOR2_X1 U613 ( .A1(n554), .A2(n553), .ZN(G171) );
  NAND2_X1 U614 ( .A1(G138), .A2(n896), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n610), .A2(G102), .ZN(n555) );
  NAND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n564) );
  AND2_X1 U617 ( .A1(G2105), .A2(G126), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U619 ( .A(KEYINPUT89), .B(n559), .Z(n561) );
  NAND2_X1 U620 ( .A1(n900), .A2(G114), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT90), .ZN(n563) );
  NOR2_X1 U623 ( .A1(n564), .A2(n563), .ZN(G164) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(KEYINPUT74), .Z(n568) );
  XOR2_X1 U625 ( .A(KEYINPUT10), .B(KEYINPUT73), .Z(n566) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n565) );
  XOR2_X1 U627 ( .A(n566), .B(n565), .Z(n829) );
  NAND2_X1 U628 ( .A1(G567), .A2(n829), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n568), .B(n567), .ZN(G234) );
  NAND2_X1 U630 ( .A1(n653), .A2(G43), .ZN(n569) );
  XNOR2_X1 U631 ( .A(KEYINPUT76), .B(n569), .ZN(n579) );
  XNOR2_X1 U632 ( .A(KEYINPUT75), .B(KEYINPUT13), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n649), .A2(G81), .ZN(n570) );
  XNOR2_X1 U634 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G68), .A2(n650), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(n574), .B(n573), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n654), .A2(G56), .ZN(n575) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n575), .Z(n576) );
  NOR2_X1 U640 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n579), .A2(n578), .ZN(n977) );
  INV_X1 U642 ( .A(G860), .ZN(n600) );
  OR2_X1 U643 ( .A1(n977), .A2(n600), .ZN(G153) );
  INV_X1 U644 ( .A(G171), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U646 ( .A1(G92), .A2(n649), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G66), .A2(n654), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G54), .A2(n653), .ZN(n583) );
  NAND2_X1 U650 ( .A1(G79), .A2(n650), .ZN(n582) );
  NAND2_X1 U651 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U652 ( .A(KEYINPUT77), .B(n584), .Z(n585) );
  NOR2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n587), .Z(n973) );
  OR2_X1 U655 ( .A1(n973), .A2(G868), .ZN(n588) );
  NAND2_X1 U656 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G53), .A2(n653), .ZN(n591) );
  NAND2_X1 U658 ( .A1(G65), .A2(n654), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U660 ( .A(KEYINPUT72), .B(n592), .ZN(n595) );
  NAND2_X1 U661 ( .A1(G78), .A2(n650), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT71), .B(n593), .ZN(n594) );
  NOR2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n649), .A2(G91), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n597), .A2(n596), .ZN(G299) );
  NAND2_X1 U666 ( .A1(G868), .A2(G286), .ZN(n599) );
  INV_X1 U667 ( .A(G299), .ZN(n712) );
  OR2_X1 U668 ( .A1(n712), .A2(G868), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U671 ( .A1(n601), .A2(n973), .ZN(n602) );
  XNOR2_X1 U672 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n977), .ZN(n605) );
  NAND2_X1 U674 ( .A1(G868), .A2(n973), .ZN(n603) );
  NOR2_X1 U675 ( .A1(G559), .A2(n603), .ZN(n604) );
  NOR2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X1 U677 ( .A(KEYINPUT81), .B(n606), .Z(G282) );
  NAND2_X1 U678 ( .A1(n903), .A2(G123), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G111), .A2(n900), .ZN(n608) );
  NAND2_X1 U681 ( .A1(n609), .A2(n608), .ZN(n615) );
  INV_X1 U682 ( .A(n610), .ZN(n611) );
  INV_X1 U683 ( .A(n611), .ZN(n894) );
  NAND2_X1 U684 ( .A1(n894), .A2(G99), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G135), .A2(n896), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n922) );
  XNOR2_X1 U688 ( .A(n922), .B(G2096), .ZN(n616) );
  INV_X1 U689 ( .A(G2100), .ZN(n849) );
  NAND2_X1 U690 ( .A1(n616), .A2(n849), .ZN(G156) );
  NAND2_X1 U691 ( .A1(n973), .A2(G559), .ZN(n666) );
  XNOR2_X1 U692 ( .A(n977), .B(n666), .ZN(n617) );
  NOR2_X1 U693 ( .A1(n617), .A2(G860), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G55), .A2(n653), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G67), .A2(n654), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G93), .A2(n649), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G80), .A2(n650), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n668) );
  XNOR2_X1 U701 ( .A(n624), .B(n668), .ZN(G145) );
  NAND2_X1 U702 ( .A1(n653), .A2(G47), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n625), .B(KEYINPUT68), .ZN(n632) );
  NAND2_X1 U704 ( .A1(G85), .A2(n649), .ZN(n627) );
  NAND2_X1 U705 ( .A1(G72), .A2(n650), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G60), .A2(n654), .ZN(n628) );
  XNOR2_X1 U708 ( .A(KEYINPUT67), .B(n628), .ZN(n629) );
  NOR2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U710 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U711 ( .A1(G61), .A2(n654), .ZN(n633) );
  XNOR2_X1 U712 ( .A(n633), .B(KEYINPUT82), .ZN(n642) );
  NAND2_X1 U713 ( .A1(G73), .A2(n650), .ZN(n634) );
  XNOR2_X1 U714 ( .A(n634), .B(KEYINPUT84), .ZN(n635) );
  XNOR2_X1 U715 ( .A(n635), .B(KEYINPUT2), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G48), .A2(n653), .ZN(n636) );
  NAND2_X1 U717 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U718 ( .A1(G86), .A2(n649), .ZN(n638) );
  XNOR2_X1 U719 ( .A(KEYINPUT83), .B(n638), .ZN(n639) );
  NOR2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G49), .A2(n653), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U725 ( .A1(n654), .A2(n645), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n646), .A2(G87), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(G288) );
  NAND2_X1 U728 ( .A1(G88), .A2(n649), .ZN(n652) );
  NAND2_X1 U729 ( .A1(G75), .A2(n650), .ZN(n651) );
  NAND2_X1 U730 ( .A1(n652), .A2(n651), .ZN(n658) );
  NAND2_X1 U731 ( .A1(G50), .A2(n653), .ZN(n656) );
  NAND2_X1 U732 ( .A1(G62), .A2(n654), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U734 ( .A1(n658), .A2(n657), .ZN(G166) );
  INV_X1 U735 ( .A(G166), .ZN(G303) );
  XOR2_X1 U736 ( .A(G299), .B(G290), .Z(n659) );
  XNOR2_X1 U737 ( .A(n659), .B(G305), .ZN(n662) );
  XOR2_X1 U738 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n660) );
  XNOR2_X1 U739 ( .A(G288), .B(n660), .ZN(n661) );
  XOR2_X1 U740 ( .A(n662), .B(n661), .Z(n664) );
  XOR2_X1 U741 ( .A(G303), .B(n668), .Z(n663) );
  XNOR2_X1 U742 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(n977), .ZN(n911) );
  XOR2_X1 U744 ( .A(n911), .B(n666), .Z(n667) );
  NAND2_X1 U745 ( .A1(G868), .A2(n667), .ZN(n670) );
  OR2_X1 U746 ( .A1(n668), .A2(G868), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G235), .A2(G236), .ZN(n675) );
  XNOR2_X1 U755 ( .A(n675), .B(KEYINPUT87), .ZN(n676) );
  NOR2_X1 U756 ( .A1(G238), .A2(n676), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G57), .A2(n677), .ZN(n833) );
  NAND2_X1 U758 ( .A1(n833), .A2(G567), .ZN(n683) );
  NOR2_X1 U759 ( .A1(G220), .A2(G219), .ZN(n678) );
  XNOR2_X1 U760 ( .A(KEYINPUT22), .B(n678), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n679), .A2(G96), .ZN(n680) );
  NOR2_X1 U762 ( .A1(G218), .A2(n680), .ZN(n681) );
  XOR2_X1 U763 ( .A(KEYINPUT86), .B(n681), .Z(n834) );
  NAND2_X1 U764 ( .A1(n834), .A2(G2106), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n683), .A2(n682), .ZN(n835) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n684) );
  NOR2_X1 U767 ( .A1(n835), .A2(n684), .ZN(n832) );
  NAND2_X1 U768 ( .A1(n832), .A2(G36), .ZN(n685) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(n685), .ZN(G176) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n759) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n758) );
  INV_X1 U772 ( .A(n758), .ZN(n688) );
  AND2_X1 U773 ( .A1(n688), .A2(G1996), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n759), .A2(n686), .ZN(n687) );
  XNOR2_X1 U775 ( .A(n687), .B(KEYINPUT26), .ZN(n690) );
  AND2_X2 U776 ( .A1(n688), .A2(n759), .ZN(n700) );
  NAND2_X1 U777 ( .A1(G1341), .A2(n732), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U779 ( .A(KEYINPUT94), .B(n691), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n692), .A2(n977), .ZN(n693) );
  XNOR2_X1 U781 ( .A(n693), .B(KEYINPUT64), .ZN(n705) );
  NAND2_X1 U782 ( .A1(n705), .A2(n973), .ZN(n698) );
  NAND2_X1 U783 ( .A1(G1348), .A2(n732), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G2067), .A2(n700), .ZN(n694) );
  NAND2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U786 ( .A(KEYINPUT95), .B(n696), .Z(n697) );
  NAND2_X1 U787 ( .A1(n698), .A2(n697), .ZN(n704) );
  NAND2_X1 U788 ( .A1(n700), .A2(G2072), .ZN(n699) );
  XNOR2_X1 U789 ( .A(n699), .B(KEYINPUT27), .ZN(n702) );
  INV_X1 U790 ( .A(G1956), .ZN(n858) );
  NOR2_X1 U791 ( .A1(n858), .A2(n700), .ZN(n701) );
  NOR2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n711) );
  NOR2_X1 U793 ( .A1(n712), .A2(n711), .ZN(n703) );
  XOR2_X1 U794 ( .A(n703), .B(KEYINPUT28), .Z(n710) );
  AND2_X1 U795 ( .A1(n704), .A2(n710), .ZN(n709) );
  NOR2_X1 U796 ( .A1(n973), .A2(n705), .ZN(n707) );
  XNOR2_X1 U797 ( .A(n707), .B(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n716) );
  INV_X1 U799 ( .A(n710), .ZN(n714) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  OR2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U803 ( .A(n717), .B(KEYINPUT29), .ZN(n721) );
  XNOR2_X1 U804 ( .A(G2078), .B(KEYINPUT25), .ZN(n948) );
  NOR2_X1 U805 ( .A1(n732), .A2(n948), .ZN(n719) );
  AND2_X1 U806 ( .A1(n732), .A2(G1961), .ZN(n718) );
  NOR2_X1 U807 ( .A1(n719), .A2(n718), .ZN(n726) );
  AND2_X1 U808 ( .A1(G171), .A2(n726), .ZN(n720) );
  XNOR2_X1 U809 ( .A(n722), .B(KEYINPUT97), .ZN(n731) );
  NAND2_X1 U810 ( .A1(G8), .A2(n732), .ZN(n802) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n802), .ZN(n745) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n732), .ZN(n741) );
  NOR2_X1 U813 ( .A1(n745), .A2(n741), .ZN(n723) );
  NAND2_X1 U814 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U815 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U817 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U818 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U819 ( .A(KEYINPUT31), .B(n729), .Z(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n743) );
  NAND2_X1 U821 ( .A1(n743), .A2(G286), .ZN(n738) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n802), .ZN(n734) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U825 ( .A1(n735), .A2(G303), .ZN(n736) );
  XNOR2_X1 U826 ( .A(n736), .B(KEYINPUT98), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n739), .A2(G8), .ZN(n740) );
  XOR2_X1 U829 ( .A(KEYINPUT32), .B(n740), .Z(n795) );
  NAND2_X1 U830 ( .A1(G8), .A2(n741), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n793) );
  NOR2_X1 U833 ( .A1(n795), .A2(n793), .ZN(n746) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n747) );
  XNOR2_X1 U836 ( .A(n747), .B(KEYINPUT99), .ZN(n749) );
  INV_X1 U837 ( .A(KEYINPUT33), .ZN(n748) );
  AND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n757) );
  INV_X1 U840 ( .A(n802), .ZN(n792) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n991) );
  AND2_X1 U842 ( .A1(n792), .A2(n991), .ZN(n752) );
  NOR2_X1 U843 ( .A1(KEYINPUT33), .A2(n752), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n993), .A2(KEYINPUT33), .ZN(n753) );
  NOR2_X1 U845 ( .A1(n753), .A2(n802), .ZN(n754) );
  NOR2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n756) );
  AND2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n790) );
  XOR2_X1 U848 ( .A(G1981), .B(G305), .Z(n984) );
  NOR2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n824) );
  NAND2_X1 U850 ( .A1(n894), .A2(G104), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G140), .A2(n896), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U853 ( .A(KEYINPUT34), .B(n762), .ZN(n767) );
  NAND2_X1 U854 ( .A1(G128), .A2(n903), .ZN(n764) );
  NAND2_X1 U855 ( .A1(G116), .A2(n900), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U857 ( .A(KEYINPUT35), .B(n765), .Z(n766) );
  NOR2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U859 ( .A(KEYINPUT36), .B(n768), .Z(n884) );
  XOR2_X1 U860 ( .A(G2067), .B(KEYINPUT37), .Z(n821) );
  AND2_X1 U861 ( .A1(n884), .A2(n821), .ZN(n927) );
  NAND2_X1 U862 ( .A1(n824), .A2(n927), .ZN(n819) );
  AND2_X1 U863 ( .A1(n984), .A2(n819), .ZN(n788) );
  NAND2_X1 U864 ( .A1(G129), .A2(n903), .ZN(n770) );
  NAND2_X1 U865 ( .A1(G117), .A2(n900), .ZN(n769) );
  NAND2_X1 U866 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U867 ( .A1(G105), .A2(n894), .ZN(n771) );
  XNOR2_X1 U868 ( .A(n771), .B(KEYINPUT91), .ZN(n772) );
  XNOR2_X1 U869 ( .A(n772), .B(KEYINPUT38), .ZN(n773) );
  NOR2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U871 ( .A(n775), .B(KEYINPUT92), .ZN(n777) );
  NAND2_X1 U872 ( .A1(G141), .A2(n896), .ZN(n776) );
  NAND2_X1 U873 ( .A1(n777), .A2(n776), .ZN(n883) );
  AND2_X1 U874 ( .A1(n883), .A2(G1996), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n894), .A2(G95), .ZN(n779) );
  NAND2_X1 U876 ( .A1(G131), .A2(n896), .ZN(n778) );
  NAND2_X1 U877 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U878 ( .A1(G119), .A2(n903), .ZN(n781) );
  NAND2_X1 U879 ( .A1(G107), .A2(n900), .ZN(n780) );
  NAND2_X1 U880 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U881 ( .A1(n783), .A2(n782), .ZN(n891) );
  INV_X1 U882 ( .A(G1991), .ZN(n864) );
  NOR2_X1 U883 ( .A1(n891), .A2(n864), .ZN(n784) );
  NOR2_X1 U884 ( .A1(n785), .A2(n784), .ZN(n929) );
  INV_X1 U885 ( .A(n824), .ZN(n786) );
  NOR2_X1 U886 ( .A1(n929), .A2(n786), .ZN(n816) );
  XOR2_X1 U887 ( .A(KEYINPUT93), .B(n816), .Z(n808) );
  INV_X1 U888 ( .A(n808), .ZN(n787) );
  AND2_X1 U889 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U890 ( .A1(n790), .A2(n789), .ZN(n810) );
  INV_X1 U891 ( .A(n819), .ZN(n791) );
  OR2_X1 U892 ( .A1(n792), .A2(n791), .ZN(n796) );
  OR2_X1 U893 ( .A1(n793), .A2(n796), .ZN(n794) );
  NOR2_X1 U894 ( .A1(n795), .A2(n794), .ZN(n806) );
  INV_X1 U895 ( .A(n796), .ZN(n799) );
  NAND2_X1 U896 ( .A1(G166), .A2(G8), .ZN(n797) );
  NOR2_X1 U897 ( .A1(G2090), .A2(n797), .ZN(n798) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n800) );
  XOR2_X1 U899 ( .A(n800), .B(KEYINPUT24), .Z(n801) );
  NOR2_X1 U900 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n819), .A2(n803), .ZN(n804) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  OR2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n812) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n981) );
  NAND2_X1 U906 ( .A1(n981), .A2(n824), .ZN(n811) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n827) );
  NOR2_X1 U908 ( .A1(G1996), .A2(n883), .ZN(n935) );
  AND2_X1 U909 ( .A1(n864), .A2(n891), .ZN(n923) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n813) );
  XNOR2_X1 U911 ( .A(KEYINPUT100), .B(n813), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n923), .A2(n814), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U914 ( .A1(n935), .A2(n817), .ZN(n818) );
  XNOR2_X1 U915 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n823) );
  NOR2_X1 U917 ( .A1(n821), .A2(n884), .ZN(n822) );
  XNOR2_X1 U918 ( .A(n822), .B(KEYINPUT101), .ZN(n941) );
  NAND2_X1 U919 ( .A1(n823), .A2(n941), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n828), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U924 ( .A(n829), .ZN(G223) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U926 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n834), .A2(n833), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n835), .ZN(G319) );
  XNOR2_X1 U934 ( .A(G1341), .B(G1348), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n836), .B(G2427), .ZN(n846) );
  XOR2_X1 U936 ( .A(KEYINPUT104), .B(G2430), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2446), .B(G2451), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U939 ( .A(KEYINPUT102), .B(G2438), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2435), .B(G2454), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U943 ( .A(KEYINPUT103), .B(G2443), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  NAND2_X1 U946 ( .A1(n847), .A2(G14), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n848), .B(KEYINPUT105), .ZN(G401) );
  XNOR2_X1 U948 ( .A(n849), .B(G2096), .ZN(n851) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U951 ( .A(KEYINPUT43), .B(G2090), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U954 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U955 ( .A(G2078), .B(G2084), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(G227) );
  XOR2_X1 U957 ( .A(G1976), .B(G1971), .Z(n860) );
  XOR2_X1 U958 ( .A(G1986), .B(n858), .Z(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U960 ( .A(n861), .B(KEYINPUT41), .Z(n863) );
  XNOR2_X1 U961 ( .A(G1966), .B(G1981), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n863), .B(n862), .ZN(n868) );
  XOR2_X1 U963 ( .A(G2474), .B(G1961), .Z(n866) );
  XOR2_X1 U964 ( .A(G1996), .B(n864), .Z(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(G229) );
  NAND2_X1 U967 ( .A1(n903), .A2(G124), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G112), .A2(n900), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n894), .A2(G100), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G136), .A2(n896), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U974 ( .A1(n875), .A2(n874), .ZN(G162) );
  NAND2_X1 U975 ( .A1(n894), .A2(G103), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G139), .A2(n896), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G127), .A2(n903), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G115), .A2(n900), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n930) );
  XOR2_X1 U983 ( .A(n922), .B(n930), .Z(n886) );
  XOR2_X1 U984 ( .A(n884), .B(n883), .Z(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT108), .Z(n888) );
  XNOR2_X1 U987 ( .A(G162), .B(KEYINPUT46), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n890), .B(n889), .Z(n893) );
  XNOR2_X1 U990 ( .A(G160), .B(n891), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n893), .B(n892), .ZN(n909) );
  NAND2_X1 U992 ( .A1(n894), .A2(G106), .ZN(n895) );
  XOR2_X1 U993 ( .A(KEYINPUT107), .B(n895), .Z(n898) );
  NAND2_X1 U994 ( .A1(G142), .A2(n896), .ZN(n897) );
  NAND2_X1 U995 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U996 ( .A(n899), .B(KEYINPUT45), .ZN(n902) );
  NAND2_X1 U997 ( .A1(G118), .A2(n900), .ZN(n901) );
  NAND2_X1 U998 ( .A1(n902), .A2(n901), .ZN(n906) );
  NAND2_X1 U999 ( .A1(n903), .A2(G130), .ZN(n904) );
  XOR2_X1 U1000 ( .A(KEYINPUT106), .B(n904), .Z(n905) );
  NOR2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(G164), .B(n907), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1005 ( .A(G286), .B(n911), .ZN(n913) );
  XOR2_X1 U1006 ( .A(G301), .B(n973), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(KEYINPUT109), .B(KEYINPUT49), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n919) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(n917), .B(KEYINPUT110), .ZN(n918) );
  NAND2_X1 U1014 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n920), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n921), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1019 ( .A(KEYINPUT111), .B(KEYINPUT52), .Z(n944) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n925) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1022 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1024 ( .A1(n929), .A2(n928), .ZN(n940) );
  XOR2_X1 U1025 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(KEYINPUT50), .B(n933), .ZN(n938) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(n944), .B(n943), .ZN(n945) );
  NOR2_X1 U1036 ( .A1(KEYINPUT55), .A2(n945), .ZN(n946) );
  XOR2_X1 U1037 ( .A(KEYINPUT112), .B(n946), .Z(n947) );
  NAND2_X1 U1038 ( .A1(G29), .A2(n947), .ZN(n1033) );
  XOR2_X1 U1039 ( .A(G2090), .B(G35), .Z(n963) );
  XNOR2_X1 U1040 ( .A(G27), .B(n948), .ZN(n952) );
  XNOR2_X1 U1041 ( .A(G2067), .B(G26), .ZN(n950) );
  XNOR2_X1 U1042 ( .A(G2072), .B(G33), .ZN(n949) );
  NOR2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(KEYINPUT114), .B(G1996), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G32), .B(n953), .ZN(n954) );
  NOR2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n959) );
  XOR2_X1 U1048 ( .A(G1991), .B(G25), .Z(n956) );
  NAND2_X1 U1049 ( .A1(n956), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT113), .ZN(n958) );
  NAND2_X1 U1051 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1052 ( .A(KEYINPUT115), .B(n960), .Z(n961) );
  XNOR2_X1 U1053 ( .A(n961), .B(KEYINPUT53), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(n963), .A2(n962), .ZN(n968) );
  XOR2_X1 U1055 ( .A(G34), .B(KEYINPUT117), .Z(n965) );
  XNOR2_X1 U1056 ( .A(G2084), .B(KEYINPUT54), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n966), .B(KEYINPUT116), .ZN(n967) );
  NOR2_X1 U1059 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1060 ( .A(KEYINPUT55), .B(n969), .ZN(n971) );
  INV_X1 U1061 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(n972), .A2(G11), .ZN(n1031) );
  INV_X1 U1064 ( .A(G16), .ZN(n1027) );
  XOR2_X1 U1065 ( .A(n1027), .B(KEYINPUT56), .Z(n999) );
  XNOR2_X1 U1066 ( .A(n973), .B(G1348), .ZN(n975) );
  XOR2_X1 U1067 ( .A(G301), .B(G1961), .Z(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT119), .B(n976), .ZN(n983) );
  XOR2_X1 U1070 ( .A(n977), .B(G1341), .Z(n979) );
  XOR2_X1 U1071 ( .A(G299), .B(G1956), .Z(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n989) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1077 ( .A(KEYINPUT118), .B(n986), .Z(n987) );
  XNOR2_X1 U1078 ( .A(KEYINPUT57), .B(n987), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n997) );
  XOR2_X1 U1080 ( .A(G303), .B(G1971), .Z(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(KEYINPUT120), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1084 ( .A(KEYINPUT121), .B(n995), .Z(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1029) );
  XOR2_X1 U1087 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n1006) );
  XNOR2_X1 U1088 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1004) );
  XOR2_X1 U1091 ( .A(G1986), .B(KEYINPUT126), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(G24), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1006), .B(n1005), .ZN(n1024) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1981), .B(G6), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(KEYINPUT122), .B(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(G1956), .B(G20), .Z(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  XNOR2_X1 U1101 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(n1012), .B(G4), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(n1013), .B(G1348), .ZN(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1016), .Z(n1018) );
  XNOR2_X1 U1106 ( .A(G1966), .B(G21), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1108 ( .A(KEYINPUT124), .B(n1019), .Z(n1021) );
  XNOR2_X1 U1109 ( .A(G1961), .B(G5), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(n1022), .B(KEYINPUT125), .ZN(n1023) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1034), .ZN(G150) );
  INV_X1 U1119 ( .A(G150), .ZN(G311) );
endmodule

