

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597;

  NOR2_X1 U323 ( .A1(n477), .A2(n595), .ZN(n480) );
  XOR2_X1 U324 ( .A(n330), .B(n329), .Z(n580) );
  AND2_X1 U325 ( .A1(n370), .A2(n369), .ZN(n372) );
  NOR2_X1 U326 ( .A1(n475), .A2(n474), .ZN(n506) );
  XNOR2_X1 U327 ( .A(n489), .B(n488), .ZN(n548) );
  AND2_X1 U328 ( .A1(n566), .A2(n580), .ZN(n332) );
  INV_X1 U329 ( .A(KEYINPUT86), .ZN(n439) );
  XNOR2_X1 U330 ( .A(n440), .B(n439), .ZN(n441) );
  INV_X1 U331 ( .A(KEYINPUT31), .ZN(n295) );
  XNOR2_X1 U332 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U333 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U334 ( .A(n448), .B(n447), .ZN(n449) );
  INV_X1 U335 ( .A(KEYINPUT37), .ZN(n478) );
  XNOR2_X1 U336 ( .A(n450), .B(n449), .ZN(n454) );
  XNOR2_X1 U337 ( .A(n478), .B(KEYINPUT102), .ZN(n479) );
  INV_X1 U338 ( .A(KEYINPUT116), .ZN(n418) );
  XNOR2_X1 U339 ( .A(n480), .B(n479), .ZN(n487) );
  XNOR2_X1 U340 ( .A(n419), .B(n418), .ZN(n560) );
  XNOR2_X1 U341 ( .A(n392), .B(n391), .ZN(n393) );
  AND2_X1 U342 ( .A1(n487), .A2(n507), .ZN(n483) );
  NOR2_X1 U343 ( .A1(n537), .A2(n499), .ZN(n575) );
  XNOR2_X1 U344 ( .A(n394), .B(n393), .ZN(n546) );
  XNOR2_X1 U345 ( .A(n500), .B(G176GAT), .ZN(n501) );
  XNOR2_X1 U346 ( .A(n458), .B(G120GAT), .ZN(n459) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n484) );
  XNOR2_X1 U348 ( .A(n502), .B(n501), .ZN(G1349GAT) );
  XNOR2_X1 U349 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  XNOR2_X1 U350 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n291) );
  XNOR2_X1 U351 ( .A(n291), .B(KEYINPUT72), .ZN(n339) );
  XOR2_X1 U352 ( .A(G85GAT), .B(G99GAT), .Z(n353) );
  XNOR2_X1 U353 ( .A(n339), .B(n353), .ZN(n292) );
  INV_X1 U354 ( .A(n292), .ZN(n294) );
  NAND2_X1 U355 ( .A1(G230GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U356 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U357 ( .A(G120GAT), .B(G71GAT), .Z(n428) );
  XNOR2_X1 U358 ( .A(n428), .B(KEYINPUT32), .ZN(n296) );
  XNOR2_X1 U359 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U360 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n300) );
  XNOR2_X1 U361 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n299) );
  XNOR2_X1 U362 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U363 ( .A(n302), .B(n301), .Z(n308) );
  XOR2_X1 U364 ( .A(KEYINPUT73), .B(G78GAT), .Z(n304) );
  XNOR2_X1 U365 ( .A(G148GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U366 ( .A(n304), .B(n303), .ZN(n442) );
  XOR2_X1 U367 ( .A(G176GAT), .B(G204GAT), .Z(n306) );
  XNOR2_X1 U368 ( .A(G92GAT), .B(G64GAT), .ZN(n305) );
  XNOR2_X1 U369 ( .A(n306), .B(n305), .ZN(n384) );
  XNOR2_X1 U370 ( .A(n442), .B(n384), .ZN(n307) );
  XNOR2_X1 U371 ( .A(n308), .B(n307), .ZN(n584) );
  NAND2_X1 U372 ( .A1(n584), .A2(KEYINPUT64), .ZN(n312) );
  INV_X1 U373 ( .A(n584), .ZN(n310) );
  INV_X1 U374 ( .A(KEYINPUT64), .ZN(n309) );
  NAND2_X1 U375 ( .A1(n310), .A2(n309), .ZN(n311) );
  NAND2_X1 U376 ( .A1(n312), .A2(n311), .ZN(n313) );
  XOR2_X2 U377 ( .A(n313), .B(KEYINPUT41), .Z(n566) );
  XOR2_X1 U378 ( .A(KEYINPUT71), .B(G197GAT), .Z(n315) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(G141GAT), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n330) );
  XOR2_X1 U381 ( .A(KEYINPUT70), .B(KEYINPUT69), .Z(n317) );
  XNOR2_X1 U382 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n316) );
  XNOR2_X1 U383 ( .A(n317), .B(n316), .ZN(n323) );
  XOR2_X1 U384 ( .A(G43GAT), .B(KEYINPUT7), .Z(n319) );
  XNOR2_X1 U385 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n318) );
  XNOR2_X1 U386 ( .A(n319), .B(n318), .ZN(n352) );
  XOR2_X1 U387 ( .A(n352), .B(KEYINPUT29), .Z(n321) );
  NAND2_X1 U388 ( .A1(G229GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U389 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U390 ( .A(n323), .B(n322), .ZN(n328) );
  XOR2_X1 U391 ( .A(G8GAT), .B(G169GAT), .Z(n392) );
  XNOR2_X1 U392 ( .A(G1GAT), .B(G15GAT), .ZN(n324) );
  XNOR2_X1 U393 ( .A(n324), .B(G22GAT), .ZN(n336) );
  XOR2_X1 U394 ( .A(n392), .B(n336), .Z(n326) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(G50GAT), .ZN(n325) );
  XNOR2_X1 U396 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U397 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U398 ( .A(KEYINPUT46), .B(KEYINPUT114), .ZN(n331) );
  XNOR2_X1 U399 ( .A(n332), .B(n331), .ZN(n333) );
  OR2_X1 U400 ( .A1(n333), .A2(KEYINPUT113), .ZN(n335) );
  NAND2_X1 U401 ( .A1(KEYINPUT113), .A2(n333), .ZN(n334) );
  NAND2_X1 U402 ( .A1(n335), .A2(n334), .ZN(n370) );
  XOR2_X1 U403 ( .A(G183GAT), .B(KEYINPUT78), .Z(n388) );
  XOR2_X1 U404 ( .A(n336), .B(n388), .Z(n338) );
  XNOR2_X1 U405 ( .A(G127GAT), .B(G71GAT), .ZN(n337) );
  XNOR2_X1 U406 ( .A(n338), .B(n337), .ZN(n343) );
  XOR2_X1 U407 ( .A(n339), .B(KEYINPUT79), .Z(n341) );
  NAND2_X1 U408 ( .A1(G231GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U410 ( .A(n343), .B(n342), .Z(n351) );
  XOR2_X1 U411 ( .A(G8GAT), .B(G211GAT), .Z(n345) );
  XNOR2_X1 U412 ( .A(G155GAT), .B(G78GAT), .ZN(n344) );
  XNOR2_X1 U413 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U414 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n347) );
  XNOR2_X1 U415 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n346) );
  XNOR2_X1 U416 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U417 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U418 ( .A(n351), .B(n350), .Z(n503) );
  XOR2_X1 U419 ( .A(G162GAT), .B(G50GAT), .Z(n444) );
  XNOR2_X1 U420 ( .A(n352), .B(n444), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n359) );
  XNOR2_X1 U422 ( .A(G36GAT), .B(KEYINPUT77), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n355), .B(G190GAT), .ZN(n381) );
  XOR2_X1 U424 ( .A(n381), .B(G92GAT), .Z(n357) );
  NAND2_X1 U425 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U427 ( .A(n359), .B(n358), .Z(n367) );
  XOR2_X1 U428 ( .A(KEYINPUT11), .B(G106GAT), .Z(n361) );
  XNOR2_X1 U429 ( .A(G134GAT), .B(G218GAT), .ZN(n360) );
  XNOR2_X1 U430 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U431 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n363) );
  XNOR2_X1 U432 ( .A(KEYINPUT65), .B(KEYINPUT10), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U435 ( .A(n367), .B(n366), .Z(n574) );
  INV_X1 U436 ( .A(n574), .ZN(n368) );
  AND2_X1 U437 ( .A1(n503), .A2(n368), .ZN(n369) );
  XNOR2_X1 U438 ( .A(KEYINPUT115), .B(KEYINPUT47), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n377) );
  XOR2_X1 U440 ( .A(KEYINPUT36), .B(n574), .Z(n595) );
  NOR2_X1 U441 ( .A1(n595), .A2(n503), .ZN(n373) );
  XNOR2_X1 U442 ( .A(n373), .B(KEYINPUT45), .ZN(n374) );
  INV_X1 U443 ( .A(n580), .ZN(n481) );
  NAND2_X1 U444 ( .A1(n374), .A2(n481), .ZN(n375) );
  NOR2_X1 U445 ( .A1(n584), .A2(n375), .ZN(n376) );
  NOR2_X1 U446 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U447 ( .A(n378), .B(KEYINPUT48), .ZN(n494) );
  XOR2_X1 U448 ( .A(G197GAT), .B(KEYINPUT21), .Z(n380) );
  XNOR2_X1 U449 ( .A(G218GAT), .B(G211GAT), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n380), .B(n379), .ZN(n451) );
  XNOR2_X1 U451 ( .A(n381), .B(n451), .ZN(n386) );
  XNOR2_X1 U452 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n382), .B(KEYINPUT18), .ZN(n429) );
  INV_X1 U454 ( .A(n429), .ZN(n383) );
  XNOR2_X1 U455 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U456 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U457 ( .A(n387), .B(KEYINPUT93), .ZN(n390) );
  XOR2_X1 U458 ( .A(n388), .B(KEYINPUT92), .Z(n389) );
  XNOR2_X1 U459 ( .A(n390), .B(n389), .ZN(n394) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XOR2_X1 U461 ( .A(n546), .B(KEYINPUT27), .Z(n466) );
  XOR2_X1 U462 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n396) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n396), .B(n395), .ZN(n405) );
  XOR2_X1 U465 ( .A(KEYINPUT90), .B(KEYINPUT88), .Z(n403) );
  XOR2_X1 U466 ( .A(KEYINPUT0), .B(G134GAT), .Z(n398) );
  XNOR2_X1 U467 ( .A(G127GAT), .B(G113GAT), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U469 ( .A(KEYINPUT80), .B(n399), .Z(n433) );
  XOR2_X1 U470 ( .A(G141GAT), .B(G155GAT), .Z(n401) );
  XNOR2_X1 U471 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n400) );
  XNOR2_X1 U472 ( .A(n401), .B(n400), .ZN(n452) );
  XNOR2_X1 U473 ( .A(n433), .B(n452), .ZN(n402) );
  XNOR2_X1 U474 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U475 ( .A(n405), .B(n404), .ZN(n417) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n411) );
  XOR2_X1 U477 ( .A(G57GAT), .B(G148GAT), .Z(n407) );
  XNOR2_X1 U478 ( .A(G85GAT), .B(G120GAT), .ZN(n406) );
  XNOR2_X1 U479 ( .A(n407), .B(n406), .ZN(n409) );
  XOR2_X1 U480 ( .A(G29GAT), .B(G162GAT), .Z(n408) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U482 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U483 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n413) );
  XNOR2_X1 U484 ( .A(KEYINPUT87), .B(KEYINPUT1), .ZN(n412) );
  XNOR2_X1 U485 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U486 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U487 ( .A(n417), .B(n416), .Z(n544) );
  INV_X1 U488 ( .A(n544), .ZN(n531) );
  OR2_X1 U489 ( .A1(n466), .A2(n531), .ZN(n470) );
  NOR2_X1 U490 ( .A1(n494), .A2(n470), .ZN(n419) );
  XOR2_X1 U491 ( .A(G169GAT), .B(G176GAT), .Z(n421) );
  XNOR2_X1 U492 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n420) );
  XNOR2_X1 U493 ( .A(n421), .B(n420), .ZN(n437) );
  XOR2_X1 U494 ( .A(G183GAT), .B(G99GAT), .Z(n423) );
  XNOR2_X1 U495 ( .A(G190GAT), .B(G43GAT), .ZN(n422) );
  XNOR2_X1 U496 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U497 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n425) );
  XNOR2_X1 U498 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n424) );
  XNOR2_X1 U499 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U500 ( .A(n427), .B(n426), .Z(n435) );
  XOR2_X1 U501 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U502 ( .A1(G227GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U503 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U504 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U505 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U506 ( .A(n437), .B(n436), .Z(n549) );
  INV_X1 U507 ( .A(n549), .ZN(n537) );
  NOR2_X1 U508 ( .A1(n560), .A2(n537), .ZN(n438) );
  XNOR2_X1 U509 ( .A(n438), .B(KEYINPUT117), .ZN(n457) );
  INV_X1 U510 ( .A(KEYINPUT28), .ZN(n456) );
  NAND2_X1 U511 ( .A1(G228GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U512 ( .A(n443), .B(KEYINPUT22), .ZN(n450) );
  XOR2_X1 U513 ( .A(n444), .B(KEYINPUT24), .Z(n448) );
  XOR2_X1 U514 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n446) );
  XNOR2_X1 U515 ( .A(G22GAT), .B(G204GAT), .ZN(n445) );
  XOR2_X1 U516 ( .A(n446), .B(n445), .Z(n447) );
  XNOR2_X1 U517 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(n497) );
  XNOR2_X1 U519 ( .A(n497), .B(KEYINPUT67), .ZN(n455) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(n515) );
  NOR2_X1 U521 ( .A1(n457), .A2(n515), .ZN(n557) );
  NAND2_X1 U522 ( .A1(n557), .A2(n566), .ZN(n460) );
  XOR2_X1 U523 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n458) );
  XNOR2_X1 U524 ( .A(n460), .B(n459), .ZN(G1341GAT) );
  INV_X1 U525 ( .A(n503), .ZN(n588) );
  INV_X1 U526 ( .A(n546), .ZN(n534) );
  NOR2_X1 U527 ( .A1(n534), .A2(n537), .ZN(n461) );
  XNOR2_X1 U528 ( .A(n461), .B(KEYINPUT96), .ZN(n462) );
  NOR2_X1 U529 ( .A1(n497), .A2(n462), .ZN(n463) );
  XNOR2_X1 U530 ( .A(n463), .B(KEYINPUT25), .ZN(n464) );
  XNOR2_X1 U531 ( .A(n464), .B(KEYINPUT97), .ZN(n468) );
  NAND2_X1 U532 ( .A1(n537), .A2(n497), .ZN(n465) );
  XNOR2_X1 U533 ( .A(n465), .B(KEYINPUT26), .ZN(n579) );
  NOR2_X1 U534 ( .A1(n579), .A2(n466), .ZN(n467) );
  NOR2_X1 U535 ( .A1(n468), .A2(n467), .ZN(n469) );
  NOR2_X1 U536 ( .A1(n544), .A2(n469), .ZN(n475) );
  NOR2_X1 U537 ( .A1(n470), .A2(n515), .ZN(n471) );
  XNOR2_X1 U538 ( .A(KEYINPUT94), .B(n471), .ZN(n472) );
  AND2_X1 U539 ( .A1(n472), .A2(n537), .ZN(n473) );
  XOR2_X1 U540 ( .A(n473), .B(KEYINPUT95), .Z(n474) );
  NOR2_X1 U541 ( .A1(n588), .A2(n506), .ZN(n476) );
  XNOR2_X1 U542 ( .A(n476), .B(KEYINPUT101), .ZN(n477) );
  NOR2_X1 U543 ( .A1(n584), .A2(n481), .ZN(n507) );
  INV_X1 U544 ( .A(KEYINPUT38), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n525) );
  NOR2_X1 U546 ( .A1(n531), .A2(n525), .ZN(n485) );
  INV_X1 U547 ( .A(KEYINPUT110), .ZN(n489) );
  INV_X1 U548 ( .A(n566), .ZN(n486) );
  NOR2_X1 U549 ( .A1(n580), .A2(n486), .ZN(n530) );
  NAND2_X1 U550 ( .A1(n530), .A2(n487), .ZN(n488) );
  NAND2_X1 U551 ( .A1(n548), .A2(n515), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n491) );
  INV_X1 U553 ( .A(G106GAT), .ZN(n490) );
  XNOR2_X1 U554 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U555 ( .A(n493), .B(n492), .ZN(G1339GAT) );
  NOR2_X1 U556 ( .A1(n534), .A2(n494), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(KEYINPUT54), .ZN(n496) );
  NAND2_X1 U558 ( .A1(n496), .A2(n531), .ZN(n578) );
  NOR2_X1 U559 ( .A1(n497), .A2(n578), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(KEYINPUT55), .ZN(n499) );
  NAND2_X1 U561 ( .A1(n575), .A2(n566), .ZN(n502) );
  XOR2_X1 U562 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n500) );
  NOR2_X1 U563 ( .A1(n574), .A2(n503), .ZN(n504) );
  XOR2_X1 U564 ( .A(KEYINPUT16), .B(n504), .Z(n505) );
  NOR2_X1 U565 ( .A1(n506), .A2(n505), .ZN(n529) );
  NAND2_X1 U566 ( .A1(n507), .A2(n529), .ZN(n516) );
  NOR2_X1 U567 ( .A1(n531), .A2(n516), .ZN(n508) );
  XOR2_X1 U568 ( .A(KEYINPUT34), .B(n508), .Z(n509) );
  XNOR2_X1 U569 ( .A(G1GAT), .B(n509), .ZN(G1324GAT) );
  NOR2_X1 U570 ( .A1(n534), .A2(n516), .ZN(n510) );
  XOR2_X1 U571 ( .A(G8GAT), .B(n510), .Z(G1325GAT) );
  NOR2_X1 U572 ( .A1(n516), .A2(n537), .ZN(n514) );
  XOR2_X1 U573 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n512) );
  XNOR2_X1 U574 ( .A(G15GAT), .B(KEYINPUT99), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(n514), .B(n513), .ZN(G1326GAT) );
  INV_X1 U577 ( .A(n515), .ZN(n541) );
  NOR2_X1 U578 ( .A1(n541), .A2(n516), .ZN(n517) );
  XOR2_X1 U579 ( .A(KEYINPUT100), .B(n517), .Z(n518) );
  XNOR2_X1 U580 ( .A(G22GAT), .B(n518), .ZN(G1327GAT) );
  XNOR2_X1 U581 ( .A(G36GAT), .B(KEYINPUT103), .ZN(n520) );
  NOR2_X1 U582 ( .A1(n534), .A2(n525), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1329GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n522) );
  XNOR2_X1 U585 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n524) );
  NOR2_X1 U587 ( .A1(n525), .A2(n537), .ZN(n523) );
  XOR2_X1 U588 ( .A(n524), .B(n523), .Z(G1330GAT) );
  NOR2_X1 U589 ( .A1(n541), .A2(n525), .ZN(n526) );
  XOR2_X1 U590 ( .A(G50GAT), .B(n526), .Z(G1331GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n528) );
  XNOR2_X1 U592 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n540) );
  NOR2_X1 U595 ( .A1(n531), .A2(n540), .ZN(n532) );
  XOR2_X1 U596 ( .A(n533), .B(n532), .Z(G1332GAT) );
  NOR2_X1 U597 ( .A1(n534), .A2(n540), .ZN(n535) );
  XOR2_X1 U598 ( .A(KEYINPUT108), .B(n535), .Z(n536) );
  XNOR2_X1 U599 ( .A(G64GAT), .B(n536), .ZN(G1333GAT) );
  NOR2_X1 U600 ( .A1(n537), .A2(n540), .ZN(n539) );
  XNOR2_X1 U601 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n539), .B(n538), .ZN(G1334GAT) );
  NOR2_X1 U603 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U604 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(G1335GAT) );
  NAND2_X1 U606 ( .A1(n548), .A2(n544), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n545), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U608 ( .A1(n546), .A2(n548), .ZN(n547) );
  XNOR2_X1 U609 ( .A(n547), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U610 ( .A(G99GAT), .B(KEYINPUT111), .Z(n551) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n551), .B(n550), .ZN(G1338GAT) );
  NAND2_X1 U613 ( .A1(n580), .A2(n557), .ZN(n552) );
  XNOR2_X1 U614 ( .A(G113GAT), .B(n552), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(KEYINPUT50), .Z(n554) );
  NAND2_X1 U616 ( .A1(n557), .A2(n588), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n554), .B(n553), .ZN(n556) );
  XNOR2_X1 U618 ( .A(G127GAT), .B(KEYINPUT119), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(G1342GAT) );
  XOR2_X1 U620 ( .A(G134GAT), .B(KEYINPUT51), .Z(n559) );
  NAND2_X1 U621 ( .A1(n557), .A2(n574), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(G1343GAT) );
  XOR2_X1 U623 ( .A(G141GAT), .B(KEYINPUT121), .Z(n562) );
  NOR2_X1 U624 ( .A1(n579), .A2(n560), .ZN(n570) );
  NAND2_X1 U625 ( .A1(n570), .A2(n580), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n562), .B(n561), .ZN(G1344GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U630 ( .A(KEYINPUT52), .B(n565), .Z(n568) );
  NAND2_X1 U631 ( .A1(n570), .A2(n566), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n588), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U637 ( .A1(n580), .A2(n575), .ZN(n572) );
  XNOR2_X1 U638 ( .A(G169GAT), .B(n572), .ZN(G1348GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n588), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1351GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n582) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n593) );
  NAND2_X1 U646 ( .A1(n593), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U650 ( .A1(n593), .A2(n584), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n587), .ZN(G1353GAT) );
  XOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT125), .Z(n590) );
  NAND2_X1 U654 ( .A1(n593), .A2(n588), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n592) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n592), .B(n591), .ZN(n597) );
  INV_X1 U659 ( .A(n593), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U661 ( .A(n597), .B(n596), .Z(G1355GAT) );
endmodule

