//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n547, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g041(.A1(new_n466), .A2(KEYINPUT64), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(KEYINPUT64), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT3), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n463), .A2(KEYINPUT65), .A3(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n479), .A2(new_n462), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n475), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n485), .A2(G124), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n476), .A2(new_n478), .A3(G138), .A4(new_n462), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n463), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n462), .B2(G114), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G102), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(new_n462), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n498), .A2(new_n500), .A3(G2104), .A4(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n476), .A2(new_n478), .A3(G126), .A4(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n496), .A2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n513), .A2(G88), .B1(G62), .B2(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n510), .A2(new_n512), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n515), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G51), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n513), .A2(G89), .A3(new_n518), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n526), .A2(KEYINPUT68), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g104(.A(KEYINPUT68), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n522), .B(new_n525), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G168));
  NOR2_X1   g107(.A1(new_n523), .A2(new_n519), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G90), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n524), .A2(G52), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n511), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n533), .A2(G81), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n524), .A2(G43), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n511), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  AND3_X1   g121(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G36), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n547), .A2(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n513), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n524), .A2(new_n555), .A3(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n533), .A2(G91), .ZN(new_n558));
  OR2_X1    g133(.A1(KEYINPUT69), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(KEYINPUT69), .A2(G65), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n518), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n511), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n557), .A2(new_n558), .A3(new_n564), .ZN(G299));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n531), .B(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n524), .A2(G49), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n533), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n513), .A2(G48), .B1(G73), .B2(G651), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n515), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n513), .A2(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(G61), .A2(G651), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n519), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n511), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT71), .Z(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(G85), .B2(new_n533), .ZN(new_n584));
  XOR2_X1   g159(.A(KEYINPUT72), .B(G47), .Z(new_n585));
  NAND2_X1  g160(.A1(new_n524), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n513), .A2(new_n518), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n592), .A2(new_n593), .B1(G54), .B2(new_n524), .ZN(new_n594));
  NOR2_X1   g169(.A1(KEYINPUT74), .A2(G66), .ZN(new_n595));
  AND2_X1   g170(.A1(KEYINPUT74), .A2(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n518), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT73), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(KEYINPUT75), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(KEYINPUT75), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n588), .B1(new_n606), .B2(G868), .ZN(G284));
  XNOR2_X1  g182(.A(G284), .B(KEYINPUT76), .ZN(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n567), .B2(new_n609), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n567), .B2(new_n609), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT77), .ZN(G148));
  INV_X1    g190(.A(new_n605), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n613), .B1(new_n616), .B2(new_n603), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n483), .A2(G135), .ZN(new_n621));
  OR2_X1    g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n475), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n485), .A2(G123), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n628));
  NOR3_X1   g203(.A1(new_n477), .A2(new_n475), .A3(G2105), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT13), .B(G2100), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n627), .A2(new_n632), .ZN(G156));
  NOR2_X1   g208(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  AOI21_X1  g213(.A(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(KEYINPUT79), .B2(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n641), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  OAI21_X1  g232(.A(KEYINPUT17), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n657), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n659), .A2(new_n655), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n654), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n662), .C1(new_n660), .C2(new_n654), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(new_n662), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n668), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  AOI22_X1  g249(.A1(new_n672), .A2(KEYINPUT20), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n674), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n668), .A3(new_n671), .ZN(new_n677));
  OAI211_X1 g252(.A(new_n675), .B(new_n677), .C1(KEYINPUT20), .C2(new_n672), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT87), .ZN(new_n679));
  XOR2_X1   g254(.A(G1991), .B(G1996), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n681), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G24), .ZN(new_n690));
  INV_X1    g265(.A(G290), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G1986), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n689), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n689), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1971), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT32), .B(G1981), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n689), .A2(G6), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n579), .B2(new_n689), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n696), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(KEYINPUT90), .B1(G16), .B2(G23), .ZN(new_n702));
  OR3_X1    g277(.A1(KEYINPUT90), .A2(G16), .A3(G23), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n702), .B(new_n703), .C1(G288), .C2(new_n689), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n701), .B(new_n706), .C1(new_n697), .C2(new_n700), .ZN(new_n707));
  AOI211_X1 g282(.A(KEYINPUT91), .B(new_n693), .C1(new_n707), .C2(KEYINPUT34), .ZN(new_n708));
  INV_X1    g283(.A(G25), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT88), .B1(new_n709), .B2(G29), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n709), .A2(KEYINPUT88), .A3(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n483), .A2(G131), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(G107), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n475), .B1(new_n714), .B2(G2105), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n485), .A2(G119), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n710), .B(new_n711), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT35), .B(G1991), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n708), .B(new_n722), .C1(KEYINPUT34), .C2(new_n707), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n719), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT29), .B(G2090), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n723), .A2(new_n724), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n689), .A2(G21), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G168), .B2(new_n689), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1966), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n689), .A2(G20), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G299), .B2(G16), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G1956), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n719), .A2(G27), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G164), .B2(new_n719), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2078), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n545), .A2(new_n689), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n689), .B2(G19), .ZN(new_n743));
  INV_X1    g318(.A(G1341), .ZN(new_n744));
  NOR2_X1   g319(.A1(G5), .A2(G16), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G171), .B2(G16), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n743), .A2(new_n744), .B1(G1961), .B2(new_n746), .ZN(new_n747));
  NOR4_X1   g322(.A1(new_n733), .A2(new_n738), .A3(new_n741), .A4(new_n747), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n743), .A2(new_n744), .B1(G1961), .B2(new_n746), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G11), .ZN(new_n750));
  AND2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NOR2_X1   g326(.A1(KEYINPUT24), .A2(G34), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n751), .A2(new_n752), .A3(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n472), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2084), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n626), .A2(G29), .ZN(new_n757));
  AND2_X1   g332(.A1(KEYINPUT30), .A2(G28), .ZN(new_n758));
  NOR2_X1   g333(.A1(KEYINPUT30), .A2(G28), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n719), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G32), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n483), .A2(G141), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT26), .Z(new_n765));
  NOR2_X1   g340(.A1(new_n475), .A2(G2105), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n485), .A2(G129), .B1(G105), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n763), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n762), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT27), .B(G1996), .Z(new_n771));
  AOI21_X1  g346(.A(new_n761), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n749), .A2(new_n750), .A3(new_n756), .A4(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n719), .A2(G33), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n483), .A2(G139), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT94), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2105), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n766), .A2(G103), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT25), .Z(new_n781));
  NAND3_X1  g356(.A1(new_n776), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n774), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT96), .B(G2072), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n754), .A2(new_n755), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n783), .A2(new_n784), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n770), .B2(new_n771), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n773), .A2(new_n785), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n748), .A2(new_n790), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n719), .A2(G26), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n485), .A2(G128), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n462), .A2(G116), .ZN(new_n794));
  OR3_X1    g369(.A1(KEYINPUT92), .A2(G104), .A3(G2105), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT92), .B1(G104), .B2(G2105), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n795), .A2(G2104), .A3(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n793), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G140), .B2(new_n483), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT93), .Z(new_n800));
  AOI21_X1  g375(.A(new_n792), .B1(new_n800), .B2(G29), .ZN(new_n801));
  MUX2_X1   g376(.A(new_n792), .B(new_n801), .S(KEYINPUT28), .Z(new_n802));
  INV_X1    g377(.A(G2067), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NOR2_X1   g380(.A1(G4), .A2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n606), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1348), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n791), .A2(new_n804), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n725), .A2(new_n729), .A3(new_n730), .A4(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  AOI22_X1  g386(.A1(G55), .A2(new_n524), .B1(new_n533), .B2(G93), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT99), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G651), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n606), .A2(G559), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n816), .B(new_n544), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT39), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n818), .B1(new_n823), .B2(G860), .ZN(G145));
  XNOR2_X1  g399(.A(new_n800), .B(new_n768), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n782), .A2(KEYINPUT102), .A3(new_n717), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n503), .A2(KEYINPUT101), .A3(new_n504), .ZN(new_n828));
  AOI21_X1  g403(.A(KEYINPUT101), .B1(new_n503), .B2(new_n504), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n494), .B(new_n495), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n717), .B1(new_n782), .B2(KEYINPUT102), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n827), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n505), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n503), .A2(KEYINPUT101), .A3(new_n504), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n496), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n782), .A2(KEYINPUT102), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n718), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n838), .B2(new_n826), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n825), .B1(new_n832), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n825), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n836), .A3(new_n826), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n830), .B1(new_n827), .B2(new_n831), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n485), .A2(G130), .ZN(new_n846));
  NOR2_X1   g421(.A1(G106), .A2(G2105), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n848));
  INV_X1    g423(.A(G142), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n846), .B1(new_n847), .B2(new_n848), .C1(new_n482), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n630), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n840), .A2(new_n851), .A3(new_n844), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n490), .B(KEYINPUT100), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n472), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n626), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT103), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT103), .A4(new_n857), .ZN(new_n861));
  AOI21_X1  g436(.A(G37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n853), .A2(new_n854), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(new_n857), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n867));
  INV_X1    g442(.A(new_n821), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n617), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n821), .B1(new_n606), .B2(new_n613), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n563), .B1(new_n554), .B2(new_n556), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n602), .A2(new_n558), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(G299), .A2(new_n601), .A3(new_n594), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n602), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n877), .A2(KEYINPUT104), .A3(G299), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n873), .A2(new_n874), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(KEYINPUT41), .ZN(new_n882));
  XOR2_X1   g457(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n884), .B1(new_n876), .B2(new_n878), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n869), .A2(new_n870), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n867), .B1(new_n880), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n880), .A2(new_n867), .ZN(new_n889));
  XNOR2_X1  g464(.A(G166), .B(G288), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n579), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n579), .ZN(new_n893));
  OAI21_X1  g468(.A(G290), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n691), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT42), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n888), .A2(new_n889), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n897), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n889), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n887), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G868), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n906));
  INV_X1    g481(.A(new_n816), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(G868), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n609), .B1(new_n899), .B2(new_n903), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT107), .B1(new_n911), .B2(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(G295));
  NAND2_X1  g488(.A1(new_n905), .A2(new_n909), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n531), .A2(G171), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n821), .B(new_n917), .C1(new_n567), .C2(G301), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n531), .A2(KEYINPUT70), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n531), .A2(KEYINPUT70), .ZN(new_n922));
  OAI21_X1  g497(.A(G171), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n821), .A4(new_n917), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n529), .A2(new_n530), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(new_n566), .A3(new_n522), .A4(new_n525), .ZN(new_n927));
  AOI21_X1  g502(.A(G301), .B1(new_n927), .B2(new_n920), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n868), .B1(new_n928), .B2(new_n916), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n919), .A2(new_n879), .A3(new_n925), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n821), .B1(new_n923), .B2(new_n917), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n928), .A2(new_n868), .A3(new_n916), .ZN(new_n932));
  OAI22_X1  g507(.A1(new_n931), .A2(new_n932), .B1(new_n882), .B2(new_n885), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n897), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT109), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n933), .ZN(new_n936));
  INV_X1    g511(.A(new_n897), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G37), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n930), .A2(new_n933), .A3(new_n940), .A4(new_n897), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n935), .A2(new_n938), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n935), .A2(new_n939), .A3(new_n941), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n919), .A2(new_n929), .A3(new_n925), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n876), .A2(new_n878), .A3(new_n884), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT110), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n881), .A2(KEYINPUT41), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n876), .A2(new_n950), .A3(new_n878), .A4(new_n884), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n929), .A2(new_n879), .A3(new_n918), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n897), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n945), .A2(KEYINPUT43), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n915), .B1(new_n944), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n942), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n945), .A2(new_n958), .A3(new_n955), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n957), .A2(new_n961), .ZN(G397));
  NOR2_X1   g537(.A1(new_n836), .A2(G1384), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n467), .A2(new_n471), .A3(G40), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n800), .B(new_n803), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(new_n769), .ZN(new_n969));
  INV_X1    g544(.A(new_n967), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT127), .B(KEYINPUT46), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  NOR2_X1   g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT111), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(new_n967), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT48), .Z(new_n981));
  XNOR2_X1  g556(.A(new_n768), .B(new_n971), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n968), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n717), .B(new_n721), .Z(new_n984));
  OAI21_X1  g559(.A(new_n970), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n718), .A2(new_n721), .ZN(new_n987));
  OAI22_X1  g562(.A1(new_n983), .A2(new_n987), .B1(G2067), .B2(new_n800), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n970), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n977), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT113), .B1(new_n836), .B2(G1384), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n993));
  INV_X1    g568(.A(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n830), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n966), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G8), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  OAI21_X1  g575(.A(G1981), .B1(new_n575), .B2(new_n578), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n575), .A2(new_n578), .A3(G1981), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1000), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1003), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(KEYINPUT49), .A3(new_n1001), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n999), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n1009));
  INV_X1    g584(.A(G1976), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G288), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n998), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n1014));
  INV_X1    g589(.A(G288), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G1976), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n999), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1013), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1012), .A2(new_n1014), .A3(new_n999), .A4(new_n1016), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1008), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(G8), .B1(new_n516), .B2(new_n520), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n1021), .B(KEYINPUT55), .Z(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n965), .B1(new_n996), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n994), .B1(new_n496), .B2(new_n505), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G2090), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n966), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1971), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1022), .B(G8), .C1(new_n1028), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1020), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1007), .A2(new_n1010), .A3(new_n1015), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1003), .B(KEYINPUT115), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n999), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT116), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1038), .A2(new_n1045), .A3(new_n1042), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT63), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1022), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n992), .A2(new_n995), .A3(KEYINPUT50), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n966), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1034), .B1(G2090), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1048), .A2(new_n1036), .A3(new_n1055), .A4(new_n1007), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n992), .A2(new_n995), .A3(new_n1030), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n965), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1966), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1024), .A2(new_n755), .A3(new_n1026), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1060), .A2(KEYINPUT117), .A3(new_n1061), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(G8), .A3(new_n567), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1047), .B1(new_n1056), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1047), .B1(new_n1070), .B2(new_n1049), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1068), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1020), .A2(new_n1071), .A3(new_n1036), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1044), .A2(new_n1046), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  XOR2_X1   g649(.A(KEYINPUT118), .B(G1956), .Z(new_n1075));
  NAND2_X1  g650(.A1(new_n1052), .A2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT119), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1029), .A2(new_n966), .A3(new_n1031), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G299), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n872), .A2(KEYINPUT57), .A3(new_n558), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1080), .A2(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1024), .A2(KEYINPUT120), .A3(new_n1026), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT120), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n1086), .A2(new_n1087), .A3(G1348), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n965), .B1(new_n992), .B2(new_n995), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n803), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n877), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1093), .A2(new_n1076), .A3(new_n1079), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1085), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1085), .A2(KEYINPUT122), .A3(new_n1094), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT61), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1080), .A2(new_n1084), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1097), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1086), .A2(new_n1087), .A3(G1348), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n877), .A4(new_n1090), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT58), .B(G1341), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1032), .A2(G1996), .B1(new_n1089), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT121), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  OAI221_X1 g683(.A(new_n1108), .B1(new_n1089), .B2(new_n1105), .C1(new_n1032), .C2(G1996), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n545), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT59), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1107), .A2(new_n1109), .A3(new_n1112), .A4(new_n545), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1101), .A2(new_n1104), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1102), .A2(new_n602), .A3(new_n1090), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1103), .B1(new_n1116), .B2(new_n1092), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1085), .A2(KEYINPUT61), .A3(new_n1094), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT123), .Z(new_n1120));
  AOI21_X1  g695(.A(new_n1096), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1086), .A2(new_n1087), .A3(G1961), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G2078), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1057), .A2(KEYINPUT53), .A3(new_n1059), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1123), .A2(KEYINPUT125), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1125), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1122), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1130), .B1(new_n1032), .B2(G2078), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(G301), .B(KEYINPUT54), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n466), .A2(new_n470), .ZN(new_n1135));
  AND4_X1   g710(.A1(KEYINPUT53), .A2(new_n1029), .A3(new_n1124), .A4(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(G40), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n964), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1133), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1123), .A2(new_n1131), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1056), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1067), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1064), .A2(KEYINPUT124), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1145), .A2(G8), .A3(new_n531), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1064), .A2(G168), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1147), .A2(new_n1148), .A3(G8), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1143), .A2(G168), .A3(new_n1144), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1151), .B2(G8), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1134), .B(new_n1141), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1074), .B1(new_n1121), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1132), .A2(G171), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n1056), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1150), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1151), .A2(G8), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT51), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1149), .ZN(new_n1161));
  AOI21_X1  g736(.A(G168), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(G8), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT62), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1156), .B1(new_n1158), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT126), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(new_n1156), .C1(new_n1158), .C2(new_n1164), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1154), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n979), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n985), .B1(new_n1171), .B2(new_n967), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1172), .B(KEYINPUT112), .Z(new_n1173));
  OAI21_X1  g748(.A(new_n991), .B1(new_n1169), .B2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g749(.A(new_n955), .ZN(new_n1176));
  NAND4_X1  g750(.A1(new_n1176), .A2(new_n939), .A3(new_n941), .A4(new_n935), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n943), .B1(new_n1177), .B2(KEYINPUT43), .ZN(new_n1178));
  INV_X1    g752(.A(G227), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n652), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n862), .B2(new_n864), .ZN(new_n1181));
  NOR2_X1   g755(.A1(G229), .A2(new_n460), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n1178), .A2(new_n1181), .A3(new_n1182), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


