//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT84), .ZN(new_n189));
  INV_X1    g003(.A(G113), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n190), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT5), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G116), .B(G119), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT2), .A2(G113), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT67), .B1(new_n202), .B2(new_n190), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n204), .A2(KEYINPUT2), .A3(G113), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n200), .B(new_n201), .C1(new_n203), .C2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n199), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(G107), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n208), .A2(G107), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n207), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n201), .B1(new_n205), .B2(new_n203), .ZN(new_n221));
  INV_X1    g035(.A(new_n200), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n209), .A2(new_n212), .A3(new_n214), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G101), .ZN(new_n226));
  AOI22_X1  g040(.A1(new_n223), .A2(new_n206), .B1(new_n226), .B2(new_n215), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(G101), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT78), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n225), .A2(new_n228), .A3(new_n231), .A4(G101), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n220), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT83), .A2(KEYINPUT6), .ZN(new_n236));
  NOR3_X1   g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n220), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n230), .A2(new_n232), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n223), .A2(new_n206), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n226), .A2(new_n215), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n238), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n235), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n238), .B(new_n235), .C1(new_n239), .C2(new_n242), .ZN(new_n246));
  INV_X1    g060(.A(new_n236), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n237), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT1), .B1(new_n250), .B2(G146), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(G146), .ZN(new_n252));
  INV_X1    g066(.A(G146), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n253), .A2(G143), .ZN(new_n254));
  OAI211_X1 g068(.A(G128), .B(new_n251), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n250), .A2(G146), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n256), .B(new_n257), .C1(KEYINPUT1), .C2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G125), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(KEYINPUT0), .A2(G128), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n256), .A2(new_n257), .B1(new_n263), .B2(KEYINPUT64), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  OR2_X1    g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G143), .B(G146), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n264), .A2(new_n268), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G224), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n272), .B(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n189), .B1(new_n249), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n236), .B1(new_n234), .B2(new_n235), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n234), .A2(new_n235), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT84), .A3(new_n275), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n274), .A2(KEYINPUT86), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n274), .A2(KEYINPUT7), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n262), .A2(new_n271), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT7), .B(new_n274), .C1(new_n272), .C2(KEYINPUT86), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n194), .A2(KEYINPUT85), .ZN(new_n289));
  OAI21_X1  g103(.A(G113), .B1(new_n196), .B2(KEYINPUT5), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT85), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n289), .A2(new_n198), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n219), .B1(new_n293), .B2(new_n206), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n235), .B(KEYINPUT8), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n215), .A2(new_n218), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n207), .B2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n287), .B(new_n288), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n246), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n284), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n188), .B1(new_n283), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n188), .ZN(new_n303));
  AOI211_X1 g117(.A(new_n303), .B(new_n300), .C1(new_n277), .C2(new_n282), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n187), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT9), .B(G234), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT72), .B(G217), .Z(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n273), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n250), .A2(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n258), .A2(G143), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G134), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n311), .A3(G134), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT89), .ZN(new_n317));
  INV_X1    g131(.A(G122), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G116), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n191), .A2(KEYINPUT89), .A3(G122), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n191), .A2(G122), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n211), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n319), .A2(new_n320), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT14), .ZN(new_n327));
  OAI211_X1 g141(.A(KEYINPUT90), .B(new_n323), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT90), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n319), .B2(new_n320), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n322), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n327), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n325), .B1(new_n333), .B2(G107), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT13), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n311), .A2(new_n335), .A3(G134), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n314), .A2(new_n315), .A3(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n310), .A2(new_n311), .A3(new_n335), .A4(G134), .ZN(new_n338));
  INV_X1    g152(.A(new_n324), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n211), .B1(new_n321), .B2(new_n323), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n309), .B1(new_n334), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n309), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n330), .A2(new_n322), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n345), .A2(KEYINPUT90), .B1(new_n327), .B2(new_n326), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n211), .B1(new_n346), .B2(new_n331), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n341), .B(new_n344), .C1(new_n347), .C2(new_n325), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n334), .A2(new_n342), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT91), .B1(new_n351), .B2(new_n344), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n284), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G478), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(KEYINPUT15), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(KEYINPUT15), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n359), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n284), .B(new_n361), .C1(new_n350), .C2(new_n352), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G113), .B(G122), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n364), .B(new_n208), .ZN(new_n365));
  NOR2_X1   g179(.A1(G237), .A2(G953), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(G143), .A3(G214), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(G143), .B1(new_n366), .B2(G214), .ZN(new_n369));
  OAI21_X1  g183(.A(G131), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n369), .ZN(new_n371));
  INV_X1    g185(.A(G131), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n367), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT17), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(KEYINPUT17), .B(G131), .C1(new_n368), .C2(new_n369), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT16), .ZN(new_n379));
  INV_X1    g193(.A(G140), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n261), .A2(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n381), .B1(new_n384), .B2(new_n379), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n253), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n387));
  OAI211_X1 g201(.A(G146), .B(new_n381), .C1(new_n384), .C2(new_n379), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(KEYINPUT73), .A3(new_n253), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n378), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G125), .B(G140), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n253), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT18), .B(G131), .C1(new_n368), .C2(new_n369), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT18), .A2(G131), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n371), .A2(new_n367), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n365), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n365), .ZN(new_n400));
  INV_X1    g214(.A(new_n398), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n400), .B(new_n401), .C1(new_n378), .C2(new_n391), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n284), .B1(new_n399), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G475), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n273), .A2(G952), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(G234), .B2(G237), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT21), .B(G898), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(KEYINPUT93), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n284), .B(new_n273), .C1(G234), .C2(G237), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n370), .A2(new_n373), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT19), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n393), .B(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n415), .B(new_n388), .C1(G146), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n365), .B1(new_n418), .B2(new_n398), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n401), .B1(new_n378), .B2(new_n391), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n419), .B1(new_n420), .B2(new_n365), .ZN(new_n421));
  NOR2_X1   g235(.A1(G475), .A2(G902), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n414), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n389), .A2(new_n390), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n365), .B(new_n398), .C1(new_n425), .C2(new_n377), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n398), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n400), .ZN(new_n428));
  AOI211_X1 g242(.A(KEYINPUT20), .B(new_n423), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n424), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR4_X1   g245(.A1(new_n421), .A2(KEYINPUT88), .A3(KEYINPUT20), .A4(new_n423), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n404), .B(new_n412), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n305), .A2(new_n363), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G472), .ZN(new_n435));
  INV_X1    g249(.A(G137), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G134), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT11), .B1(new_n313), .B2(G137), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT11), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n436), .A3(G134), .ZN(new_n440));
  AOI211_X1 g254(.A(G131), .B(new_n437), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n440), .ZN(new_n442));
  INV_X1    g256(.A(new_n437), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n372), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n270), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n436), .B2(G134), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n436), .A2(G134), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n313), .A2(KEYINPUT65), .A3(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G131), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n439), .B1(G134), .B2(new_n436), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n313), .A2(KEYINPUT11), .A3(G137), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n372), .B(new_n443), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n451), .A2(new_n454), .A3(new_n259), .A4(new_n255), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n445), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n240), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n445), .A2(new_n223), .A3(new_n206), .A4(new_n455), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(KEYINPUT71), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(new_n460), .A3(new_n240), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(KEYINPUT28), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n458), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n463), .A2(KEYINPUT28), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n366), .A2(G210), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT26), .B(G101), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n462), .A2(KEYINPUT29), .A3(new_n464), .A4(new_n470), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n471), .A2(new_n284), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT66), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n445), .B1(new_n474), .B2(new_n455), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n451), .A2(new_n454), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT66), .B1(new_n476), .B2(new_n260), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n473), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n445), .A2(KEYINPUT30), .A3(new_n455), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n240), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n458), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n469), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT29), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT69), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n469), .B(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n455), .A2(new_n474), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n260), .A2(KEYINPUT66), .A3(new_n454), .A4(new_n451), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n445), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n463), .B1(new_n240), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n491));
  OAI211_X1 g305(.A(new_n486), .B(new_n464), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n484), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n435), .B1(new_n472), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n481), .A2(new_n458), .A3(new_n470), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT31), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n481), .A2(KEYINPUT31), .A3(new_n458), .A4(new_n470), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n464), .B1(new_n490), .B2(new_n491), .ZN(new_n499));
  INV_X1    g313(.A(new_n486), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G472), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT32), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n500), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n479), .B1(new_n489), .B2(new_n473), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n463), .B1(new_n506), .B2(new_n240), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT31), .B1(new_n507), .B2(new_n470), .ZN(new_n508));
  AND4_X1   g322(.A1(KEYINPUT31), .A2(new_n481), .A3(new_n458), .A4(new_n470), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT32), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n502), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n494), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G234), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n308), .B1(new_n514), .B2(G902), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT23), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n516), .B1(new_n195), .B2(G128), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n517), .B(new_n518), .C1(G119), .C2(new_n258), .ZN(new_n519));
  XNOR2_X1  g333(.A(G119), .B(G128), .ZN(new_n520));
  XOR2_X1   g334(.A(KEYINPUT24), .B(G110), .Z(new_n521));
  AOI22_X1  g335(.A1(new_n519), .A2(G110), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n389), .A2(new_n390), .A3(new_n522), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n519), .A2(G110), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n524), .B(new_n388), .C1(G146), .C2(new_n384), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G137), .ZN(new_n527));
  INV_X1    g341(.A(G221), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n528), .A2(new_n514), .A3(G953), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n527), .B(new_n529), .Z(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n523), .A2(new_n525), .A3(new_n530), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT25), .ZN(new_n534));
  AOI21_X1  g348(.A(G902), .B1(new_n534), .B2(KEYINPUT74), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n515), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n537), .B2(new_n536), .ZN(new_n539));
  AND2_X1   g353(.A1(new_n532), .A2(new_n533), .ZN(new_n540));
  AOI21_X1  g354(.A(G902), .B1(new_n308), .B2(new_n514), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n513), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n380), .A2(G110), .ZN(new_n545));
  INV_X1    g359(.A(G110), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G140), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G110), .B(G140), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n550), .B2(new_n552), .ZN(new_n556));
  INV_X1    g370(.A(G227), .ZN(new_n557));
  OAI22_X1  g371(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(G953), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n548), .A2(new_n549), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n551), .A2(KEYINPUT75), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT76), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n561), .A2(G227), .A3(new_n273), .A4(new_n554), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n269), .A2(new_n265), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n252), .A2(new_n254), .B1(new_n266), .B2(new_n267), .ZN(new_n565));
  INV_X1    g379(.A(new_n265), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n263), .B2(KEYINPUT64), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n215), .B2(new_n226), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT10), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n260), .A2(new_n296), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n255), .A2(new_n215), .A3(new_n218), .A4(new_n259), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT10), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n569), .A2(new_n233), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n441), .A2(new_n444), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n563), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n575), .B2(new_n574), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n255), .A2(new_n259), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n219), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n572), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n441), .A2(new_n444), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(KEYINPUT12), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT79), .A4(KEYINPUT12), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n575), .B1(new_n581), .B2(KEYINPUT80), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT80), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n580), .A2(new_n589), .A3(new_n572), .ZN(new_n590));
  AOI21_X1  g404(.A(KEYINPUT12), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT81), .B(new_n578), .C1(new_n587), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n563), .ZN(new_n593));
  INV_X1    g407(.A(new_n572), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n259), .A2(new_n255), .B1(new_n215), .B2(new_n218), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT80), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n582), .A3(new_n590), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT12), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n599), .A2(new_n585), .A3(new_n586), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT81), .B1(new_n600), .B2(new_n578), .ZN(new_n601));
  OAI211_X1 g415(.A(G469), .B(new_n577), .C1(new_n593), .C2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G469), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n284), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n576), .B1(new_n587), .B2(new_n591), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n569), .A2(new_n233), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n571), .A2(new_n573), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n606), .A2(new_n607), .A3(new_n575), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n575), .B1(new_n606), .B2(new_n607), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n563), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n604), .B1(new_n611), .B2(new_n603), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n528), .B1(new_n307), .B2(new_n284), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT82), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT82), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n617), .B(new_n614), .C1(new_n602), .C2(new_n612), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n434), .A2(new_n544), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT94), .B(G101), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G3));
  NAND2_X1  g436(.A1(new_n613), .A2(new_n615), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n617), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n435), .B1(new_n510), .B2(new_n284), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n501), .A2(new_n503), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n625), .A2(new_n626), .A3(new_n543), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n614), .B1(new_n602), .B2(new_n612), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT82), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n624), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n619), .A2(KEYINPUT95), .A3(new_n627), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n635));
  INV_X1    g449(.A(new_n187), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n281), .A2(KEYINPUT84), .A3(new_n275), .ZN(new_n637));
  AOI21_X1  g451(.A(KEYINPUT84), .B1(new_n281), .B2(new_n275), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n301), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n303), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n188), .B(new_n301), .C1(new_n637), .C2(new_n638), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n636), .B(new_n411), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n404), .B1(new_n431), .B2(new_n432), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n348), .A2(new_n349), .ZN(new_n644));
  INV_X1    g458(.A(new_n334), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n645), .A2(KEYINPUT91), .A3(new_n341), .A4(new_n344), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n644), .A2(new_n646), .A3(new_n343), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n344), .A2(KEYINPUT96), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n648), .B1(new_n351), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n351), .B2(new_n650), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n354), .A2(G902), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n353), .A2(new_n354), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n643), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n635), .B1(new_n642), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n187), .B(new_n412), .C1(new_n302), .C2(new_n304), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n660), .A2(KEYINPUT97), .A3(new_n657), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n634), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT34), .B(G104), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  INV_X1    g479(.A(KEYINPUT98), .ZN(new_n666));
  INV_X1    g480(.A(new_n362), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n361), .B1(new_n647), .B2(new_n284), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n426), .A2(new_n428), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n422), .A3(new_n413), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n424), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n404), .A3(new_n412), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n666), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  AOI22_X1  g488(.A1(new_n424), .A2(new_n671), .B1(new_n403), .B2(G475), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n363), .A2(KEYINPUT98), .A3(new_n412), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n305), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n632), .A2(new_n633), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT35), .B(G107), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  OR2_X1    g495(.A1(new_n625), .A2(new_n626), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n531), .A2(KEYINPUT36), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n526), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n541), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n539), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n434), .A2(new_n619), .A3(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n406), .B1(new_n410), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n675), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n363), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n305), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n504), .A2(new_n512), .ZN(new_n698));
  INV_X1    g512(.A(new_n494), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n687), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n697), .A2(new_n619), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G128), .ZN(G30));
  NAND2_X1  g516(.A1(new_n640), .A2(new_n641), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n459), .A2(new_n461), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI22_X1  g521(.A1(new_n500), .A2(new_n707), .B1(new_n507), .B2(new_n470), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n708), .B2(G902), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n698), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n643), .A2(new_n363), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n686), .A2(new_n636), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n705), .A2(new_n710), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT40), .ZN(new_n715));
  XOR2_X1   g529(.A(new_n693), .B(KEYINPUT39), .Z(new_n716));
  NAND3_X1  g530(.A1(new_n624), .A2(new_n629), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(KEYINPUT100), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n619), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n715), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n717), .A2(KEYINPUT100), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n619), .A2(new_n719), .A3(new_n716), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT40), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n714), .B1(new_n721), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n250), .ZN(G45));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n643), .A2(new_n656), .A3(new_n694), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n305), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n643), .A2(new_n656), .A3(new_n694), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n730), .A2(new_n703), .A3(KEYINPUT101), .A4(new_n187), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n729), .A2(new_n619), .A3(new_n731), .A4(new_n700), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NOR2_X1   g547(.A1(new_n611), .A2(new_n603), .ZN(new_n734));
  AOI211_X1 g548(.A(G469), .B(G902), .C1(new_n605), .C2(new_n610), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n734), .A2(new_n735), .A3(new_n614), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n513), .A2(new_n543), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n738), .B1(new_n659), .B2(new_n661), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n678), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  INV_X1    g557(.A(KEYINPUT102), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n501), .A2(KEYINPUT32), .A3(new_n503), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n511), .B1(new_n510), .B2(new_n502), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n699), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n686), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n433), .A2(new_n363), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n703), .A3(new_n187), .A4(new_n736), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n744), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n187), .B(new_n736), .C1(new_n302), .C2(new_n304), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(new_n700), .A3(KEYINPUT102), .A4(new_n749), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  NAND2_X1  g570(.A1(new_n736), .A2(new_n412), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n305), .A2(new_n757), .A3(new_n711), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n497), .A2(new_n498), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n462), .A2(new_n464), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n500), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n503), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT103), .ZN(new_n763));
  AOI21_X1  g577(.A(G902), .B1(new_n759), .B2(new_n505), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n763), .B1(new_n764), .B2(new_n435), .ZN(new_n765));
  OAI211_X1 g579(.A(KEYINPUT103), .B(G472), .C1(new_n501), .C2(G902), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n543), .B(new_n762), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  AOI211_X1 g583(.A(new_n687), .B(new_n762), .C1(new_n765), .C2(new_n766), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n752), .A2(new_n728), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G125), .ZN(G27));
  OAI21_X1  g587(.A(KEYINPUT104), .B1(new_n745), .B2(new_n746), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n504), .A2(new_n512), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n699), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n640), .A2(new_n187), .A3(new_n641), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(new_n623), .A3(new_n728), .ZN(new_n779));
  INV_X1    g593(.A(new_n543), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n777), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT42), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n778), .A2(new_n623), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n728), .A2(KEYINPUT42), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n544), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n372), .ZN(G33));
  INV_X1    g601(.A(KEYINPUT105), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n696), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n544), .A3(new_n783), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  OR2_X1    g605(.A1(new_n593), .A2(new_n601), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(KEYINPUT106), .A3(KEYINPUT45), .A4(new_n577), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT106), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n577), .B1(new_n593), .B2(new_n601), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n603), .B1(new_n795), .B2(new_n796), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n604), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n735), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n802), .B2(new_n801), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n615), .A3(new_n716), .ZN(new_n805));
  INV_X1    g619(.A(new_n643), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT107), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n643), .A2(KEYINPUT107), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n656), .A2(KEYINPUT43), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT43), .B1(new_n806), .B2(new_n656), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT44), .A3(new_n682), .A4(new_n686), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT44), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n643), .B(new_n807), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n812), .B1(new_n817), .B2(new_n810), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n682), .A2(new_n686), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n778), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n815), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n805), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n436), .ZN(G39));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n513), .A3(new_n543), .A4(new_n730), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n615), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT47), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n799), .A2(KEYINPUT46), .A3(new_n800), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT46), .B1(new_n799), .B2(new_n800), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n828), .A2(new_n829), .A3(new_n735), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n827), .B1(new_n830), .B2(new_n614), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n825), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(new_n380), .ZN(G42));
  NOR2_X1   g647(.A1(new_n734), .A2(new_n735), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT49), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n543), .A2(new_n614), .A3(new_n636), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(new_n656), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n817), .ZN(new_n838));
  OR4_X1    g652(.A1(new_n705), .A2(new_n837), .A3(new_n710), .A4(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n778), .A2(new_n737), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n814), .A2(new_n406), .A3(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n770), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n780), .A2(new_n406), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n710), .A2(new_n737), .A3(new_n778), .A4(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n806), .A3(new_n655), .A4(new_n654), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT51), .B1(new_n846), .B2(KEYINPUT109), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n814), .A2(new_n406), .A3(new_n767), .ZN(new_n848));
  NOR4_X1   g662(.A1(new_n848), .A2(new_n187), .A3(new_n705), .A4(new_n737), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT50), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n826), .A2(new_n831), .ZN(new_n851));
  INV_X1    g665(.A(new_n834), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n615), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n848), .A2(new_n778), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n850), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n847), .B(new_n857), .C1(KEYINPUT109), .C2(new_n846), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n783), .A2(new_n860), .A3(new_n686), .A4(new_n730), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n695), .A2(new_n669), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n778), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n619), .A2(new_n700), .A3(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n657), .B1(new_n669), .B2(new_n643), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n642), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n632), .A2(new_n633), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n434), .B(new_n619), .C1(new_n688), .C2(new_n544), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AND4_X1   g684(.A1(new_n747), .A2(new_n624), .A3(new_n629), .A4(new_n686), .ZN(new_n871));
  AOI22_X1  g685(.A1(new_n871), .A2(new_n697), .B1(new_n770), .B2(new_n771), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  INV_X1    g687(.A(new_n305), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n628), .A2(new_n687), .A3(new_n694), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n710), .A4(new_n712), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n872), .A2(new_n873), .A3(new_n732), .A4(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n782), .A2(new_n785), .A3(new_n790), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n732), .A2(new_n701), .A3(new_n772), .A4(new_n876), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n870), .A2(new_n877), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n767), .A2(new_n758), .B1(new_n738), .B2(new_n678), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n755), .A2(new_n739), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT108), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT108), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n739), .A2(new_n755), .A3(new_n882), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n859), .B1(new_n881), .B2(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n881), .A2(new_n887), .ZN(new_n889));
  INV_X1    g703(.A(new_n772), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n697), .A2(new_n619), .A3(new_n700), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT52), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n892), .A2(new_n859), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n888), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT54), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n892), .A2(KEYINPUT53), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n883), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n782), .A2(new_n785), .A3(new_n790), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n897), .A2(new_n877), .A3(new_n880), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n888), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n895), .B1(KEYINPUT54), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n857), .A2(new_n846), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n904), .A2(KEYINPUT51), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n777), .A2(new_n780), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n841), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT48), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n405), .B1(new_n844), .B2(new_n658), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n908), .B(new_n909), .C1(new_n752), .C2(new_n848), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT110), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n858), .A2(new_n903), .A3(new_n905), .A4(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(G952), .A2(G953), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n839), .B1(new_n912), .B2(new_n913), .ZN(G75));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n249), .B(KEYINPUT111), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT112), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n275), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n284), .B1(new_n888), .B2(new_n901), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(G210), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n915), .B(new_n919), .C1(new_n921), .C2(KEYINPUT113), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(KEYINPUT113), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n273), .A2(G952), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT114), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT56), .B1(new_n920), .B2(G210), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n919), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n923), .A2(new_n927), .ZN(G51));
  INV_X1    g742(.A(KEYINPUT115), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n284), .B(new_n799), .C1(new_n888), .C2(new_n901), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n604), .B(KEYINPUT57), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n605), .A2(new_n610), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n930), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n936), .B2(new_n924), .ZN(new_n937));
  INV_X1    g751(.A(new_n924), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n902), .B(KEYINPUT54), .ZN(new_n939));
  AOI22_X1  g753(.A1(new_n939), .A2(new_n931), .B1(new_n610), .B2(new_n605), .ZN(new_n940));
  OAI211_X1 g754(.A(KEYINPUT115), .B(new_n938), .C1(new_n940), .C2(new_n930), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n937), .A2(new_n941), .ZN(G54));
  NAND3_X1  g756(.A1(new_n920), .A2(KEYINPUT58), .A3(G475), .ZN(new_n943));
  OR3_X1    g757(.A1(new_n943), .A2(KEYINPUT116), .A3(new_n421), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT116), .B1(new_n943), .B2(new_n421), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n924), .B1(new_n943), .B2(new_n421), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G60));
  AND2_X1   g761(.A1(new_n649), .A2(new_n652), .ZN(new_n948));
  XNOR2_X1  g762(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n949));
  NAND2_X1  g763(.A1(G478), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n903), .B2(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n939), .A2(new_n948), .A3(new_n951), .ZN(new_n953));
  INV_X1    g767(.A(new_n925), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G63));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n888), .B2(new_n901), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n684), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n925), .B1(new_n958), .B2(new_n540), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n961), .A2(KEYINPUT118), .B1(new_n684), .B2(new_n958), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT118), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n925), .C1(new_n958), .C2(new_n540), .ZN(new_n965));
  AOI211_X1 g779(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT119), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n961), .A2(KEYINPUT118), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n965), .A3(new_n959), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n962), .B1(new_n966), .B2(new_n971), .ZN(G66));
  AOI21_X1  g786(.A(new_n273), .B1(new_n408), .B2(G224), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT120), .ZN(new_n974));
  AND4_X1   g788(.A1(new_n884), .A2(new_n886), .A3(new_n868), .A4(new_n869), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(G953), .ZN(new_n976));
  INV_X1    g790(.A(G898), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n916), .B1(new_n977), .B2(G953), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n976), .B(new_n978), .Z(G69));
  OAI21_X1  g793(.A(G953), .B1(new_n557), .B2(new_n692), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT124), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n872), .A2(new_n732), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n724), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT40), .B1(new_n722), .B2(new_n723), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n985), .B(KEYINPUT62), .C1(new_n988), .C2(new_n714), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n725), .B2(new_n984), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n544), .A2(new_n821), .A3(new_n866), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n718), .A2(new_n720), .A3(new_n993), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n832), .A2(new_n823), .A3(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n992), .A2(KEYINPUT122), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT122), .B1(new_n992), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n273), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n506), .B(KEYINPUT121), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(new_n417), .Z(new_n1000));
  AOI21_X1  g814(.A(new_n983), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  OAI22_X1  g816(.A1(new_n851), .A2(new_n825), .B1(new_n805), .B2(new_n822), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n906), .A2(new_n874), .A3(new_n712), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n985), .B(new_n878), .C1(new_n805), .C2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1005), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n832), .A2(new_n823), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1007), .A2(new_n1008), .A3(KEYINPUT125), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1006), .A2(new_n1009), .A3(new_n273), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1000), .B1(G900), .B2(G953), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1001), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n998), .A2(new_n983), .A3(new_n1000), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n982), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n992), .A2(new_n995), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT122), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n992), .A2(KEYINPUT122), .A3(new_n995), .ZN(new_n1021));
  AOI21_X1  g835(.A(G953), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1000), .ZN(new_n1023));
  OAI21_X1  g837(.A(KEYINPUT123), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1025));
  AND4_X1   g839(.A1(new_n982), .A2(new_n1024), .A3(new_n1025), .A4(new_n1016), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1017), .A2(new_n1026), .ZN(G72));
  NAND3_X1  g841(.A1(new_n1020), .A2(new_n975), .A3(new_n1021), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  AOI211_X1 g844(.A(new_n469), .B(new_n507), .C1(new_n1028), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT127), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1030), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n483), .B2(new_n495), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n894), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1032), .B1(new_n894), .B2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n938), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1006), .A2(new_n1009), .A3(new_n975), .ZN(new_n1038));
  AOI211_X1 g852(.A(new_n470), .B(new_n482), .C1(new_n1038), .C2(new_n1030), .ZN(new_n1039));
  NOR3_X1   g853(.A1(new_n1031), .A2(new_n1037), .A3(new_n1039), .ZN(G57));
endmodule


