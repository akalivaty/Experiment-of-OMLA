//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT65), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n466), .A2(new_n467), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n464), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(new_n468), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n478), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n464), .A2(G2105), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n487), .A2(G124), .B1(G136), .B2(new_n488), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n467), .C2(G112), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT68), .ZN(G162));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n483), .B2(new_n484), .ZN(new_n494));
  AND2_X1   g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(G138), .B1(new_n462), .B2(new_n463), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(new_n478), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n485), .A2(new_n467), .A3(KEYINPUT4), .A4(G138), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n469), .A2(G102), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n496), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G651), .ZN(new_n507));
  AND2_X1   g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n505), .A2(new_n507), .A3(G543), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(new_n504), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n514), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(new_n510), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT70), .B(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n508), .A2(new_n522), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n513), .A2(KEYINPUT69), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G51), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n509), .A2(G63), .ZN(new_n526));
  NAND2_X1  g101(.A1(G76), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(G651), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n527), .B2(new_n504), .ZN(new_n531));
  NAND4_X1  g106(.A1(new_n521), .A2(new_n525), .A3(new_n530), .A4(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  XOR2_X1   g108(.A(KEYINPUT5), .B(G543), .Z(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  INV_X1    g110(.A(G77), .ZN(new_n536));
  INV_X1    g111(.A(G543), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n534), .A2(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT71), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI221_X1 g115(.A(KEYINPUT71), .B1(new_n536), .B2(new_n537), .C1(new_n534), .C2(new_n535), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n540), .A2(G651), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n540), .A2(KEYINPUT72), .A3(new_n541), .A4(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n519), .A2(G90), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n523), .A2(G52), .A3(new_n524), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  AND3_X1   g126(.A1(new_n523), .A2(G43), .A3(new_n524), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n553), .A2(new_n504), .B1(new_n510), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g135(.A1(G319), .A2(G483), .A3(G661), .A4(new_n560), .ZN(G188));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n513), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n519), .A2(G91), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n504), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(G299));
  NAND2_X1  g144(.A1(new_n519), .A2(G87), .ZN(new_n570));
  INV_X1    g145(.A(new_n513), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n534), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G48), .B2(new_n571), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n519), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  NAND3_X1  g155(.A1(new_n523), .A2(G47), .A3(new_n524), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n519), .A2(G85), .ZN(new_n582));
  INV_X1    g157(.A(G60), .ZN(new_n583));
  INV_X1    g158(.A(G72), .ZN(new_n584));
  OAI22_X1  g159(.A1(new_n534), .A2(new_n583), .B1(new_n584), .B2(new_n537), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT73), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(KEYINPUT73), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n581), .B(new_n582), .C1(new_n587), .C2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n504), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n523), .A2(G54), .A3(new_n524), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n593), .A2(KEYINPUT74), .A3(new_n594), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n510), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n597), .A2(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT75), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n602), .A2(new_n601), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT74), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT74), .B1(new_n593), .B2(new_n594), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT75), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n591), .B1(new_n612), .B2(new_n590), .ZN(G284));
  AOI21_X1  g188(.A(new_n591), .B1(new_n612), .B2(new_n590), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  OAI21_X1  g195(.A(G868), .B1(new_n611), .B2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n556), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n485), .A2(new_n469), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT76), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2100), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT77), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n478), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  AND2_X1   g210(.A1(new_n487), .A2(G123), .ZN(new_n636));
  AOI211_X1 g211(.A(new_n635), .B(new_n636), .C1(G135), .C2(new_n488), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n628), .A2(new_n629), .A3(new_n638), .ZN(G156));
  XOR2_X1   g214(.A(KEYINPUT15), .B(G2435), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2438), .ZN(new_n641));
  XOR2_X1   g216(.A(G2427), .B(G2430), .Z(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT80), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT81), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n652), .A2(new_n655), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n658), .A2(G14), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT82), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n662), .A3(new_n659), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n661), .A2(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT17), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  OR3_X1    g245(.A1(new_n667), .A2(new_n665), .A3(new_n668), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n665), .A3(new_n668), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G2096), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2100), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1981), .B(G1986), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT83), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  NOR2_X1   g271(.A1(G16), .A2(G23), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  INV_X1    g273(.A(G288), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT89), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n701));
  NAND2_X1  g276(.A1(G288), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G16), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n698), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT33), .B(G1976), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G305), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(new_n704), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G6), .B2(new_n704), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT32), .B(G1981), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n704), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n704), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(G1971), .Z(new_n717));
  NAND4_X1  g292(.A1(new_n707), .A2(new_n713), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT34), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n487), .A2(G119), .B1(G131), .B2(new_n488), .ZN(new_n722));
  OAI221_X1 g297(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n467), .C2(G107), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT84), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n721), .B1(new_n725), .B2(new_n720), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT85), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT86), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(KEYINPUT86), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n704), .A2(G24), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT87), .Z(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G290), .B2(G16), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1986), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n730), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  OR3_X1    g311(.A1(new_n719), .A2(KEYINPUT36), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(KEYINPUT36), .B1(new_n719), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT31), .B(G11), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G28), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT96), .Z(new_n743));
  OAI21_X1  g318(.A(new_n720), .B1(new_n741), .B2(G28), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n637), .A2(G29), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(KEYINPUT95), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n720), .B1(KEYINPUT24), .B2(G34), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(KEYINPUT24), .B2(G34), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n480), .B2(G29), .ZN(new_n751));
  OAI221_X1 g326(.A(new_n747), .B1(KEYINPUT95), .B2(new_n746), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n704), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n704), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n720), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT28), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n487), .A2(G128), .ZN(new_n758));
  OAI221_X1 g333(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n467), .C2(G116), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n488), .A2(G140), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n757), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n754), .A2(G1966), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n755), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n751), .A2(new_n748), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n752), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(G162), .A2(new_n720), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n720), .B2(G35), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT29), .B(G2090), .Z(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n704), .A2(G20), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT23), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n616), .B2(new_n704), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G1956), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n770), .A2(new_n771), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n768), .A2(new_n772), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n779));
  NAND2_X1  g354(.A1(G103), .A2(G2104), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n478), .B2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n781), .A2(new_n782), .B1(new_n488), .B2(G139), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT92), .Z(new_n784));
  AOI22_X1  g359(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(new_n467), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n784), .A2(KEYINPUT93), .A3(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT93), .B1(new_n784), .B2(new_n786), .ZN(new_n789));
  OAI21_X1  g364(.A(G29), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G33), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(G29), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n792), .A2(G2072), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n720), .A2(G32), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n487), .A2(G129), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n488), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT26), .Z(new_n798));
  NAND3_X1  g373(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n794), .B1(new_n800), .B2(new_n720), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT27), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1996), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n720), .A2(G27), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT98), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n502), .B2(G29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2078), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n803), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G171), .A2(new_n704), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G5), .B2(new_n704), .ZN(new_n813));
  INV_X1    g388(.A(G1961), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n814), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n704), .A2(G19), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n556), .B2(new_n704), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT91), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT90), .B(G1341), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n815), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n778), .A2(new_n793), .A3(new_n811), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n792), .A2(G2072), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT94), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n704), .A2(G4), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n612), .B2(new_n704), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1348), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n739), .A2(new_n823), .A3(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NAND2_X1  g406(.A1(G80), .A2(G543), .ZN(new_n832));
  INV_X1    g407(.A(G67), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n534), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n519), .A2(G93), .B1(new_n834), .B2(G651), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n523), .A2(G55), .A3(new_n524), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n835), .A2(KEYINPUT100), .A3(new_n836), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n556), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n556), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n842), .A2(new_n837), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n612), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  INV_X1    g423(.A(G860), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n849), .B1(new_n839), .B2(new_n840), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(G145));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n637), .B(G160), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(G162), .Z(new_n857));
  OAI21_X1  g432(.A(G164), .B1(new_n788), .B2(new_n789), .ZN(new_n858));
  INV_X1    g433(.A(new_n789), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n859), .A2(new_n502), .A3(new_n787), .ZN(new_n860));
  INV_X1    g435(.A(new_n761), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n861), .B1(new_n858), .B2(new_n860), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n487), .A2(G130), .B1(G142), .B2(new_n488), .ZN(new_n865));
  OAI221_X1 g440(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n467), .C2(G118), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n625), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n863), .A2(new_n864), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n858), .A2(new_n860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n761), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n870), .B1(new_n872), .B2(new_n862), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n857), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n724), .B(new_n799), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n868), .B1(new_n863), .B2(new_n864), .ZN(new_n876));
  INV_X1    g451(.A(new_n857), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n872), .A2(new_n862), .A3(new_n870), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(KEYINPUT101), .B(G37), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n875), .B1(new_n874), .B2(new_n879), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n855), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n885), .A2(KEYINPUT40), .A3(new_n880), .A4(new_n881), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n884), .A2(new_n886), .ZN(G395));
  NAND2_X1  g462(.A1(new_n608), .A2(new_n616), .ZN(new_n888));
  OAI211_X1 g463(.A(G299), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n889), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n890), .A2(KEYINPUT103), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n844), .B1(new_n611), .B2(G559), .ZN(new_n898));
  INV_X1    g473(.A(new_n843), .ZN(new_n899));
  INV_X1    g474(.A(new_n840), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT100), .B1(new_n835), .B2(new_n836), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n842), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n903), .A2(new_n619), .A3(new_n610), .A4(new_n604), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n890), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n888), .B2(new_n889), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n898), .A3(new_n904), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n906), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n908), .A2(new_n909), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n905), .A2(new_n914), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n895), .A2(new_n896), .B1(new_n898), .B2(new_n904), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G290), .B(G166), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n700), .A2(G305), .A3(new_n702), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G305), .B1(new_n700), .B2(new_n702), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  XNOR2_X1  g498(.A(G290), .B(G303), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n919), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n913), .A2(new_n917), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n913), .B2(new_n917), .ZN(new_n929));
  OAI21_X1  g504(.A(G868), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT104), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n590), .B1(new_n900), .B2(new_n901), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n930), .B2(new_n932), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(G295));
  NAND2_X1  g510(.A1(new_n930), .A2(new_n932), .ZN(G331));
  AOI21_X1  g511(.A(new_n548), .B1(new_n543), .B2(new_n542), .ZN(new_n937));
  AOI21_X1  g512(.A(G286), .B1(new_n937), .B2(new_n545), .ZN(new_n938));
  AND4_X1   g513(.A1(G286), .A2(new_n544), .A3(new_n545), .A4(new_n549), .ZN(new_n939));
  OAI22_X1  g514(.A1(new_n938), .A2(new_n939), .B1(new_n841), .B2(new_n843), .ZN(new_n940));
  NAND2_X1  g515(.A1(G301), .A2(G168), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(G286), .A3(new_n545), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n899), .A2(new_n941), .A3(new_n902), .A4(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n895), .A3(new_n896), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n943), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n890), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n926), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n926), .B1(new_n945), .B2(new_n947), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n950), .A2(G37), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n881), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n926), .B1(new_n910), .B2(new_n946), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n944), .A2(new_n892), .A3(new_n894), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n949), .B1(new_n956), .B2(new_n948), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT44), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n956), .A2(new_n949), .A3(new_n948), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n945), .A2(new_n926), .A3(new_n947), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n962), .A2(new_n951), .A3(G37), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n960), .B(new_n961), .C1(new_n963), .C2(new_n949), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n958), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n959), .B1(new_n958), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(G397));
  XNOR2_X1  g542(.A(KEYINPUT106), .B(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n502), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n470), .A2(G40), .A3(new_n479), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n761), .B(G2067), .Z(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n800), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT46), .ZN(new_n977));
  INV_X1    g552(.A(G1996), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n977), .B2(new_n979), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n982));
  XNOR2_X1  g557(.A(new_n981), .B(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n799), .B(new_n978), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n974), .B1(new_n975), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT107), .Z(new_n986));
  XOR2_X1   g561(.A(new_n724), .B(new_n728), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n973), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n974), .A2(G1986), .A3(G290), .ZN(new_n990));
  XOR2_X1   g565(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n991));
  XNOR2_X1  g566(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n983), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n725), .A2(new_n728), .ZN(new_n994));
  XOR2_X1   g569(.A(new_n994), .B(KEYINPUT124), .Z(new_n995));
  NAND2_X1  g570(.A1(new_n986), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G2067), .B2(new_n761), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n974), .B1(new_n997), .B2(KEYINPUT125), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT4), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n501), .B1(new_n498), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G138), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n483), .B2(new_n484), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT4), .B1(new_n1004), .B2(new_n467), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n1006), .B2(new_n496), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n470), .A2(G40), .A3(new_n479), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G8), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT113), .Z(new_n1011));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n1012));
  OR3_X1    g587(.A1(G305), .A2(new_n1012), .A3(G1981), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(G305), .B2(G1981), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT112), .B(G86), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n578), .B1(new_n510), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G1981), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT49), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(new_n1010), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1015), .A2(KEYINPUT49), .A3(new_n1018), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n699), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1011), .B1(new_n1024), .B2(new_n1015), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1008), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1029));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n502), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(KEYINPUT108), .A3(new_n970), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1027), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G1971), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n502), .A2(new_n1036), .A3(new_n1030), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1035), .A2(new_n1008), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1038), .A2(G2090), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G303), .A2(G8), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1041), .B(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(G8), .B(new_n1009), .C1(new_n703), .C2(new_n1023), .ZN(new_n1045));
  NAND2_X1  g620(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n699), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1048), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n1047), .A2(new_n1049), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1025), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1044), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1053));
  INV_X1    g628(.A(G1966), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n972), .B1(new_n1031), .B2(new_n970), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n502), .A2(KEYINPUT114), .A3(KEYINPUT45), .A4(new_n1030), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n1030), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n502), .A2(new_n1036), .A3(new_n1030), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1036), .B1(new_n502), .B2(new_n1030), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(new_n1062), .A3(new_n972), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1054), .A2(new_n1060), .B1(new_n1063), .B2(new_n748), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1064), .A2(new_n1065), .A3(G286), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1052), .A2(new_n1050), .A3(new_n1053), .A4(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT63), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1051), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G2078), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT53), .B1(new_n1033), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1038), .A2(new_n814), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1055), .A2(new_n1059), .A3(new_n1056), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(G171), .B1(new_n1073), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT122), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(G171), .C1(new_n1073), .C2(new_n1078), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1026), .A2(new_n1008), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(new_n1076), .A3(new_n971), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1074), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT108), .B1(new_n1031), .B2(new_n970), .ZN(new_n1086));
  AOI211_X1 g661(.A(new_n1028), .B(KEYINPUT45), .C1(new_n502), .C2(new_n1030), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1083), .B(new_n1072), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1085), .B1(new_n1075), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G301), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1080), .A2(new_n1082), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1093));
  AND3_X1   g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1065), .B1(new_n1064), .B2(G168), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1098), .B2(KEYINPUT51), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1060), .A2(new_n1054), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1063), .A2(new_n748), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(G8), .B1(new_n1102), .B2(G286), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1103), .A2(KEYINPUT120), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1064), .A2(KEYINPUT119), .ZN(new_n1108));
  AOI21_X1  g683(.A(G286), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1099), .B(new_n1105), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1107), .A2(new_n1108), .A3(G8), .A4(G286), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n1114));
  XNOR2_X1  g689(.A(G299), .B(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1083), .B(new_n1117), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT115), .B(G1956), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1038), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n972), .B1(new_n1031), .B2(KEYINPUT50), .ZN(new_n1122));
  AOI21_X1  g697(.A(G1348), .B1(new_n1122), .B2(new_n1037), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1031), .A2(new_n972), .A3(G2067), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n603), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1116), .A2(new_n1121), .B1(new_n1125), .B2(KEYINPUT116), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1118), .A2(new_n1115), .A3(new_n1120), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1127), .A2(KEYINPUT61), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(new_n603), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1088), .A2(new_n1075), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1132), .A2(G301), .A3(new_n1074), .A4(new_n1077), .ZN(new_n1133));
  OAI211_X1 g708(.A(KEYINPUT54), .B(new_n1133), .C1(new_n1089), .C2(G301), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1127), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1121), .A2(new_n1116), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1125), .A2(KEYINPUT116), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1140), .A2(new_n1141), .A3(new_n1130), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1139), .B1(new_n1127), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1135), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1127), .ZN(new_n1145));
  INV_X1    g720(.A(G1348), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1124), .B1(new_n1038), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n608), .B1(new_n1147), .B2(KEYINPUT60), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n1149));
  NOR4_X1   g724(.A1(new_n1123), .A2(new_n603), .A3(new_n1149), .A4(new_n1124), .ZN(new_n1150));
  OAI22_X1  g725(.A1(new_n1148), .A2(new_n1150), .B1(KEYINPUT60), .B2(new_n1147), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1083), .B(new_n978), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  AOI22_X1  g728(.A1(new_n1152), .A2(KEYINPUT117), .B1(new_n1009), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1033), .A2(new_n1155), .A3(new_n978), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n842), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1151), .B1(new_n1157), .B2(KEYINPUT59), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1145), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1113), .A2(new_n1144), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1111), .A2(new_n1162), .A3(new_n1112), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1162), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1096), .A2(new_n1161), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1052), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1071), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(G290), .B(G1986), .Z(new_n1170));
  OAI211_X1 g745(.A(new_n986), .B(new_n988), .C1(new_n974), .C2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1000), .B1(new_n1169), .B2(new_n1171), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g747(.A1(new_n885), .A2(new_n881), .A3(new_n880), .ZN(new_n1174));
  NOR2_X1   g748(.A1(G227), .A2(new_n460), .ZN(new_n1175));
  NAND2_X1  g749(.A1(new_n695), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1176), .B1(new_n661), .B2(new_n663), .ZN(new_n1177));
  OAI21_X1  g751(.A(new_n961), .B1(new_n963), .B2(new_n949), .ZN(new_n1178));
  NAND3_X1  g752(.A1(new_n1174), .A2(new_n1177), .A3(new_n1178), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


