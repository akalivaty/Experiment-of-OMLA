//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n566, new_n567,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT67), .A2(KEYINPUT3), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT67), .A2(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(G2104), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT68), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(KEYINPUT68), .B(G2104), .C1(new_n462), .C2(new_n463), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G137), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G2105), .B1(G101), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n469), .A2(G136), .ZN(new_n482));
  INV_X1    g057(.A(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n483), .B1(new_n467), .B2(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n483), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(new_n473), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT67), .A2(KEYINPUT3), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n465), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n466), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n468), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n495), .A2(new_n483), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G126), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  OR3_X1    g079(.A1(new_n504), .A2(new_n483), .A3(G114), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n504), .B1(new_n483), .B2(G114), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n503), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n472), .A2(new_n474), .A3(new_n483), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n496), .B1(new_n509), .B2(new_n497), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n499), .A2(new_n502), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  OR3_X1    g090(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT71), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n515), .B1(new_n514), .B2(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT70), .ZN(new_n525));
  INV_X1    g100(.A(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(new_n518), .ZN(new_n529));
  INV_X1    g104(.A(G88), .ZN(new_n530));
  INV_X1    g105(.A(G50), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(G543), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n522), .B1(new_n529), .B2(new_n530), .C1(new_n531), .C2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND2_X1  g109(.A1(new_n525), .A2(new_n527), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n515), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G51), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n519), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT72), .B(G89), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(G63), .A2(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n518), .A2(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n537), .A2(new_n540), .A3(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n548), .A2(new_n532), .B1(new_n529), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n526), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n550), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AOI22_X1  g129(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n526), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n536), .A2(G43), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n538), .A2(G81), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n559), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(G53), .ZN(new_n570));
  OAI211_X1 g145(.A(KEYINPUT74), .B(new_n569), .C1(new_n532), .C2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT74), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n570), .B1(new_n572), .B2(KEYINPUT9), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n536), .B(new_n573), .C1(new_n572), .C2(KEYINPUT9), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n575));
  OR2_X1    g150(.A1(new_n575), .A2(new_n526), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n538), .A2(G91), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n571), .A2(new_n574), .A3(new_n576), .A4(new_n577), .ZN(G299));
  NAND2_X1  g153(.A1(new_n536), .A2(G49), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n538), .A2(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT75), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n579), .A2(new_n580), .A3(new_n584), .A4(new_n581), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G288));
  AOI22_X1  g162(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n526), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(G86), .B2(new_n538), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n525), .A2(G48), .A3(G543), .A4(new_n527), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT76), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n526), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n536), .A2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n538), .A2(G85), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n538), .A2(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n519), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(G54), .A2(new_n536), .B1(new_n606), .B2(G651), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT78), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT78), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n603), .A2(new_n610), .A3(new_n607), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n600), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n600), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT79), .ZN(G148));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n562), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n609), .A2(new_n611), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n623), .B1(new_n625), .B2(new_n622), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g203(.A1(new_n509), .A2(new_n465), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n469), .A2(G135), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n484), .A2(G123), .ZN(new_n635));
  NOR2_X1   g210(.A1(new_n483), .A2(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(G2096), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT82), .ZN(new_n655));
  OAI21_X1  g230(.A(G14), .B1(new_n652), .B2(new_n653), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT17), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n665), .B(new_n662), .C1(new_n658), .C2(new_n660), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n661), .A2(new_n658), .A3(new_n660), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2096), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT85), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NOR3_X1   g256(.A1(new_n675), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n675), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  NAND2_X1  g266(.A1(new_n469), .A2(G139), .ZN(new_n692));
  INV_X1    g267(.A(G127), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n475), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G115), .B2(G2104), .ZN(new_n695));
  NAND2_X1  g270(.A1(G103), .A2(G2104), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(G2105), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n697), .A2(KEYINPUT25), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT25), .ZN(new_n699));
  NOR3_X1   g274(.A1(new_n696), .A2(new_n699), .A3(G2105), .ZN(new_n700));
  OAI221_X1 g275(.A(new_n692), .B1(new_n695), .B2(new_n483), .C1(new_n698), .C2(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G33), .B(new_n701), .S(G29), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT95), .B(G2072), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G5), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G171), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G1961), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n705), .A2(G21), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G168), .B2(new_n705), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  INV_X1    g287(.A(G34), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(KEYINPUT24), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(KEYINPUT24), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G160), .B2(new_n712), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n709), .B1(G1966), .B2(new_n711), .C1(G2084), .C2(new_n717), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n704), .B(new_n718), .C1(G2084), .C2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n712), .A2(G35), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G162), .B2(new_n712), .ZN(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n712), .A2(G26), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT94), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n469), .A2(G140), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n484), .A2(G128), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n483), .A2(G116), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n728), .B1(new_n733), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G2067), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n719), .A2(new_n725), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n705), .A2(G19), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT93), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n563), .B2(new_n705), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1341), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n712), .A2(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n712), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT99), .Z(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n740), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n612), .A2(new_n705), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G4), .B2(new_n705), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n705), .A2(G20), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT23), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n616), .B2(new_n705), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT101), .B(G1956), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT31), .B(G11), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n638), .A2(new_n712), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT30), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n712), .B1(new_n760), .B2(G28), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n761), .A2(KEYINPUT98), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(KEYINPUT98), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n760), .B2(G28), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n758), .B(new_n759), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n711), .A2(G1966), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT27), .B(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n712), .A2(G32), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n469), .A2(G141), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n484), .A2(G129), .ZN(new_n771));
  NAND3_X1  g346(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT26), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(G105), .B2(new_n478), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n770), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n769), .B1(new_n777), .B2(G29), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n765), .B(new_n766), .C1(new_n768), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n757), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n768), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT97), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n751), .A2(new_n752), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n736), .A2(new_n747), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(G6), .A2(G16), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G305), .B2(new_n705), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1981), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n705), .A2(G23), .ZN(new_n789));
  INV_X1    g364(.A(new_n582), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(new_n705), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT33), .B(G1976), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n705), .A2(G22), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT90), .Z(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G166), .B2(new_n705), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT91), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n793), .B1(new_n797), .B2(G1971), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n788), .B(new_n798), .C1(G1971), .C2(new_n797), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n801));
  OR2_X1    g376(.A1(G16), .A2(G24), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G290), .B2(new_n705), .ZN(new_n803));
  INV_X1    g378(.A(G1986), .ZN(new_n804));
  OAI21_X1  g379(.A(KEYINPUT92), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n712), .A2(G25), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT86), .Z(new_n807));
  NAND2_X1  g382(.A1(new_n469), .A2(G131), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT87), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(new_n483), .B2(G107), .ZN(new_n810));
  OR3_X1    g385(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n811));
  OAI21_X1  g386(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n484), .B2(G119), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n807), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT89), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n805), .B(new_n819), .C1(new_n804), .C2(new_n803), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n800), .A2(new_n801), .A3(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n822), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n784), .A2(new_n823), .A3(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  AOI22_X1  g401(.A1(G55), .A2(new_n536), .B1(new_n538), .B2(G93), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n526), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n612), .A2(G559), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n562), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g409(.A(KEYINPUT102), .B(new_n556), .C1(new_n560), .C2(new_n561), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n829), .A3(new_n835), .ZN(new_n836));
  OR3_X1    g411(.A1(new_n562), .A2(new_n829), .A3(new_n833), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n838));
  AND3_X1   g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n832), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n837), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(KEYINPUT38), .ZN(new_n843));
  INV_X1    g418(.A(new_n832), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n846), .A3(KEYINPUT39), .ZN(new_n847));
  INV_X1    g422(.A(G860), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n839), .A2(new_n840), .A3(new_n832), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT103), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(new_n850), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n849), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT104), .ZN(new_n859));
  AOI211_X1 g434(.A(new_n859), .B(new_n849), .C1(new_n854), .C2(new_n856), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n831), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g438(.A(KEYINPUT105), .B(new_n831), .C1(new_n858), .C2(new_n860), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(G145));
  XNOR2_X1  g440(.A(new_n815), .B(new_n630), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n469), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n484), .A2(G130), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(G2104), .C1(G118), .C2(new_n483), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n866), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT108), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n701), .B(new_n777), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n733), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n509), .A2(new_n497), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n469), .A2(new_n498), .B1(new_n496), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n500), .B1(new_n467), .B2(new_n468), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT106), .B1(new_n878), .B2(new_n507), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n502), .A2(new_n880), .A3(new_n508), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(KEYINPUT107), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n877), .A2(new_n879), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n875), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n873), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n638), .B(new_n480), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n488), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT109), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n888), .B2(new_n872), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n873), .B(new_n887), .ZN(new_n895));
  INV_X1    g470(.A(new_n891), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g473(.A1(new_n829), .A2(new_n622), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n608), .B(G299), .ZN(new_n900));
  XNOR2_X1  g475(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(KEYINPUT110), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n608), .A2(new_n616), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(KEYINPUT110), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n902), .B1(new_n905), .B2(KEYINPUT41), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n625), .B(new_n842), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n900), .B2(new_n907), .ZN(new_n909));
  XNOR2_X1  g484(.A(G303), .B(new_n790), .ZN(new_n910));
  XNOR2_X1  g485(.A(G305), .B(G290), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n910), .B(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT42), .Z(new_n913));
  XNOR2_X1  g488(.A(new_n909), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n899), .B1(new_n914), .B2(new_n622), .ZN(G295));
  OAI21_X1  g490(.A(new_n899), .B1(new_n914), .B2(new_n622), .ZN(G331));
  XNOR2_X1  g491(.A(G301), .B(G168), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n842), .B(new_n917), .Z(new_n918));
  AND3_X1   g493(.A1(new_n918), .A2(KEYINPUT41), .A3(new_n905), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n900), .B1(new_n918), .B2(new_n901), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n912), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n842), .B(new_n917), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n900), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n906), .B2(new_n922), .ZN(new_n924));
  INV_X1    g499(.A(new_n912), .ZN(new_n925));
  AOI21_X1  g500(.A(G37), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n924), .A2(new_n925), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT43), .B1(new_n930), .B2(new_n926), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT44), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n928), .B1(new_n930), .B2(new_n926), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n932), .A2(new_n936), .ZN(G397));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n883), .A2(new_n938), .A3(new_n885), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n470), .A2(G40), .A3(new_n479), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT112), .B1(G290), .B2(G1986), .ZN(new_n944));
  NAND2_X1  g519(.A1(G290), .A2(G1986), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n944), .B(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n817), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n815), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G2067), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n733), .B(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1996), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n777), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n809), .A2(new_n814), .A3(new_n817), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n948), .A2(new_n950), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n943), .B1(new_n946), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT123), .ZN(new_n956));
  NAND2_X1  g531(.A1(G286), .A2(G8), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1966), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT45), .B1(new_n882), .B2(new_n938), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n938), .ZN(new_n962));
  INV_X1    g537(.A(new_n942), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n511), .A2(new_n938), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n942), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n882), .A2(new_n968), .A3(new_n938), .ZN(new_n969));
  XOR2_X1   g544(.A(KEYINPUT116), .B(G2084), .Z(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n959), .B1(new_n972), .B2(G8), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n965), .A2(KEYINPUT122), .A3(new_n971), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT122), .B1(new_n965), .B2(new_n971), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n975), .A2(new_n976), .A3(G286), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n958), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n974), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT122), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n972), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n965), .A2(KEYINPUT122), .A3(new_n971), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n957), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n956), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(G168), .A3(new_n984), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n973), .B1(new_n988), .B2(new_n979), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n989), .A2(KEYINPUT123), .A3(new_n985), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT62), .B1(new_n987), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n981), .A2(new_n956), .A3(new_n986), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT123), .B1(new_n989), .B2(new_n985), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n938), .A4(new_n885), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n966), .A2(new_n940), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n963), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1971), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n967), .A2(new_n969), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(G2090), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n978), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT114), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1002), .B1(new_n998), .B2(new_n999), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  NOR4_X1   g586(.A1(new_n1010), .A2(new_n1007), .A3(new_n1011), .A4(new_n978), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n590), .A2(new_n1015), .A3(new_n592), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1015), .B1(new_n590), .B2(new_n592), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1018), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n882), .A2(new_n938), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(new_n942), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(new_n978), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n790), .A2(G1976), .ZN(new_n1027));
  INV_X1    g602(.A(G1976), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n583), .A2(new_n1028), .A3(new_n585), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1026), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n963), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(KEYINPUT50), .B2(new_n1022), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n998), .A2(new_n999), .B1(new_n1035), .B2(new_n722), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1007), .B1(new_n1036), .B2(new_n978), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n996), .A2(new_n744), .A3(new_n963), .A4(new_n997), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT124), .B(G1961), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1001), .A2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n961), .A2(new_n964), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1040), .A2(G2078), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(G171), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1013), .A2(new_n1038), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n991), .A2(new_n995), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT127), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT127), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n991), .A2(new_n1050), .A3(new_n1053), .A4(new_n995), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n978), .B(G286), .C1(new_n965), .C2(new_n971), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1033), .B(new_n1055), .C1(new_n1004), .C2(new_n1008), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(KEYINPUT63), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1024), .B(KEYINPUT115), .Z(new_n1058));
  AND3_X1   g633(.A1(new_n1025), .A2(new_n1028), .A3(new_n586), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n1017), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1037), .A2(new_n1062), .A3(new_n1055), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1061), .B1(new_n1033), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1052), .A2(new_n1054), .A3(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n941), .A2(new_n963), .A3(new_n996), .A4(new_n1046), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1041), .A2(new_n1067), .A3(G301), .A4(new_n1044), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT54), .B1(new_n1049), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n992), .B2(new_n993), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1013), .A2(new_n1038), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT126), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1041), .A2(new_n1044), .A3(new_n1067), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G171), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT125), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(G171), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1048), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(G301), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1072), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1073), .A2(new_n1076), .A3(G171), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1076), .B1(new_n1073), .B2(G171), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1081), .B(new_n1072), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1070), .B(new_n1071), .C1(new_n1082), .C2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT58), .B(G1341), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n998), .A2(G1996), .B1(new_n1023), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n563), .ZN(new_n1090));
  XOR2_X1   g665(.A(new_n1090), .B(KEYINPUT59), .Z(new_n1091));
  AOI21_X1  g666(.A(G1348), .B1(new_n967), .B2(new_n969), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1022), .A2(G2067), .A3(new_n942), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT60), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n624), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n612), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1096), .B1(new_n1095), .B2(new_n1097), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT60), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1100), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT60), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n1098), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1091), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1106));
  XNOR2_X1  g681(.A(G299), .B(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1107), .B(KEYINPUT119), .Z(new_n1108));
  XOR2_X1   g683(.A(KEYINPUT56), .B(G2072), .Z(new_n1109));
  OR2_X1    g684(.A1(new_n998), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1035), .A2(G1956), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1110), .B2(KEYINPUT118), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1110), .A2(KEYINPUT118), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1107), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(new_n1111), .A3(new_n1113), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1118), .A3(KEYINPUT61), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT120), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(new_n1118), .A3(new_n1121), .A4(KEYINPUT61), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1107), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1118), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1105), .A2(new_n1120), .A3(new_n1122), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1115), .A2(new_n1097), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1118), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1087), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n955), .B1(new_n1066), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n950), .A2(new_n952), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1132), .A2(new_n953), .B1(G2067), .B2(new_n733), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1133), .A2(new_n943), .ZN(new_n1134));
  INV_X1    g709(.A(new_n950), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n943), .B1(new_n777), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n943), .A2(new_n951), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1137), .A2(KEYINPUT46), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(KEYINPUT46), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT47), .Z(new_n1141));
  NOR2_X1   g716(.A1(G290), .A2(G1986), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n943), .A2(KEYINPUT48), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT48), .B1(new_n943), .B2(new_n1142), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1144), .B1(new_n943), .B2(new_n954), .ZN(new_n1145));
  AOI211_X1 g720(.A(new_n1134), .B(new_n1141), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1131), .A2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g722(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1149));
  OAI211_X1 g723(.A(new_n897), .B(new_n1149), .C1(new_n934), .C2(new_n935), .ZN(G225));
  INV_X1    g724(.A(G225), .ZN(G308));
endmodule


