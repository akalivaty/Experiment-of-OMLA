//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n440, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  AND2_X1   g014(.A1(KEYINPUT65), .A2(G57), .ZN(new_n440));
  NOR2_X1   g015(.A1(KEYINPUT65), .A2(G57), .ZN(new_n441));
  NOR2_X1   g016(.A1(new_n440), .A2(new_n441), .ZN(G237));
  XOR2_X1   g017(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n455), .A2(KEYINPUT67), .A3(G567), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n458), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n466), .B2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n468), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n475), .A2(new_n476), .A3(new_n465), .A4(new_n467), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT69), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(new_n473), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n472), .B1(new_n480), .B2(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G112), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT71), .Z(new_n492));
  AND4_X1   g067(.A1(G2105), .A2(new_n475), .A3(new_n467), .A4(new_n476), .ZN(new_n493));
  AOI211_X1 g068(.A(new_n486), .B(new_n492), .C1(G124), .C2(new_n493), .ZN(G162));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n493), .B2(G126), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n475), .A2(new_n476), .A3(new_n500), .A4(new_n467), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n467), .A2(new_n469), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n498), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  OR2_X1    g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n511), .A2(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n519), .A2(new_n520), .B1(G651), .B2(new_n524), .ZN(G166));
  INV_X1    g100(.A(new_n513), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g107(.A(new_n527), .B(new_n529), .C1(new_n532), .C2(KEYINPUT74), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n532), .A2(KEYINPUT74), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n513), .A2(new_n539), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n537), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n513), .A2(new_n545), .B1(new_n515), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  NAND2_X1  g128(.A1(new_n511), .A2(G65), .ZN(new_n554));
  INV_X1    g129(.A(G78), .ZN(new_n555));
  INV_X1    g130(.A(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OR3_X1    g132(.A1(new_n555), .A2(new_n556), .A3(KEYINPUT76), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n526), .A2(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n512), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(new_n565), .A3(G53), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n515), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(KEYINPUT75), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT75), .B1(new_n566), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n563), .B1(new_n570), .B2(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n524), .A2(G651), .ZN(new_n575));
  INV_X1    g150(.A(new_n520), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n576), .B2(new_n518), .ZN(G303));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(new_n515), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n511), .A2(new_n512), .A3(G87), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n582), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n564), .A2(G49), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT77), .A4(new_n579), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G288));
  NAND2_X1  g163(.A1(new_n511), .A2(G61), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n537), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n511), .A2(new_n512), .A3(G86), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n512), .A2(G48), .A3(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n564), .A2(G47), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT78), .B(G85), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n513), .B2(new_n598), .C1(new_n537), .C2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n511), .A2(new_n512), .A3(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n511), .A2(G66), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT79), .B1(new_n605), .B2(new_n556), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n605), .A2(new_n556), .A3(KEYINPUT79), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n564), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n603), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  XNOR2_X1  g187(.A(G321), .B(KEYINPUT80), .ZN(G284));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(new_n571), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n562), .B1(new_n615), .B2(new_n569), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n614), .B1(new_n616), .B2(G868), .ZN(G280));
  XNOR2_X1  g193(.A(KEYINPUT81), .B(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n611), .B1(G860), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g196(.A1(new_n611), .A2(new_n619), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g200(.A1(new_n465), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n628), .B1(KEYINPUT83), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n629), .A2(KEYINPUT83), .ZN(new_n631));
  MUX2_X1   g206(.A(new_n630), .B(new_n628), .S(new_n631), .Z(new_n632));
  NAND4_X1  g207(.A1(new_n475), .A2(new_n476), .A3(G2105), .A4(new_n467), .ZN(new_n633));
  INV_X1    g208(.A(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(KEYINPUT84), .B1(new_n465), .B2(G111), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(G2104), .A3(new_n636), .ZN(new_n637));
  NOR3_X1   g212(.A1(new_n465), .A2(KEYINPUT84), .A3(G111), .ZN(new_n638));
  OAI22_X1  g213(.A1(new_n633), .A2(new_n634), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n490), .B2(G135), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(G2096), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n632), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT85), .ZN(G156));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2427), .B(G2430), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n648), .B2(new_n649), .ZN(new_n652));
  XOR2_X1   g227(.A(G2443), .B(G2446), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(G14), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n656), .B2(new_n657), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT17), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2084), .B(G2090), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT87), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n665), .A2(new_n666), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n670), .B(new_n667), .C1(new_n664), .C2(new_n666), .ZN(new_n671));
  INV_X1    g246(.A(new_n667), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n664), .A3(new_n666), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n679), .A2(new_n680), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(new_n683), .A3(new_n681), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n686), .B(new_n688), .C1(new_n683), .C2(new_n687), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n696), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G2090), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G35), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G162), .B2(new_n701), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT29), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n611), .A2(G16), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G4), .B2(G16), .ZN(new_n708));
  INV_X1    g283(.A(G1348), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n712), .A2(G28), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n701), .B1(new_n712), .B2(G28), .ZN(new_n714));
  AND2_X1   g289(.A1(KEYINPUT31), .A2(G11), .ZN(new_n715));
  NOR2_X1   g290(.A1(KEYINPUT31), .A2(G11), .ZN(new_n716));
  OAI22_X1  g291(.A1(new_n713), .A2(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NOR2_X1   g293(.A1(G171), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G5), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1961), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n717), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n710), .A2(new_n711), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT25), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n727));
  INV_X1    g302(.A(G139), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n726), .B1(new_n465), .B2(new_n727), .C1(new_n489), .C2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G33), .B(new_n729), .S(G29), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2072), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n640), .A2(G29), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT98), .Z(new_n733));
  NOR3_X1   g308(.A1(new_n723), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G27), .A2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G164), .B2(G29), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(G2078), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G19), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n548), .B2(G16), .ZN(new_n739));
  OAI22_X1  g314(.A1(new_n720), .A2(new_n721), .B1(G1341), .B2(new_n739), .ZN(new_n740));
  AOI211_X1 g315(.A(new_n737), .B(new_n740), .C1(G1341), .C2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n718), .A2(G21), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G168), .B2(new_n718), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n743), .A2(G1966), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT99), .Z(new_n745));
  AOI22_X1  g320(.A1(new_n743), .A2(G1966), .B1(G2078), .B2(new_n736), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n734), .A2(new_n741), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n701), .A2(G26), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT94), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT28), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n493), .A2(G128), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n465), .A2(G116), .ZN(new_n752));
  OAI21_X1  g327(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n751), .B1(new_n752), .B2(new_n753), .C1(new_n489), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT95), .B(G2067), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G34), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n701), .B1(new_n759), .B2(G34), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(KEYINPUT96), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(KEYINPUT96), .B2(new_n761), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G160), .B2(G29), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n758), .B1(G2084), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT101), .B(KEYINPUT23), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n718), .A2(G20), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n616), .B2(new_n718), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n765), .B(new_n771), .C1(G2084), .C2(new_n764), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n706), .A2(new_n747), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G6), .A2(G16), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n595), .B2(G16), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT32), .B(G1981), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n718), .A2(G23), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n581), .A2(new_n582), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n779), .B2(new_n718), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT92), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n780), .B(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(G166), .A2(G16), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G16), .B2(G22), .ZN(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n777), .B(new_n783), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n490), .A2(G131), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n493), .A2(G119), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT90), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n465), .A2(G107), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n790), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT35), .B(G1991), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G16), .A2(G24), .ZN(new_n799));
  XNOR2_X1  g374(.A(G290), .B(KEYINPUT91), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G16), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G1986), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n797), .B2(new_n796), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n789), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT93), .B(KEYINPUT36), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n701), .A2(G32), .ZN(new_n807));
  NAND3_X1  g382(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT26), .Z(new_n809));
  NAND3_X1  g384(.A1(new_n465), .A2(G105), .A3(G2104), .ZN(new_n810));
  INV_X1    g385(.A(G129), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n633), .ZN(new_n812));
  INV_X1    g387(.A(G141), .ZN(new_n813));
  OR3_X1    g388(.A1(new_n489), .A2(KEYINPUT97), .A3(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT97), .B1(new_n489), .B2(new_n813), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n812), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n807), .B1(new_n816), .B2(new_n701), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT27), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1996), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT36), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(KEYINPUT93), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n789), .A2(new_n798), .A3(new_n803), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n773), .A2(new_n806), .A3(new_n819), .A4(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n704), .A2(new_n700), .A3(new_n705), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT100), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n825), .ZN(G311));
  XOR2_X1   g401(.A(new_n824), .B(KEYINPUT100), .Z(new_n827));
  AND2_X1   g402(.A1(new_n806), .A2(new_n822), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n827), .A2(new_n819), .A3(new_n773), .A4(new_n828), .ZN(G150));
  NAND2_X1  g404(.A1(new_n611), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n537), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  INV_X1    g409(.A(G55), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n513), .A2(new_n834), .B1(new_n515), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n548), .A2(new_n837), .ZN(new_n838));
  OAI22_X1  g413(.A1(new_n544), .A2(new_n547), .B1(new_n833), .B2(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n831), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  INV_X1    g418(.A(G860), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n837), .A2(new_n844), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n795), .B(new_n627), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n490), .A2(KEYINPUT103), .A3(G142), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  INV_X1    g428(.A(G142), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n489), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n857), .A2(KEYINPUT104), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(KEYINPUT104), .B2(new_n857), .ZN(new_n860));
  INV_X1    g435(.A(G130), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n633), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n729), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n816), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n816), .A2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n816), .A2(new_n865), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n856), .A2(new_n862), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n866), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n755), .B(G164), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n873), .B1(new_n869), .B2(new_n872), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n851), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(new_n872), .ZN(new_n878));
  INV_X1    g453(.A(new_n873), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n880), .A2(new_n850), .A3(new_n874), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n877), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n640), .B(G160), .Z(new_n884));
  XNOR2_X1  g459(.A(G162), .B(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(new_n885), .B2(new_n883), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g463(.A(new_n840), .B(KEYINPUT106), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n622), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n616), .A2(new_n610), .ZN(new_n891));
  NAND2_X1  g466(.A1(G299), .A2(new_n611), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(G299), .A2(new_n611), .A3(KEYINPUT107), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n891), .A2(new_n892), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n898), .B1(new_n890), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  XNOR2_X1  g482(.A(G303), .B(G290), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n779), .B(new_n595), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n906), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n906), .B2(new_n907), .ZN(new_n913));
  OAI21_X1  g488(.A(G868), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n837), .A2(G868), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(G295));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n915), .ZN(G331));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n840), .A2(G171), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n840), .A2(G171), .ZN(new_n921));
  AOI21_X1  g496(.A(G168), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n923), .A2(new_n919), .A3(G286), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n894), .A2(new_n901), .A3(new_n895), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n926), .A2(KEYINPUT108), .B1(KEYINPUT41), .B2(new_n900), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n926), .A2(KEYINPUT108), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n897), .B1(new_n924), .B2(new_n922), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n911), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n922), .A2(new_n924), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(new_n899), .A3(new_n902), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n910), .A3(new_n930), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n934), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n910), .B1(new_n936), .B2(new_n930), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT43), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n939), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n918), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n946), .B1(new_n947), .B2(new_n933), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(G397));
  XNOR2_X1  g525(.A(KEYINPUT116), .B(G8), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT115), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n507), .B2(new_n955), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n501), .A2(KEYINPUT4), .B1(new_n503), .B2(new_n504), .ZN(new_n957));
  INV_X1    g532(.A(new_n495), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G114), .B2(new_n465), .ZN(new_n959));
  INV_X1    g534(.A(G126), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n633), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n954), .B(new_n955), .C1(new_n957), .C2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n953), .B1(new_n956), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT119), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n955), .B1(new_n957), .B2(new_n961), .ZN(new_n966));
  XNOR2_X1  g541(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(new_n967), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n507), .A2(KEYINPUT119), .A3(new_n955), .A4(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G40), .ZN(new_n972));
  AOI211_X1 g547(.A(new_n972), .B(new_n472), .C1(new_n480), .C2(new_n482), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n964), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1966), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(KEYINPUT120), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n966), .A2(KEYINPUT115), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT50), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n978), .A3(new_n962), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n973), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2084), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n472), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n476), .A2(new_n467), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(G137), .A3(new_n465), .A4(new_n475), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n481), .B1(new_n988), .B2(new_n473), .ZN(new_n989));
  INV_X1    g564(.A(new_n482), .ZN(new_n990));
  OAI211_X1 g565(.A(G40), .B(new_n986), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n977), .A2(new_n962), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(new_n953), .ZN(new_n993));
  AOI21_X1  g568(.A(G1966), .B1(new_n993), .B2(new_n971), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(KEYINPUT120), .ZN(new_n995));
  OAI211_X1 g570(.A(G286), .B(new_n952), .C1(new_n985), .C2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n994), .A2(KEYINPUT120), .B1(new_n983), .B2(new_n982), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n974), .A2(new_n975), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT120), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n997), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G168), .A2(new_n951), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n996), .B(KEYINPUT51), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n952), .B1(new_n985), .B2(new_n995), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1003), .A2(KEYINPUT51), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(KEYINPUT62), .A3(new_n1007), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(G166), .B2(new_n997), .ZN(new_n1013));
  NAND3_X1  g588(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n966), .A2(new_n1016), .A3(new_n967), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n966), .B2(new_n967), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n955), .C1(new_n957), .C2(new_n961), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n991), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(G1971), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AND4_X1   g599(.A1(new_n700), .A2(new_n979), .A3(new_n973), .A4(new_n980), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1015), .B(G8), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(G1981), .B1(new_n591), .B2(new_n594), .ZN(new_n1027));
  INV_X1    g602(.A(G61), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n509), .B2(new_n510), .ZN(new_n1029));
  INV_X1    g604(.A(new_n590), .ZN(new_n1030));
  OAI21_X1  g605(.A(G651), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n592), .A4(new_n593), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1027), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT49), .B1(new_n1027), .B2(new_n1033), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n977), .A2(G160), .A3(G40), .A4(new_n962), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(new_n952), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1036), .A2(KEYINPUT117), .A3(new_n952), .A4(new_n1037), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n779), .A2(G1976), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n952), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT52), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n583), .A2(new_n586), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(new_n952), .A3(new_n1037), .A4(new_n1043), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1026), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G2078), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n966), .A2(new_n967), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT114), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1023), .A2(new_n1053), .A3(new_n1055), .A4(new_n1017), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n1057), .B1(new_n981), .B2(new_n721), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n993), .A2(KEYINPUT53), .A3(new_n1053), .A4(new_n971), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1015), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n978), .B1(new_n977), .B2(new_n962), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n978), .B(new_n955), .C1(new_n957), .C2(new_n961), .ZN(new_n1063));
  NAND3_X1  g638(.A1(G160), .A2(G40), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1055), .A2(new_n973), .A3(new_n1021), .A4(new_n1017), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1065), .A2(new_n700), .B1(new_n1066), .B2(new_n786), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1067), .B2(new_n951), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1052), .A2(new_n1060), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1010), .A2(new_n1011), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1023), .A2(new_n1055), .A3(new_n1017), .A4(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n770), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n566), .A2(new_n568), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n563), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1072), .A2(new_n1073), .A3(KEYINPUT123), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1076), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT124), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1076), .A2(new_n1085), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1037), .A2(KEYINPUT122), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n973), .A2(new_n1088), .A3(new_n977), .A4(new_n962), .ZN(new_n1089));
  AOI21_X1  g664(.A(G2067), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n991), .B1(KEYINPUT50), .B2(new_n966), .ZN(new_n1091));
  AOI21_X1  g666(.A(G1348), .B1(new_n1091), .B2(new_n979), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n611), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1084), .A2(new_n1086), .A3(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1072), .A2(new_n1073), .A3(new_n1077), .A4(new_n1080), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1074), .B2(new_n1081), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1098), .B2(KEYINPUT61), .ZN(new_n1099));
  NAND2_X1  g674(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g676(.A(KEYINPUT58), .B(G1341), .Z(new_n1102));
  NAND3_X1  g677(.A1(new_n1087), .A2(new_n1089), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1996), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1020), .A2(new_n1104), .A3(new_n1023), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n548), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT59), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1109), .A3(new_n548), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1090), .A2(new_n1092), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1112), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n611), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1100), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1113), .A2(new_n610), .B1(new_n1095), .B2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1101), .A2(new_n1111), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1096), .A2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1057), .B1(new_n1066), .B2(G2078), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n981), .A2(new_n721), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1023), .A2(KEYINPUT53), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(G171), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1058), .A2(G301), .A3(new_n1059), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT54), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(new_n1052), .A3(new_n1068), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1124), .A2(G171), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1060), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT126), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n1129), .C1(new_n1130), .C2(new_n1060), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1128), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1120), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1068), .A2(new_n1026), .A3(new_n1042), .A4(new_n1051), .ZN(new_n1139));
  OAI211_X1 g714(.A(G168), .B(new_n952), .C1(new_n985), .C2(new_n995), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT121), .B(new_n1138), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1144));
  OAI21_X1  g719(.A(G8), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1138), .B1(new_n1145), .B2(new_n1061), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1052), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1143), .B(new_n1144), .C1(new_n1140), .C2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1037), .A2(new_n952), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT118), .ZN(new_n1150));
  AOI211_X1 g725(.A(G1976), .B(G288), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1033), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1026), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1070), .A2(new_n1137), .A3(new_n1148), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1054), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n973), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT112), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n755), .B(G2067), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1159), .A2(G1996), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1160), .A2(new_n1161), .B1(new_n816), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1160), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n795), .B(new_n797), .Z(new_n1165));
  OR3_X1    g740(.A1(new_n1164), .A2(new_n1104), .A3(new_n816), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT113), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1169));
  OAI221_X1 g744(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1159), .A2(G1986), .A3(G290), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1159), .ZN(new_n1172));
  AND2_X1   g747(.A1(G290), .A2(G1986), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT111), .Z(new_n1175));
  NOR2_X1   g750(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1157), .A2(new_n1176), .ZN(new_n1177));
  XOR2_X1   g752(.A(new_n1162), .B(KEYINPUT46), .Z(new_n1178));
  NAND2_X1  g753(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1178), .B(new_n1179), .C1(new_n816), .C2(new_n1164), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT47), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1171), .B(KEYINPUT48), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1170), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n795), .A2(new_n797), .ZN(new_n1184));
  OAI211_X1 g759(.A(new_n1184), .B(new_n1163), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n755), .A2(G2067), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1164), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1177), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g764(.A1(G227), .A2(new_n463), .ZN(new_n1191));
  AOI21_X1  g765(.A(new_n1191), .B1(new_n697), .B2(new_n698), .ZN(new_n1192));
  OAI21_X1  g766(.A(new_n1192), .B1(new_n661), .B2(new_n662), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n1193), .A2(KEYINPUT127), .ZN(new_n1194));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n1195));
  OAI211_X1 g769(.A(new_n1192), .B(new_n1195), .C1(new_n661), .C2(new_n662), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n887), .B(new_n1197), .C1(new_n940), .C2(new_n944), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


