//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT68), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT66), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n207));
  NAND3_X1  g006(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(KEYINPUT25), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n218), .A2(KEYINPUT23), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n217), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n203), .B1(new_n214), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n212), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n226), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n228), .A2(new_n231), .A3(KEYINPUT64), .A4(new_n211), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  INV_X1    g032(.A(G176gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT23), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n235), .A2(new_n216), .A3(new_n219), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n227), .A2(new_n232), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n221), .A2(new_n222), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n213), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n240), .A2(new_n241), .A3(KEYINPUT68), .A4(new_n217), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  OR2_X1    g046(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(G113gat), .A3(new_n249), .ZN(new_n250));
  OR2_X1    g049(.A1(KEYINPUT74), .A2(G113gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT74), .A2(G113gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(G120gat), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n255), .A2(KEYINPUT72), .A3(G134gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n244), .B2(KEYINPUT72), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  INV_X1    g057(.A(G120gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT1), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n258), .B2(new_n259), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n247), .A2(new_n254), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n229), .A2(KEYINPUT27), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT27), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G183gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n265), .A3(new_n230), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n263), .A2(new_n265), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n270), .A2(KEYINPUT70), .A3(KEYINPUT28), .A4(new_n230), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n266), .B2(new_n267), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n266), .A2(new_n274), .A3(new_n267), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n269), .A2(new_n271), .A3(new_n273), .A4(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT26), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT71), .B(new_n219), .C1(new_n218), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n218), .A2(new_n277), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n219), .B1(new_n218), .B2(new_n277), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n280), .A2(new_n283), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n276), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n243), .A2(new_n262), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT75), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n243), .A2(new_n285), .A3(new_n288), .A4(new_n262), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n243), .A2(new_n285), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n247), .A2(new_n254), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n257), .A2(new_n261), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n287), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n202), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT33), .ZN(new_n299));
  XOR2_X1   g098(.A(G15gat), .B(G43gat), .Z(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT76), .ZN(new_n301));
  XNOR2_X1  g100(.A(G71gat), .B(G99gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n298), .B1(new_n299), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT33), .B1(new_n295), .B2(new_n297), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n306));
  NOR4_X1   g105(.A1(new_n298), .A2(new_n305), .A3(new_n306), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n295), .A2(new_n297), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n303), .B1(new_n308), .B2(KEYINPUT32), .ZN(new_n309));
  INV_X1    g108(.A(new_n305), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT77), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n304), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n287), .A2(new_n294), .A3(new_n296), .A4(new_n289), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314));
  OR3_X1    g113(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT34), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(KEYINPUT34), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n314), .B1(new_n313), .B2(KEYINPUT34), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT36), .ZN(new_n320));
  INV_X1    g119(.A(new_n318), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n321), .B(new_n304), .C1(new_n307), .C2(new_n311), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n320), .B1(new_n319), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT81), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n257), .A2(new_n261), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n246), .B1(new_n250), .B2(new_n253), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT81), .ZN(new_n330));
  XOR2_X1   g129(.A(G141gat), .B(G148gat), .Z(new_n331));
  INV_X1    g130(.A(G155gat), .ZN(new_n332));
  INV_X1    g131(.A(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT2), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G155gat), .B(G162gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n336), .A3(new_n334), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n329), .A2(new_n330), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n339), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n336), .B1(new_n331), .B2(new_n334), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n262), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G225gat), .A2(G233gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n347), .B(KEYINPUT82), .Z(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n342), .B2(new_n343), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n338), .A2(new_n351), .A3(new_n339), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n329), .A2(new_n350), .A3(new_n330), .A4(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n348), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n355), .B1(new_n344), .B2(new_n262), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n293), .A2(new_n340), .A3(KEYINPUT4), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n353), .B(new_n354), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n356), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n355), .A3(new_n262), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n364), .A2(new_n354), .A3(new_n353), .A4(new_n359), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT0), .ZN(new_n368));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT6), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n370), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n361), .A2(new_n372), .A3(new_n365), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n372), .B1(new_n361), .B2(new_n365), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT6), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n366), .A2(KEYINPUT6), .A3(new_n370), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT84), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n374), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(G64gat), .B(G92gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  INV_X1    g182(.A(G226gat), .ZN(new_n384));
  INV_X1    g183(.A(G233gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(KEYINPUT29), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n290), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n243), .B(new_n285), .C1(new_n384), .C2(new_n385), .ZN(new_n390));
  XNOR2_X1  g189(.A(G211gat), .B(G218gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G197gat), .B(G204gat), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT79), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(KEYINPUT79), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n392), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n399), .A2(new_n391), .A3(new_n395), .A4(new_n393), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n389), .A2(new_n390), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT80), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT80), .B1(new_n398), .B2(new_n400), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n389), .B2(new_n390), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n383), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n408), .ZN(new_n410));
  INV_X1    g209(.A(new_n383), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n403), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT30), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n383), .C1(new_n404), .C2(new_n408), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT29), .B1(new_n398), .B2(new_n400), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n417), .A2(KEYINPUT86), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n351), .B1(new_n417), .B2(KEYINPUT86), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n340), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G228gat), .A2(G233gat), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n352), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n407), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n398), .A2(new_n400), .A3(KEYINPUT85), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n427), .B(new_n392), .C1(new_n396), .C2(new_n397), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n344), .B1(new_n429), .B2(new_n351), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n423), .A2(new_n402), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n421), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G22gat), .ZN(new_n435));
  INV_X1    g234(.A(G22gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n425), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT88), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT31), .B(G50gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n439), .B1(new_n441), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n444), .ZN(new_n446));
  AOI211_X1 g245(.A(KEYINPUT88), .B(new_n446), .C1(new_n437), .C2(new_n440), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n438), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n428), .A2(new_n422), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT3), .B1(new_n449), .B2(new_n426), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n431), .B1(new_n450), .B2(new_n344), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n421), .A2(new_n451), .B1(new_n420), .B2(new_n424), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT87), .B1(new_n452), .B2(new_n436), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT88), .B1(new_n453), .B2(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(new_n438), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n441), .A2(new_n439), .A3(new_n444), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n380), .A2(new_n416), .B1(new_n448), .B2(new_n457), .ZN(new_n458));
  AND4_X1   g257(.A1(new_n376), .A2(new_n366), .A3(KEYINPUT6), .A4(new_n370), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n376), .B1(new_n375), .B2(KEYINPUT6), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT92), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n379), .A2(new_n462), .A3(new_n377), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n371), .A2(KEYINPUT89), .A3(new_n373), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT89), .B1(new_n371), .B2(new_n373), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT37), .B1(new_n410), .B2(new_n403), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(new_n383), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n410), .A2(KEYINPUT37), .A3(new_n403), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT38), .ZN(new_n472));
  INV_X1    g271(.A(new_n409), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n401), .B1(new_n389), .B2(new_n390), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(KEYINPUT91), .ZN(new_n475));
  INV_X1    g274(.A(new_n407), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n389), .A2(new_n390), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT90), .ZN(new_n478));
  OR2_X1    g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n478), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n474), .A2(KEYINPUT91), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n475), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n468), .A2(KEYINPUT38), .A3(new_n383), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n473), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n464), .A2(new_n467), .A3(new_n472), .A4(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n354), .B1(new_n364), .B2(new_n353), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n370), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n341), .A2(new_n354), .A3(new_n345), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n329), .A2(new_n330), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n350), .A2(new_n352), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n491), .A2(new_n492), .B1(new_n362), .B2(new_n363), .ZN(new_n493));
  OAI211_X1 g292(.A(KEYINPUT39), .B(new_n490), .C1(new_n493), .C2(new_n354), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT40), .B1(new_n489), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(new_n375), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n494), .A3(KEYINPUT40), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n496), .A2(new_n415), .A3(new_n413), .A4(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n498), .A2(new_n457), .A3(new_n448), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n458), .B1(new_n486), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n448), .A2(new_n457), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n459), .A2(new_n460), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n502), .A2(new_n374), .B1(new_n415), .B2(new_n413), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n319), .A2(new_n501), .A3(new_n503), .A4(new_n322), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT35), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n416), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n464), .B2(new_n467), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n508), .A2(new_n319), .A3(new_n322), .A4(new_n501), .ZN(new_n509));
  AOI22_X1  g308(.A1(new_n325), .A2(new_n500), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(G29gat), .A2(G36gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n513), .B(KEYINPUT14), .Z(new_n514));
  XNOR2_X1  g313(.A(KEYINPUT94), .B(G29gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT95), .B(G36gat), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  XOR2_X1   g316(.A(G43gat), .B(G50gat), .Z(new_n518));
  INV_X1    g317(.A(KEYINPUT15), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(KEYINPUT96), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(new_n517), .B2(new_n520), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n518), .B(new_n519), .ZN(new_n525));
  OAI22_X1  g324(.A1(new_n522), .A2(new_n524), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G15gat), .B(G22gat), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT16), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(G1gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G1gat), .B2(new_n528), .ZN(new_n531));
  INV_X1    g330(.A(G8gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n526), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT97), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n533), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(new_n527), .B2(KEYINPUT17), .ZN(new_n540));
  AOI211_X1 g339(.A(new_n512), .B(new_n534), .C1(new_n538), .C2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT98), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT18), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n538), .A2(new_n540), .ZN(new_n544));
  INV_X1    g343(.A(new_n534), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n511), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT98), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n544), .A2(new_n511), .A3(new_n545), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n527), .A2(new_n533), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n534), .B1(KEYINPUT99), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(KEYINPUT99), .B2(new_n551), .ZN(new_n553));
  XOR2_X1   g352(.A(new_n511), .B(KEYINPUT13), .Z(new_n554));
  AOI22_X1  g353(.A1(new_n549), .A2(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(G113gat), .B(G141gat), .Z(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G169gat), .B(G197gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT12), .Z(new_n561));
  AND3_X1   g360(.A1(new_n548), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n561), .B1(new_n548), .B2(new_n555), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n510), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G230gat), .A2(G233gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G85gat), .A2(G92gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT7), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  INV_X1    g369(.A(G85gat), .ZN(new_n571));
  INV_X1    g370(.A(G92gat), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G99gat), .B(G106gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT101), .ZN(new_n577));
  XOR2_X1   g376(.A(G57gat), .B(G64gat), .Z(new_n578));
  INV_X1    g377(.A(KEYINPUT9), .ZN(new_n579));
  INV_X1    g378(.A(G71gat), .ZN(new_n580));
  INV_X1    g379(.A(G78gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584));
  OR2_X1    g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT100), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n577), .A2(KEYINPUT10), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n576), .B(new_n587), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n567), .B1(new_n594), .B2(KEYINPUT102), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(KEYINPUT102), .B2(new_n594), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n591), .A2(new_n566), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(KEYINPUT103), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n594), .A2(new_n566), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n605), .B1(new_n607), .B2(new_n598), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n577), .B1(new_n527), .B2(KEYINPUT17), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n538), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n577), .A2(new_n526), .B1(KEYINPUT41), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G190gat), .B(G218gat), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n614), .A2(KEYINPUT41), .ZN(new_n619));
  XNOR2_X1  g418(.A(G134gat), .B(G162gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n612), .A2(new_n622), .A3(new_n615), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n618), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n618), .B2(new_n623), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT21), .B1(new_n585), .B2(new_n586), .ZN(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n255), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n539), .B1(new_n589), .B2(KEYINPUT21), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G155gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g435(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n632), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n626), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n565), .A2(new_n610), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n380), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  INV_X1    g447(.A(new_n416), .ZN(new_n649));
  XOR2_X1   g448(.A(KEYINPUT16), .B(G8gat), .Z(new_n650));
  AND3_X1   g449(.A1(new_n645), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n532), .B1(new_n645), .B2(new_n649), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(KEYINPUT42), .B2(new_n651), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n319), .A2(new_n322), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n645), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n325), .B1(new_n643), .B2(new_n644), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n659), .B2(new_n655), .ZN(G1326gat));
  INV_X1    g459(.A(new_n501), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT43), .B(G22gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  INV_X1    g463(.A(new_n626), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(new_n609), .A3(new_n639), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n565), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n646), .A3(new_n515), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT45), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n510), .B2(new_n665), .ZN(new_n671));
  INV_X1    g470(.A(new_n324), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n500), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n661), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n675), .A2(new_n508), .B1(new_n504), .B2(KEYINPUT35), .ZN(new_n676));
  OAI211_X1 g475(.A(KEYINPUT44), .B(new_n626), .C1(new_n674), .C2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n639), .B(KEYINPUT105), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n609), .B(KEYINPUT106), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n564), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n380), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n669), .B1(new_n515), .B2(new_n684), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n667), .A2(new_n649), .A3(new_n516), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT46), .Z(new_n687));
  NOR2_X1   g486(.A1(new_n683), .A2(new_n416), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n516), .B2(new_n688), .ZN(G1329gat));
  NAND2_X1  g488(.A1(new_n667), .A2(new_n657), .ZN(new_n690));
  INV_X1    g489(.A(G43gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n693));
  INV_X1    g492(.A(new_n325), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G43gat), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n692), .B(new_n693), .C1(new_n683), .C2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n696), .A2(KEYINPUT108), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n692), .B1(new_n683), .B2(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT47), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n698), .B2(new_n700), .ZN(G1330gat));
  INV_X1    g500(.A(G50gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n667), .A2(new_n702), .A3(new_n661), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT48), .B1(new_n703), .B2(KEYINPUT111), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(KEYINPUT111), .B2(new_n703), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n678), .A2(new_n661), .A3(new_n682), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(G50gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n703), .B(KEYINPUT110), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(G50gat), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(G1331gat));
  NAND2_X1  g511(.A1(new_n564), .A2(new_n641), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n510), .A2(new_n713), .A3(new_n680), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n646), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g515(.A(new_n416), .B(KEYINPUT112), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT113), .B(KEYINPUT114), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1333gat));
  AOI21_X1  g522(.A(new_n580), .B1(new_n714), .B2(new_n694), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n656), .A2(G71gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n714), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n714), .A2(new_n661), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT116), .B(new_n626), .C1(new_n674), .C2(new_n676), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n564), .A2(new_n640), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n325), .A2(new_n500), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n505), .A2(new_n509), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n665), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(KEYINPUT116), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n730), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT116), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n510), .B2(new_n665), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n741), .A2(new_n731), .A3(KEYINPUT51), .A4(new_n733), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n646), .A2(new_n571), .A3(new_n609), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n732), .A2(new_n610), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n671), .A2(new_n677), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n671), .A2(new_n677), .A3(KEYINPUT115), .A4(new_n746), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n749), .A2(new_n646), .A3(new_n750), .ZN(new_n751));
  OAI22_X1  g550(.A1(new_n744), .A2(new_n745), .B1(new_n751), .B2(new_n571), .ZN(G1336gat));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n749), .A2(new_n649), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n680), .A2(G92gat), .A3(new_n717), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n743), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n756), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n739), .B2(new_n742), .ZN(new_n760));
  OAI21_X1  g559(.A(G92gat), .B1(new_n747), .B2(new_n717), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n753), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT117), .B1(new_n758), .B2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n757), .A2(new_n753), .A3(new_n761), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n760), .B1(G92gat), .B2(new_n754), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n765), .B(new_n766), .C1(new_n767), .C2(new_n753), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n764), .A2(new_n768), .ZN(G1337gat));
  INV_X1    g568(.A(G99gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n657), .A2(new_n770), .A3(new_n609), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n749), .A2(new_n694), .A3(new_n750), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n744), .A2(new_n771), .B1(new_n772), .B2(new_n770), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n680), .A2(G106gat), .A3(new_n501), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n743), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G106gat), .B1(new_n747), .B2(new_n501), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n777));
  NAND3_X1  g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n749), .A2(new_n661), .A3(new_n750), .ZN(new_n779));
  AOI22_X1  g578(.A1(G106gat), .A2(new_n779), .B1(new_n743), .B2(new_n774), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(G1339gat));
  INV_X1    g581(.A(new_n679), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n602), .B1(new_n606), .B2(KEYINPUT54), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n590), .A2(new_n593), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(new_n567), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n596), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n604), .B1(new_n788), .B2(KEYINPUT55), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT102), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n566), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n594), .A2(KEYINPUT102), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n784), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT119), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n788), .A2(new_n798), .A3(KEYINPUT55), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n789), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n562), .B2(new_n563), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n548), .A2(new_n555), .A3(new_n561), .ZN(new_n802));
  INV_X1    g601(.A(new_n560), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n553), .A2(new_n554), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n511), .B1(new_n544), .B2(new_n545), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(new_n609), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n626), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n800), .A2(new_n802), .A3(new_n626), .A4(new_n806), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n783), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n713), .A2(new_n609), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n814), .A2(new_n646), .A3(new_n675), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n717), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n564), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(G113gat), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n251), .A2(new_n252), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n817), .ZN(G1340gat));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821));
  OAI21_X1  g620(.A(G120gat), .B1(new_n816), .B2(new_n680), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n609), .A2(new_n248), .A3(new_n249), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n821), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n822), .B(KEYINPUT120), .C1(new_n816), .C2(new_n824), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1341gat));
  OAI21_X1  g627(.A(G127gat), .B1(new_n816), .B2(new_n783), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n639), .A2(new_n255), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n816), .B2(new_n830), .ZN(G1342gat));
  INV_X1    g630(.A(G134gat), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n665), .A2(new_n649), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n815), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  XOR2_X1   g633(.A(new_n834), .B(KEYINPUT56), .Z(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n816), .B2(new_n665), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1343gat));
  NOR2_X1   g636(.A1(new_n694), .A2(new_n380), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n814), .A2(new_n661), .A3(new_n717), .A4(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n564), .ZN(new_n840));
  INV_X1    g639(.A(G141gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(KEYINPUT58), .B1(new_n843), .B2(KEYINPUT122), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n717), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n694), .A2(new_n380), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n501), .A2(new_n849), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n795), .A2(new_n796), .B1(new_n596), .B2(new_n603), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n798), .B1(new_n788), .B2(KEYINPUT55), .ZN(new_n852));
  AND4_X1   g651(.A1(new_n798), .A2(new_n793), .A3(KEYINPUT55), .A4(new_n794), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n542), .B1(new_n541), .B2(KEYINPUT18), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n546), .A2(KEYINPUT98), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n555), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n561), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n854), .B1(new_n859), .B2(new_n802), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n802), .A2(new_n609), .A3(new_n806), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n665), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n639), .B1(new_n862), .B2(new_n809), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n813), .B1(new_n863), .B2(KEYINPUT121), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT121), .B(new_n640), .C1(new_n808), .C2(new_n810), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n850), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n809), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n812), .B1(new_n868), .B2(new_n783), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n849), .B1(new_n869), .B2(new_n501), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n848), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n841), .B1(new_n871), .B2(new_n840), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n845), .B1(new_n872), .B2(new_n843), .ZN(new_n873));
  INV_X1    g672(.A(new_n850), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n640), .B1(new_n808), .B2(new_n810), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n812), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n874), .B1(new_n877), .B2(new_n865), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT57), .B1(new_n814), .B2(new_n661), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n847), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(G141gat), .B1(new_n880), .B2(new_n564), .ZN(new_n881));
  INV_X1    g680(.A(new_n843), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n844), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n873), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(new_n839), .ZN(new_n885));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n609), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n847), .A2(new_n609), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n661), .B1(new_n863), .B2(new_n812), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n849), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n814), .A2(new_n850), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n886), .B1(new_n893), .B2(KEYINPUT123), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n890), .A2(new_n849), .B1(new_n814), .B2(new_n850), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n889), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n888), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n888), .A2(G148gat), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n871), .B2(new_n609), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n887), .B1(new_n898), .B2(new_n900), .ZN(G1345gat));
  OAI21_X1  g700(.A(G155gat), .B1(new_n880), .B2(new_n783), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n332), .A3(new_n639), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n880), .B2(new_n665), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n814), .A2(new_n661), .A3(new_n838), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n833), .A2(new_n333), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(G1347gat));
  NAND4_X1  g707(.A1(new_n814), .A2(new_n380), .A3(new_n649), .A4(new_n675), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n233), .A3(new_n564), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n869), .A2(new_n646), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(new_n675), .A3(new_n846), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n840), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n910), .B1(new_n913), .B2(new_n233), .ZN(G1348gat));
  NAND3_X1  g713(.A1(new_n912), .A2(new_n234), .A3(new_n609), .ZN(new_n915));
  OAI21_X1  g714(.A(G176gat), .B1(new_n909), .B2(new_n680), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1349gat));
  NOR2_X1   g716(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n918));
  OAI21_X1  g717(.A(G183gat), .B1(new_n909), .B2(new_n783), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n639), .A2(new_n270), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n911), .A2(new_n675), .A3(new_n846), .A4(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n912), .A2(new_n230), .A3(new_n626), .ZN(new_n925));
  OAI21_X1  g724(.A(G190gat), .B1(new_n909), .B2(new_n665), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n926), .A2(KEYINPUT61), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n926), .A2(KEYINPUT61), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(G1351gat));
  NOR3_X1   g728(.A1(new_n694), .A2(new_n717), .A3(new_n501), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n564), .A2(G197gat), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n911), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n325), .A2(new_n380), .A3(new_n649), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n875), .A2(new_n813), .ZN(new_n935));
  AOI21_X1  g734(.A(KEYINPUT57), .B1(new_n935), .B2(new_n661), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n869), .A2(new_n874), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n840), .B(new_n934), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n932), .B1(new_n938), .B2(G197gat), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT126), .ZN(G1352gat));
  NAND2_X1  g739(.A1(new_n911), .A2(new_n930), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n941), .A2(G204gat), .A3(new_n610), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n891), .A2(new_n892), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n681), .A3(new_n934), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G204gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n946), .ZN(G1353gat));
  INV_X1    g746(.A(G211gat), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n640), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(KEYINPUT63), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n639), .A2(new_n948), .ZN(new_n953));
  OAI22_X1  g752(.A1(new_n951), .A2(new_n952), .B1(new_n941), .B2(new_n953), .ZN(G1354gat));
  INV_X1    g753(.A(new_n934), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT127), .B1(new_n896), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n626), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n896), .A2(KEYINPUT127), .A3(new_n955), .ZN(new_n958));
  OAI21_X1  g757(.A(G218gat), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n665), .A2(G218gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n941), .B2(new_n960), .ZN(G1355gat));
endmodule


