//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n467), .B1(new_n472), .B2(new_n466), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n464), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(KEYINPUT69), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(new_n464), .C1(new_n471), .C2(new_n473), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n461), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n472), .A2(new_n461), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n472), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n461), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n485), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT70), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n495));
  OAI211_X1 g070(.A(G126), .B(G2105), .C1(new_n469), .C2(new_n468), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n469), .A2(new_n468), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n461), .A2(KEYINPUT71), .A3(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT4), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n499), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n472), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n500), .B2(new_n503), .ZN(G164));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G50), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n512), .A2(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  INV_X1    g092(.A(G88), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n510), .B1(new_n521), .B2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n514), .A2(KEYINPUT73), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n531), .B(new_n533), .C1(new_n517), .C2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n528), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n539), .A2(new_n509), .B1(new_n517), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n529), .A2(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n507), .A2(G56), .ZN(new_n544));
  INV_X1    g119(.A(G68), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n545), .B2(new_n511), .ZN(new_n546));
  INV_X1    g121(.A(new_n517), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n546), .A2(G651), .B1(new_n547), .B2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT74), .ZN(G188));
  NAND2_X1  g131(.A1(new_n514), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n547), .A2(G91), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OAI211_X1 g135(.A(new_n558), .B(new_n559), .C1(new_n509), .C2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT75), .ZN(G299));
  INV_X1    g137(.A(G171), .ZN(G301));
  INV_X1    g138(.A(G168), .ZN(G286));
  OAI21_X1  g139(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  INV_X1    g141(.A(G49), .ZN(new_n567));
  INV_X1    g142(.A(new_n514), .ZN(new_n568));
  OAI221_X1 g143(.A(new_n565), .B1(new_n517), .B2(new_n566), .C1(new_n567), .C2(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n514), .A2(G48), .ZN(new_n570));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n517), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n507), .A2(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n509), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n573), .A2(new_n577), .ZN(G305));
  XNOR2_X1  g153(.A(KEYINPUT76), .B(G47), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n528), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n509), .B1(new_n517), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n547), .A2(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT10), .Z(new_n588));
  NAND2_X1  g163(.A1(new_n529), .A2(G54), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(new_n509), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n586), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n586), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n561), .B(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n595), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n592), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n484), .A2(G135), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n487), .A2(G123), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n461), .A2(G111), .ZN(new_n608));
  OAI21_X1  g183(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n606), .B(new_n607), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT77), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(G2096), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n472), .A2(new_n463), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(G156));
  XOR2_X1   g192(.A(G1341), .B(G1348), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT79), .ZN(new_n619));
  XOR2_X1   g194(.A(G2451), .B(G2454), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n619), .B(new_n621), .Z(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT78), .B(KEYINPUT14), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT15), .B(G2435), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  AOI21_X1  g201(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n625), .B2(new_n626), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n622), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2443), .B(G2446), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  AND3_X1   g207(.A1(new_n631), .A2(G14), .A3(new_n632), .ZN(G401));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  XOR2_X1   g209(.A(G2072), .B(G2078), .Z(new_n635));
  XOR2_X1   g210(.A(KEYINPUT81), .B(KEYINPUT17), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT80), .Z(new_n640));
  AOI21_X1  g215(.A(new_n634), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n635), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(new_n640), .ZN(new_n643));
  INV_X1    g218(.A(new_n634), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n639), .A3(new_n634), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n647), .A2(KEYINPUT18), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n647), .A2(KEYINPUT18), .ZN(new_n649));
  OAI221_X1 g224(.A(new_n643), .B1(new_n638), .B2(new_n645), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2096), .B(G2100), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1961), .B(G1966), .Z(new_n657));
  AND2_X1   g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT20), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n656), .A2(new_n657), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n654), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n654), .B2(new_n661), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT82), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT83), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  MUX2_X1   g247(.A(G6), .B(G305), .S(G16), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT85), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT32), .B(G1981), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(G16), .A2(G22), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G166), .B2(G16), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G23), .ZN(new_n682));
  INV_X1    g257(.A(G288), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT33), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1976), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n676), .A2(new_n680), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n681), .A2(G24), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n584), .B2(new_n681), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1986), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(G25), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n484), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n487), .A2(G119), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n461), .A2(G107), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT84), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(G29), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT35), .B(G1991), .Z(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n692), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n688), .A2(new_n689), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT36), .Z(new_n707));
  NOR2_X1   g282(.A1(G29), .A2(G35), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G162), .B2(G29), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G2090), .ZN(new_n711));
  OAI21_X1  g286(.A(KEYINPUT92), .B1(G29), .B2(G32), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n463), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT26), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n487), .B2(G129), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n717), .A2(new_n693), .ZN(new_n718));
  MUX2_X1   g293(.A(new_n712), .B(KEYINPUT92), .S(new_n718), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT27), .B(G1996), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(KEYINPUT93), .B1(G16), .B2(G21), .ZN(new_n722));
  NOR2_X1   g297(.A1(G286), .A2(new_n681), .ZN(new_n723));
  MUX2_X1   g298(.A(new_n722), .B(KEYINPUT93), .S(new_n723), .Z(new_n724));
  INV_X1    g299(.A(G1966), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AOI211_X1 g301(.A(new_n711), .B(new_n726), .C1(new_n725), .C2(new_n724), .ZN(new_n727));
  NAND2_X1  g302(.A1(G160), .A2(G29), .ZN(new_n728));
  INV_X1    g303(.A(G34), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(KEYINPUT24), .ZN(new_n730));
  AOI21_X1  g305(.A(G29), .B1(new_n729), .B2(KEYINPUT24), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(KEYINPUT89), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(KEYINPUT89), .B2(new_n731), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT90), .Z(new_n734));
  NAND3_X1  g309(.A1(new_n728), .A2(KEYINPUT91), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n735), .B1(KEYINPUT94), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(KEYINPUT91), .B1(new_n728), .B2(new_n734), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(G4), .A2(G16), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n592), .B2(G16), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT86), .B(G1348), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n693), .A2(G26), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT88), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  AOI22_X1  g323(.A1(G128), .A2(new_n487), .B1(new_n484), .B2(G140), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G116), .B2(new_n461), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT87), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n693), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n693), .A2(G33), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT25), .ZN(new_n759));
  NAND2_X1  g334(.A1(G103), .A2(G2104), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n760), .B2(G2105), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n484), .A2(G139), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n461), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n758), .B1(new_n765), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2072), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT30), .B(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n769), .A2(new_n693), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n610), .B2(new_n693), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n766), .B2(new_n767), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n693), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n693), .ZN(new_n776));
  INV_X1    g351(.A(G2078), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n757), .A2(new_n768), .A3(new_n774), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n681), .A2(G19), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n550), .B2(new_n681), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n681), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n681), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1961), .ZN(new_n785));
  NOR4_X1   g360(.A1(new_n745), .A2(new_n779), .A3(new_n782), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n681), .A2(G20), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT95), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT23), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n597), .B2(new_n681), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n710), .B2(G2090), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n727), .A2(new_n741), .A3(new_n786), .A4(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n707), .A2(new_n793), .ZN(G311));
  INV_X1    g369(.A(G311), .ZN(G150));
  NAND2_X1  g370(.A1(new_n592), .A2(G559), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT38), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n529), .A2(G55), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  INV_X1    g374(.A(G93), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n799), .A2(new_n509), .B1(new_n517), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(new_n550), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n549), .B1(new_n798), .B2(new_n801), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n797), .B(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT39), .ZN(new_n808));
  INV_X1    g383(.A(G860), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(KEYINPUT39), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n802), .A2(new_n809), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(G145));
  INV_X1    g389(.A(G37), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n498), .A2(KEYINPUT4), .A3(new_n499), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n502), .B1(new_n472), .B2(new_n501), .ZN(new_n817));
  OAI21_X1  g392(.A(KEYINPUT96), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n495), .A2(new_n496), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n497), .A2(KEYINPUT97), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n500), .A2(new_n503), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n818), .A2(new_n821), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n754), .B(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(G130), .A2(new_n487), .B1(new_n484), .B2(G142), .ZN(new_n827));
  NOR3_X1   g402(.A1(new_n461), .A2(KEYINPUT98), .A3(G118), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT98), .B1(new_n461), .B2(G118), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n826), .B(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n699), .B(new_n614), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n765), .B(new_n717), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n832), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(G160), .B(new_n610), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n492), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n815), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n837), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g417(.A(G305), .B(KEYINPUT100), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G290), .ZN(new_n844));
  XNOR2_X1  g419(.A(G303), .B(new_n683), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT42), .Z(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  NAND2_X1  g423(.A1(G299), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n597), .A2(KEYINPUT99), .ZN(new_n850));
  INV_X1    g425(.A(new_n592), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n597), .A2(KEYINPUT99), .A3(new_n592), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n805), .B(new_n602), .Z(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n853), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n852), .A2(KEYINPUT41), .A3(new_n853), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n856), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n847), .B(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G868), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(G868), .B2(new_n802), .ZN(G295));
  OAI21_X1  g440(.A(new_n864), .B1(G868), .B2(new_n802), .ZN(G331));
  INV_X1    g441(.A(KEYINPUT101), .ZN(new_n867));
  XNOR2_X1  g442(.A(G171), .B(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(G286), .ZN(new_n869));
  XNOR2_X1  g444(.A(G171), .B(KEYINPUT101), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(G168), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n805), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(G168), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n868), .A2(G286), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n806), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n859), .A2(new_n860), .A3(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(KEYINPUT102), .B(new_n805), .C1(new_n869), .C2(new_n871), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n879), .A2(new_n854), .A3(new_n880), .A4(new_n875), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n877), .A2(new_n881), .A3(KEYINPUT103), .ZN(new_n882));
  AOI21_X1  g457(.A(KEYINPUT103), .B1(new_n877), .B2(new_n881), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n882), .A2(new_n883), .A3(new_n846), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n877), .A2(new_n881), .ZN(new_n885));
  INV_X1    g460(.A(new_n846), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n815), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n889));
  INV_X1    g464(.A(new_n887), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  AND4_X1   g466(.A1(new_n853), .A2(new_n872), .A3(new_n852), .A4(new_n875), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n879), .A2(new_n880), .A3(new_n875), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n861), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(new_n895), .B2(new_n886), .ZN(new_n896));
  INV_X1    g471(.A(new_n860), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT41), .B1(new_n852), .B2(new_n853), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n879), .A2(new_n880), .A3(new_n875), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n892), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n889), .B(new_n890), .C1(new_n896), .C2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n888), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n890), .B1(new_n896), .B2(new_n902), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n906), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n895), .A2(new_n891), .A3(new_n886), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT104), .B1(new_n901), .B2(new_n846), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n887), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n911), .B2(new_n889), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n884), .A2(KEYINPUT43), .A3(new_n887), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n907), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n905), .B1(new_n914), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g490(.A(G40), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n481), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n475), .A2(new_n477), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT106), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1384), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n825), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR3_X1    g501(.A1(new_n922), .A2(new_n926), .A3(G1996), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n927), .A2(KEYINPUT46), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(KEYINPUT46), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n922), .A2(new_n926), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n754), .B(new_n756), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n931), .A2(new_n717), .ZN(new_n932));
  AOI22_X1  g507(.A1(new_n928), .A2(new_n929), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  INV_X1    g509(.A(new_n930), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n927), .A2(new_n717), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT107), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n931), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT108), .Z(new_n939));
  NAND3_X1  g514(.A1(new_n930), .A2(G1996), .A3(new_n717), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n702), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n941), .A2(new_n700), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n754), .A2(new_n756), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n935), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n699), .B(new_n942), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n930), .B2(new_n946), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n935), .A2(G1986), .A3(G290), .ZN(new_n948));
  XOR2_X1   g523(.A(new_n948), .B(KEYINPUT48), .Z(new_n949));
  AOI211_X1 g524(.A(new_n934), .B(new_n945), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n500), .A2(new_n823), .A3(new_n503), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n823), .B1(new_n500), .B2(new_n503), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n497), .B(new_n820), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n500), .A2(new_n503), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n956), .B2(new_n819), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT109), .B1(new_n957), .B2(KEYINPUT45), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n959), .B(new_n925), .C1(G164), .C2(G1384), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n955), .A2(KEYINPUT45), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(KEYINPUT110), .A3(new_n920), .A4(new_n921), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n960), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n825), .A2(KEYINPUT45), .A3(new_n923), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n963), .A2(new_n920), .A3(new_n921), .A4(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n967), .A3(new_n679), .ZN(new_n968));
  INV_X1    g543(.A(new_n957), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n971), .B1(new_n924), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(new_n922), .ZN(new_n973));
  INV_X1    g548(.A(G2090), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(G303), .A2(G8), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(G8), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1976), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT52), .B1(G288), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(G288), .A2(new_n982), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n920), .A2(new_n921), .A3(new_n955), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT112), .B(G8), .Z(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n985), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n993), .B1(new_n573), .B2(new_n577), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n572), .A2(new_n576), .A3(G1981), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT49), .ZN(new_n996));
  OAI22_X1  g571(.A1(new_n994), .A2(new_n995), .B1(KEYINPUT116), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(KEYINPUT49), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT116), .B(new_n996), .C1(new_n994), .C2(new_n995), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n999), .A2(new_n991), .A3(new_n989), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT52), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT114), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1006), .A3(KEYINPUT52), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1002), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n922), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n924), .B2(KEYINPUT50), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n974), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n990), .B1(new_n968), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n981), .B(new_n1008), .C1(new_n1013), .C2(new_n980), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT56), .B(G2072), .Z(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1009), .A2(KEYINPUT122), .A3(new_n961), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n965), .B2(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n561), .B(KEYINPUT57), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT121), .B(G1956), .Z(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1020), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1009), .A2(new_n756), .A3(new_n955), .ZN(new_n1026));
  INV_X1    g601(.A(G1348), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n972), .B2(new_n922), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT123), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1029), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n851), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1021), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1025), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT60), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1032), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT60), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n1030), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1039), .A3(new_n592), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT61), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1025), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1041), .B1(new_n1042), .B2(new_n1034), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1034), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT61), .A3(new_n1025), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT58), .B(G1341), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n989), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(G1996), .B2(new_n965), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n550), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT124), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT124), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1052), .A3(new_n550), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g631(.A(KEYINPUT60), .B(new_n851), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1051), .A2(KEYINPUT59), .A3(new_n1053), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1035), .B1(new_n1046), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n926), .B1(new_n925), .B2(new_n969), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n1063));
  OR3_X1    g638(.A1(new_n1062), .A2(new_n922), .A3(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n973), .A2(G1961), .ZN(new_n1065));
  AOI21_X1  g640(.A(G2078), .B1(new_n962), .B2(new_n967), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1064), .B(new_n1065), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(G171), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT126), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT126), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1071), .A3(G171), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n918), .A2(new_n1063), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n926), .A2(new_n1074), .A3(new_n964), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1065), .B(new_n1075), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(G171), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1061), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT118), .B(G2084), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n973), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n725), .B1(new_n1062), .B2(new_n922), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n991), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G168), .A2(new_n990), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1083), .A2(G168), .ZN(new_n1087));
  INV_X1    g662(.A(G8), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1088), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT51), .B1(new_n1089), .B2(new_n1084), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1086), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(G301), .B1(new_n1076), .B2(KEYINPUT127), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(KEYINPUT127), .B2(new_n1076), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1068), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1061), .B1(new_n1094), .B2(G301), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1091), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1060), .A2(new_n1078), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(new_n1073), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1014), .B1(new_n1097), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1083), .A2(G286), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1103), .B1(new_n1014), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT63), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1088), .B(new_n979), .C1(new_n968), .C2(new_n975), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1003), .A2(new_n1006), .A3(KEYINPUT52), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1006), .B1(new_n1003), .B2(KEYINPUT52), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1001), .B(new_n992), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1013), .A2(new_n980), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(KEYINPUT119), .A3(new_n1113), .A4(new_n1104), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1106), .A2(new_n1107), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n976), .A2(G8), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n979), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1112), .A2(KEYINPUT63), .A3(new_n1104), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1001), .A2(new_n982), .A3(new_n683), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n995), .B(KEYINPUT117), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n991), .B(new_n989), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n981), .B2(new_n1111), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT120), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n1126));
  AOI211_X1 g701(.A(new_n1126), .B(new_n1123), .C1(new_n1115), .C2(new_n1118), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1102), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n584), .B(G1986), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n947), .B1(new_n935), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n950), .B1(new_n1128), .B2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g706(.A1(new_n888), .A2(new_n903), .ZN(new_n1133));
  OR3_X1    g707(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1134));
  NOR3_X1   g708(.A1(new_n841), .A2(G229), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1135), .ZN(G225));
  INV_X1    g710(.A(G225), .ZN(G308));
endmodule


