

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755;

  BUF_X1 U373 ( .A(n574), .Z(n351) );
  XNOR2_X1 U374 ( .A(n557), .B(n388), .ZN(n574) );
  XNOR2_X1 U375 ( .A(n358), .B(n464), .ZN(n739) );
  XNOR2_X1 U376 ( .A(G128), .B(G137), .ZN(n481) );
  INV_X1 U377 ( .A(KEYINPUT99), .ZN(n429) );
  XNOR2_X1 U378 ( .A(G119), .B(KEYINPUT3), .ZN(n352) );
  XOR2_X1 U379 ( .A(KEYINPUT16), .B(G122), .Z(n364) );
  XNOR2_X1 U380 ( .A(KEYINPUT69), .B(G110), .ZN(n359) );
  XNOR2_X1 U381 ( .A(KEYINPUT69), .B(G110), .ZN(n356) );
  OR2_X2 U382 ( .A1(n414), .A2(n413), .ZN(n695) );
  XNOR2_X2 U383 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X2 U384 ( .A(n739), .B(G146), .ZN(n477) );
  INV_X1 U385 ( .A(n381), .ZN(n694) );
  NAND2_X1 U386 ( .A1(n381), .A2(n515), .ZN(n380) );
  AND2_X2 U387 ( .A1(n396), .A2(n395), .ZN(n381) );
  XNOR2_X2 U388 ( .A(n569), .B(n417), .ZN(n586) );
  XNOR2_X2 U389 ( .A(n416), .B(KEYINPUT84), .ZN(n569) );
  NOR2_X2 U390 ( .A1(G953), .A2(G237), .ZN(n471) );
  XNOR2_X1 U391 ( .A(G143), .B(G104), .ZN(n447) );
  XOR2_X1 U392 ( .A(G137), .B(G134), .Z(n463) );
  XOR2_X1 U393 ( .A(KEYINPUT11), .B(G122), .Z(n449) );
  NAND2_X1 U394 ( .A1(G234), .A2(G237), .ZN(n418) );
  XNOR2_X1 U395 ( .A(KEYINPUT10), .B(G140), .ZN(n391) );
  INV_X1 U396 ( .A(G214), .ZN(n413) );
  AND2_X2 U397 ( .A1(n366), .A2(n404), .ZN(n383) );
  NAND2_X2 U398 ( .A1(n503), .A2(n461), .ZN(n462) );
  XNOR2_X2 U399 ( .A(n426), .B(KEYINPUT0), .ZN(n503) );
  INV_X1 U400 ( .A(G143), .ZN(n623) );
  NOR2_X1 U401 ( .A1(n688), .A2(n511), .ZN(n513) );
  INV_X1 U402 ( .A(n515), .ZN(n511) );
  AND2_X1 U403 ( .A1(n605), .A2(n604), .ZN(n741) );
  BUF_X1 U404 ( .A(n393), .Z(n374) );
  NAND2_X1 U405 ( .A1(n365), .A2(n403), .ZN(n382) );
  NOR2_X1 U406 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U407 ( .A1(n574), .A2(n386), .ZN(n510) );
  XOR2_X1 U408 ( .A(n555), .B(KEYINPUT6), .Z(n361) );
  XNOR2_X1 U409 ( .A(n495), .B(n494), .ZN(n679) );
  XNOR2_X1 U410 ( .A(n384), .B(n469), .ZN(n722) );
  XNOR2_X1 U411 ( .A(n609), .B(KEYINPUT66), .ZN(n610) );
  XNOR2_X2 U412 ( .A(G119), .B(G110), .ZN(n480) );
  XNOR2_X1 U413 ( .A(G116), .B(G107), .ZN(n430) );
  XNOR2_X2 U414 ( .A(n353), .B(n352), .ZN(n475) );
  XNOR2_X2 U415 ( .A(n376), .B(n357), .ZN(n353) );
  XNOR2_X1 U416 ( .A(n475), .B(n354), .ZN(n733) );
  XNOR2_X1 U417 ( .A(n355), .B(n364), .ZN(n354) );
  XNOR2_X1 U418 ( .A(n375), .B(n356), .ZN(n355) );
  XNOR2_X2 U419 ( .A(G107), .B(G104), .ZN(n375) );
  XNOR2_X2 U420 ( .A(G101), .B(KEYINPUT85), .ZN(n357) );
  XNOR2_X1 U421 ( .A(n358), .B(n369), .ZN(n368) );
  XNOR2_X2 U422 ( .A(n435), .B(KEYINPUT4), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n375), .B(n359), .ZN(n360) );
  INV_X2 U424 ( .A(KEYINPUT18), .ZN(n367) );
  INV_X1 U425 ( .A(KEYINPUT33), .ZN(n401) );
  NAND2_X1 U426 ( .A1(n361), .A2(n401), .ZN(n399) );
  XNOR2_X1 U427 ( .A(G113), .B(G131), .ZN(n444) );
  AND2_X1 U428 ( .A1(n595), .A2(n387), .ZN(n596) );
  INV_X1 U429 ( .A(KEYINPUT44), .ZN(n392) );
  INV_X1 U430 ( .A(n684), .ZN(n386) );
  XNOR2_X1 U431 ( .A(n367), .B(KEYINPUT17), .ZN(n409) );
  XNOR2_X1 U432 ( .A(n446), .B(n411), .ZN(n370) );
  AND2_X1 U433 ( .A1(n400), .A2(n399), .ZN(n396) );
  NOR2_X1 U434 ( .A1(n361), .A2(n401), .ZN(n397) );
  INV_X1 U435 ( .A(G472), .ZN(n615) );
  XNOR2_X1 U436 ( .A(n477), .B(n476), .ZN(n616) );
  XOR2_X1 U437 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n473) );
  XOR2_X2 U438 ( .A(KEYINPUT67), .B(KEYINPUT23), .Z(n482) );
  XNOR2_X1 U439 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U440 ( .A(n451), .B(n740), .ZN(n390) );
  XNOR2_X1 U441 ( .A(n506), .B(n394), .ZN(n393) );
  INV_X1 U442 ( .A(KEYINPUT35), .ZN(n394) );
  INV_X1 U443 ( .A(KEYINPUT22), .ZN(n389) );
  INV_X1 U444 ( .A(KEYINPUT1), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n616), .B(KEYINPUT62), .ZN(n617) );
  XNOR2_X1 U446 ( .A(n552), .B(n551), .ZN(n754) );
  INV_X1 U447 ( .A(n679), .ZN(n385) );
  NOR2_X1 U448 ( .A1(n414), .A2(n627), .ZN(n362) );
  NOR2_X1 U449 ( .A1(n351), .A2(n682), .ZN(n363) );
  NAND2_X1 U450 ( .A1(n383), .A2(n382), .ZN(n530) );
  INV_X1 U451 ( .A(n652), .ZN(n365) );
  NAND2_X1 U452 ( .A1(n652), .A2(KEYINPUT82), .ZN(n366) );
  XNOR2_X2 U453 ( .A(n497), .B(KEYINPUT105), .ZN(n652) );
  XNOR2_X1 U454 ( .A(n733), .B(n368), .ZN(n628) );
  XNOR2_X1 U455 ( .A(n370), .B(n371), .ZN(n369) );
  XNOR2_X1 U456 ( .A(n409), .B(n408), .ZN(n371) );
  XNOR2_X2 U457 ( .A(n407), .B(n623), .ZN(n435) );
  BUF_X1 U458 ( .A(n435), .Z(n372) );
  NAND2_X1 U459 ( .A1(n383), .A2(n382), .ZN(n373) );
  XNOR2_X2 U460 ( .A(G116), .B(G113), .ZN(n376) );
  NAND2_X1 U461 ( .A1(n379), .A2(n377), .ZN(n505) );
  NAND2_X1 U462 ( .A1(n381), .A2(n378), .ZN(n377) );
  NOR2_X1 U463 ( .A1(n511), .A2(n504), .ZN(n378) );
  NAND2_X1 U464 ( .A1(n380), .A2(n504), .ZN(n379) );
  INV_X1 U465 ( .A(n477), .ZN(n384) );
  AND2_X1 U466 ( .A1(n351), .A2(n385), .ZN(n498) );
  OR2_X1 U467 ( .A1(n351), .A2(n385), .ZN(n507) );
  OR2_X1 U468 ( .A1(n351), .A2(n386), .ZN(n685) );
  INV_X1 U469 ( .A(n351), .ZN(n387) );
  XNOR2_X2 U470 ( .A(n440), .B(G478), .ZN(n517) );
  INV_X2 U471 ( .A(n410), .ZN(n446) );
  NAND2_X1 U472 ( .A1(n415), .A2(n695), .ZN(n416) );
  NAND2_X1 U473 ( .A1(n478), .A2(n361), .ZN(n508) );
  XNOR2_X2 U474 ( .A(n462), .B(n389), .ZN(n478) );
  XNOR2_X1 U475 ( .A(n452), .B(n390), .ZN(n645) );
  XNOR2_X1 U476 ( .A(n446), .B(n391), .ZN(n740) );
  NAND2_X1 U477 ( .A1(n374), .A2(n392), .ZN(n529) );
  NOR2_X1 U478 ( .A1(n393), .A2(n392), .ZN(n509) );
  XNOR2_X1 U479 ( .A(n374), .B(G122), .ZN(G24) );
  NAND2_X1 U480 ( .A1(n397), .A2(n398), .ZN(n395) );
  INV_X1 U481 ( .A(n510), .ZN(n398) );
  NAND2_X1 U482 ( .A1(n510), .A2(n401), .ZN(n400) );
  XNOR2_X2 U483 ( .A(n402), .B(n615), .ZN(n555) );
  NAND2_X1 U484 ( .A1(n616), .A2(n490), .ZN(n402) );
  NOR2_X1 U485 ( .A1(n626), .A2(KEYINPUT82), .ZN(n403) );
  NAND2_X1 U486 ( .A1(n626), .A2(KEYINPUT82), .ZN(n404) );
  NAND2_X1 U487 ( .A1(n530), .A2(KEYINPUT44), .ZN(n502) );
  INV_X1 U488 ( .A(n415), .ZN(n547) );
  XNOR2_X2 U489 ( .A(n405), .B(n362), .ZN(n415) );
  NAND2_X1 U490 ( .A1(n628), .A2(n534), .ZN(n405) );
  NOR2_X2 U491 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X2 U492 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X2 U493 ( .A1(n614), .A2(n676), .ZN(n643) );
  XOR2_X1 U494 ( .A(KEYINPUT78), .B(n585), .Z(n406) );
  XNOR2_X1 U495 ( .A(n463), .B(G131), .ZN(n464) );
  XNOR2_X1 U496 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U497 ( .A(n432), .B(n431), .ZN(n433) );
  INV_X1 U498 ( .A(KEYINPUT110), .ZN(n536) );
  INV_X1 U499 ( .A(KEYINPUT40), .ZN(n550) );
  XNOR2_X1 U500 ( .A(n550), .B(KEYINPUT111), .ZN(n551) );
  INV_X1 U501 ( .A(KEYINPUT63), .ZN(n621) );
  XNOR2_X2 U502 ( .A(G128), .B(KEYINPUT75), .ZN(n407) );
  XNOR2_X1 U503 ( .A(KEYINPUT86), .B(KEYINPUT74), .ZN(n408) );
  XNOR2_X2 U504 ( .A(G146), .B(G125), .ZN(n410) );
  INV_X2 U505 ( .A(G953), .ZN(n743) );
  NAND2_X1 U506 ( .A1(n743), .A2(G224), .ZN(n411) );
  XNOR2_X1 U507 ( .A(G902), .B(KEYINPUT15), .ZN(n534) );
  NOR2_X1 U508 ( .A1(G237), .A2(G902), .ZN(n412) );
  XNOR2_X1 U509 ( .A(n412), .B(KEYINPUT68), .ZN(n414) );
  INV_X1 U510 ( .A(G210), .ZN(n627) );
  XNOR2_X1 U511 ( .A(KEYINPUT71), .B(KEYINPUT19), .ZN(n417) );
  XNOR2_X1 U512 ( .A(n418), .B(KEYINPUT14), .ZN(n421) );
  NAND2_X1 U513 ( .A1(n421), .A2(G902), .ZN(n419) );
  XNOR2_X1 U514 ( .A(n419), .B(KEYINPUT87), .ZN(n538) );
  NOR2_X1 U515 ( .A1(G898), .A2(n743), .ZN(n735) );
  NAND2_X1 U516 ( .A1(n538), .A2(n735), .ZN(n420) );
  XOR2_X1 U517 ( .A(KEYINPUT88), .B(n420), .Z(n422) );
  NAND2_X1 U518 ( .A1(G952), .A2(n421), .ZN(n709) );
  NOR2_X1 U519 ( .A1(G953), .A2(n709), .ZN(n541) );
  NOR2_X1 U520 ( .A1(n422), .A2(n541), .ZN(n424) );
  INV_X1 U521 ( .A(KEYINPUT89), .ZN(n423) );
  NOR2_X2 U522 ( .A1(n586), .A2(n425), .ZN(n426) );
  XOR2_X1 U523 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n428) );
  XNOR2_X1 U524 ( .A(G134), .B(G122), .ZN(n427) );
  XNOR2_X1 U525 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U526 ( .A(n433), .B(KEYINPUT98), .Z(n439) );
  NAND2_X1 U527 ( .A1(G234), .A2(n743), .ZN(n434) );
  XOR2_X1 U528 ( .A(KEYINPUT8), .B(n434), .Z(n485) );
  AND2_X1 U529 ( .A1(n485), .A2(G217), .ZN(n437) );
  XNOR2_X1 U530 ( .A(n372), .B(KEYINPUT7), .ZN(n436) );
  XNOR2_X1 U531 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n439), .B(n438), .ZN(n640) );
  INV_X1 U533 ( .A(G902), .ZN(n490) );
  NAND2_X1 U534 ( .A1(n640), .A2(n490), .ZN(n440) );
  XOR2_X1 U535 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n442) );
  XNOR2_X1 U536 ( .A(KEYINPUT12), .B(KEYINPUT97), .ZN(n441) );
  XNOR2_X1 U537 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U538 ( .A(n443), .B(KEYINPUT95), .Z(n445) );
  XNOR2_X1 U539 ( .A(n445), .B(n444), .ZN(n452) );
  NAND2_X1 U540 ( .A1(G214), .A2(n471), .ZN(n448) );
  XNOR2_X1 U541 ( .A(n448), .B(n447), .ZN(n450) );
  NAND2_X1 U542 ( .A1(n645), .A2(n490), .ZN(n454) );
  XOR2_X1 U543 ( .A(KEYINPUT13), .B(G475), .Z(n453) );
  XNOR2_X2 U544 ( .A(n454), .B(n453), .ZN(n518) );
  NOR2_X2 U545 ( .A1(n517), .A2(n518), .ZN(n455) );
  XNOR2_X1 U546 ( .A(n455), .B(KEYINPUT103), .ZN(n698) );
  XOR2_X1 U547 ( .A(KEYINPUT21), .B(KEYINPUT90), .Z(n458) );
  NAND2_X1 U548 ( .A1(n534), .A2(G234), .ZN(n456) );
  XNOR2_X1 U549 ( .A(n456), .B(KEYINPUT20), .ZN(n491) );
  NAND2_X1 U550 ( .A1(n491), .A2(G221), .ZN(n457) );
  XNOR2_X1 U551 ( .A(n458), .B(n457), .ZN(n678) );
  INV_X1 U552 ( .A(n678), .ZN(n459) );
  NOR2_X1 U553 ( .A1(n698), .A2(n459), .ZN(n460) );
  XNOR2_X1 U554 ( .A(n460), .B(KEYINPUT104), .ZN(n461) );
  NAND2_X1 U555 ( .A1(G227), .A2(n743), .ZN(n465) );
  XNOR2_X1 U556 ( .A(n465), .B(G140), .ZN(n466) );
  XNOR2_X1 U557 ( .A(n360), .B(n466), .ZN(n467) );
  XOR2_X1 U558 ( .A(n467), .B(KEYINPUT73), .Z(n468) );
  XNOR2_X1 U559 ( .A(n468), .B(G101), .ZN(n469) );
  NOR2_X2 U560 ( .A1(n722), .A2(G902), .ZN(n470) );
  XNOR2_X2 U561 ( .A(n470), .B(G469), .ZN(n557) );
  NAND2_X1 U562 ( .A1(n471), .A2(G210), .ZN(n472) );
  XNOR2_X1 U563 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U564 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U565 ( .A1(n478), .A2(n363), .ZN(n479) );
  XNOR2_X1 U566 ( .A(n479), .B(KEYINPUT65), .ZN(n496) );
  XNOR2_X1 U567 ( .A(n480), .B(KEYINPUT24), .ZN(n484) );
  XNOR2_X1 U568 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U569 ( .A(n484), .B(n483), .Z(n489) );
  NAND2_X1 U570 ( .A1(G221), .A2(n485), .ZN(n487) );
  INV_X1 U571 ( .A(n740), .ZN(n486) );
  XNOR2_X1 U572 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U573 ( .A(n489), .B(n488), .ZN(n637) );
  NAND2_X1 U574 ( .A1(n637), .A2(n490), .ZN(n495) );
  NAND2_X1 U575 ( .A1(n491), .A2(G217), .ZN(n493) );
  XOR2_X1 U576 ( .A(KEYINPUT25), .B(KEYINPUT72), .Z(n492) );
  XNOR2_X1 U577 ( .A(n493), .B(n492), .ZN(n494) );
  NAND2_X1 U578 ( .A1(n496), .A2(n385), .ZN(n497) );
  INV_X1 U579 ( .A(n508), .ZN(n499) );
  NAND2_X1 U580 ( .A1(n499), .A2(n498), .ZN(n501) );
  INV_X1 U581 ( .A(KEYINPUT32), .ZN(n500) );
  XNOR2_X2 U582 ( .A(n501), .B(n500), .ZN(n626) );
  XNOR2_X1 U583 ( .A(n502), .B(KEYINPUT64), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n679), .A2(n678), .ZN(n684) );
  BUF_X1 U585 ( .A(n503), .Z(n515) );
  INV_X1 U586 ( .A(KEYINPUT34), .ZN(n504) );
  AND2_X1 U587 ( .A1(n517), .A2(n518), .ZN(n579) );
  NAND2_X1 U588 ( .A1(n505), .A2(n579), .ZN(n506) );
  NOR2_X1 U589 ( .A1(n508), .A2(n507), .ZN(n654) );
  NOR2_X1 U590 ( .A1(n509), .A2(n654), .ZN(n523) );
  OR2_X1 U591 ( .A1(n510), .A2(n555), .ZN(n688) );
  XOR2_X1 U592 ( .A(KEYINPUT93), .B(KEYINPUT31), .Z(n512) );
  XNOR2_X1 U593 ( .A(n513), .B(n512), .ZN(n669) );
  NOR2_X1 U594 ( .A1(n557), .A2(n684), .ZN(n514) );
  XNOR2_X1 U595 ( .A(KEYINPUT91), .B(n514), .ZN(n537) );
  INV_X1 U596 ( .A(n555), .ZN(n682) );
  NOR2_X1 U597 ( .A1(n537), .A2(n682), .ZN(n516) );
  NAND2_X1 U598 ( .A1(n516), .A2(n515), .ZN(n656) );
  NAND2_X1 U599 ( .A1(n669), .A2(n656), .ZN(n520) );
  INV_X1 U600 ( .A(n517), .ZN(n519) );
  NOR2_X1 U601 ( .A1(n519), .A2(n518), .ZN(n660) );
  XNOR2_X1 U602 ( .A(KEYINPUT101), .B(n660), .ZN(n601) );
  NAND2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n565) );
  NAND2_X1 U604 ( .A1(n601), .A2(n565), .ZN(n582) );
  NAND2_X1 U605 ( .A1(n520), .A2(n582), .ZN(n521) );
  XNOR2_X1 U606 ( .A(n521), .B(KEYINPUT102), .ZN(n522) );
  NAND2_X1 U607 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U608 ( .A(n524), .B(KEYINPUT81), .ZN(n525) );
  NAND2_X1 U609 ( .A1(n526), .A2(n525), .ZN(n528) );
  INV_X1 U610 ( .A(KEYINPUT80), .ZN(n527) );
  XNOR2_X1 U611 ( .A(n528), .B(n527), .ZN(n532) );
  OR2_X1 U612 ( .A1(n373), .A2(n529), .ZN(n531) );
  NAND2_X1 U613 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X2 U614 ( .A(n533), .B(KEYINPUT45), .ZN(n727) );
  INV_X1 U615 ( .A(n534), .ZN(n608) );
  NAND2_X1 U616 ( .A1(n727), .A2(n608), .ZN(n535) );
  XNOR2_X1 U617 ( .A(n535), .B(KEYINPUT79), .ZN(n607) );
  XNOR2_X1 U618 ( .A(n537), .B(n536), .ZN(n546) );
  NAND2_X1 U619 ( .A1(n538), .A2(G953), .ZN(n539) );
  NOR2_X1 U620 ( .A1(G900), .A2(n539), .ZN(n540) );
  NOR2_X1 U621 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U622 ( .A(KEYINPUT76), .B(n542), .ZN(n553) );
  NAND2_X1 U623 ( .A1(n682), .A2(n695), .ZN(n543) );
  XNOR2_X1 U624 ( .A(KEYINPUT30), .B(n543), .ZN(n544) );
  NOR2_X1 U625 ( .A1(n553), .A2(n544), .ZN(n545) );
  NAND2_X1 U626 ( .A1(n546), .A2(n545), .ZN(n581) );
  INV_X1 U627 ( .A(KEYINPUT38), .ZN(n548) );
  XNOR2_X1 U628 ( .A(n547), .B(n548), .ZN(n560) );
  NOR2_X1 U629 ( .A1(n581), .A2(n560), .ZN(n549) );
  XNOR2_X1 U630 ( .A(n549), .B(KEYINPUT39), .ZN(n602) );
  NOR2_X1 U631 ( .A1(n602), .A2(n565), .ZN(n552) );
  XOR2_X1 U632 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n563) );
  NOR2_X1 U633 ( .A1(n679), .A2(n553), .ZN(n554) );
  NAND2_X1 U634 ( .A1(n678), .A2(n554), .ZN(n566) );
  NOR2_X1 U635 ( .A1(n555), .A2(n566), .ZN(n556) );
  XNOR2_X1 U636 ( .A(KEYINPUT28), .B(n556), .ZN(n559) );
  INV_X1 U637 ( .A(n557), .ZN(n558) );
  NAND2_X1 U638 ( .A1(n559), .A2(n558), .ZN(n588) );
  INV_X1 U639 ( .A(n560), .ZN(n696) );
  NAND2_X1 U640 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U641 ( .A1(n698), .A2(n699), .ZN(n561) );
  XOR2_X1 U642 ( .A(KEYINPUT41), .B(n561), .Z(n692) );
  INV_X1 U643 ( .A(n692), .ZN(n712) );
  OR2_X1 U644 ( .A1(n588), .A2(n712), .ZN(n562) );
  XNOR2_X1 U645 ( .A(n563), .B(n562), .ZN(n750) );
  NOR2_X1 U646 ( .A1(n754), .A2(n750), .ZN(n564) );
  XOR2_X1 U647 ( .A(KEYINPUT46), .B(n564), .Z(n577) );
  XOR2_X1 U648 ( .A(KEYINPUT106), .B(n565), .Z(n663) );
  INV_X1 U649 ( .A(n663), .ZN(n666) );
  NOR2_X1 U650 ( .A1(n361), .A2(n566), .ZN(n567) );
  XNOR2_X1 U651 ( .A(n567), .B(KEYINPUT107), .ZN(n568) );
  NOR2_X1 U652 ( .A1(n666), .A2(n568), .ZN(n595) );
  BUF_X1 U653 ( .A(n569), .Z(n570) );
  INV_X1 U654 ( .A(n570), .ZN(n571) );
  NAND2_X1 U655 ( .A1(n595), .A2(n571), .ZN(n573) );
  XNOR2_X1 U656 ( .A(KEYINPUT36), .B(KEYINPUT83), .ZN(n572) );
  XNOR2_X1 U657 ( .A(n573), .B(n572), .ZN(n575) );
  NAND2_X1 U658 ( .A1(n575), .A2(n351), .ZN(n576) );
  XNOR2_X1 U659 ( .A(KEYINPUT113), .B(n576), .ZN(n751) );
  NOR2_X1 U660 ( .A1(n577), .A2(n751), .ZN(n593) );
  INV_X1 U661 ( .A(n547), .ZN(n578) );
  NAND2_X1 U662 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U663 ( .A1(n581), .A2(n580), .ZN(n624) );
  INV_X1 U664 ( .A(n624), .ZN(n584) );
  INV_X1 U665 ( .A(n582), .ZN(n700) );
  NAND2_X1 U666 ( .A1(n700), .A2(KEYINPUT47), .ZN(n583) );
  NAND2_X1 U667 ( .A1(n584), .A2(n583), .ZN(n585) );
  BUF_X1 U668 ( .A(n586), .Z(n587) );
  NOR2_X1 U669 ( .A1(n588), .A2(n587), .ZN(n664) );
  XOR2_X1 U670 ( .A(KEYINPUT47), .B(n664), .Z(n590) );
  NAND2_X1 U671 ( .A1(n664), .A2(n700), .ZN(n589) );
  NAND2_X1 U672 ( .A1(n590), .A2(n589), .ZN(n591) );
  AND2_X1 U673 ( .A1(n406), .A2(n591), .ZN(n592) );
  AND2_X1 U674 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U675 ( .A(n594), .B(KEYINPUT48), .ZN(n605) );
  XOR2_X1 U676 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n598) );
  NAND2_X1 U677 ( .A1(n596), .A2(n695), .ZN(n597) );
  XNOR2_X1 U678 ( .A(n598), .B(n597), .ZN(n599) );
  XNOR2_X1 U679 ( .A(n599), .B(KEYINPUT43), .ZN(n600) );
  AND2_X1 U680 ( .A1(n600), .A2(n547), .ZN(n625) );
  NOR2_X1 U681 ( .A1(n625), .A2(n603), .ZN(n604) );
  XNOR2_X1 U682 ( .A(n741), .B(KEYINPUT70), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n608), .A2(KEYINPUT2), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n614) );
  INV_X1 U686 ( .A(n741), .ZN(n613) );
  INV_X1 U687 ( .A(n727), .ZN(n612) );
  NOR2_X2 U688 ( .A1(n613), .A2(n612), .ZN(n674) );
  NAND2_X1 U689 ( .A1(n674), .A2(KEYINPUT2), .ZN(n676) );
  NOR2_X1 U690 ( .A1(n643), .A2(n615), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(n617), .ZN(n620) );
  INV_X1 U692 ( .A(G952), .ZN(n619) );
  AND2_X1 U693 ( .A1(n619), .A2(G953), .ZN(n726) );
  NOR2_X1 U694 ( .A1(n620), .A2(n726), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(G57) );
  XNOR2_X1 U696 ( .A(n624), .B(n623), .ZN(G45) );
  XOR2_X1 U697 ( .A(n625), .B(G140), .Z(G42) );
  XOR2_X1 U698 ( .A(n626), .B(G119), .Z(G21) );
  NOR2_X1 U699 ( .A1(n643), .A2(n627), .ZN(n632) );
  BUF_X1 U700 ( .A(n628), .Z(n629) );
  XOR2_X1 U701 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n630) );
  XNOR2_X1 U702 ( .A(n629), .B(n630), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n633), .A2(n726), .ZN(n635) );
  XNOR2_X1 U705 ( .A(KEYINPUT122), .B(KEYINPUT56), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G51) );
  INV_X1 U707 ( .A(n643), .ZN(n718) );
  NAND2_X1 U708 ( .A1(n718), .A2(G217), .ZN(n636) );
  XOR2_X1 U709 ( .A(n637), .B(n636), .Z(n638) );
  NOR2_X1 U710 ( .A1(n638), .A2(n726), .ZN(G66) );
  NAND2_X1 U711 ( .A1(n718), .A2(G478), .ZN(n639) );
  XOR2_X1 U712 ( .A(n640), .B(n639), .Z(n641) );
  NOR2_X1 U713 ( .A1(n641), .A2(n726), .ZN(G63) );
  INV_X1 U714 ( .A(G475), .ZN(n642) );
  XNOR2_X1 U715 ( .A(KEYINPUT125), .B(KEYINPUT59), .ZN(n644) );
  XOR2_X1 U716 ( .A(n645), .B(n644), .Z(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(n649) );
  INV_X1 U718 ( .A(n726), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n651) );
  INV_X1 U720 ( .A(KEYINPUT60), .ZN(n650) );
  XNOR2_X1 U721 ( .A(n651), .B(n650), .ZN(G60) );
  BUF_X1 U722 ( .A(n652), .Z(n653) );
  XOR2_X1 U723 ( .A(n653), .B(G110), .Z(G12) );
  XOR2_X1 U724 ( .A(G101), .B(n654), .Z(G3) );
  NOR2_X1 U725 ( .A1(n666), .A2(n656), .ZN(n655) );
  XOR2_X1 U726 ( .A(G104), .B(n655), .Z(G6) );
  INV_X1 U727 ( .A(n660), .ZN(n670) );
  NOR2_X1 U728 ( .A1(n670), .A2(n656), .ZN(n658) );
  XNOR2_X1 U729 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n657) );
  XNOR2_X1 U730 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(G107), .B(n659), .ZN(G9) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  NAND2_X1 U733 ( .A1(n664), .A2(n660), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(G30) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U736 ( .A(n665), .B(G146), .ZN(G48) );
  NOR2_X1 U737 ( .A1(n666), .A2(n669), .ZN(n667) );
  XOR2_X1 U738 ( .A(KEYINPUT114), .B(n667), .Z(n668) );
  XNOR2_X1 U739 ( .A(G113), .B(n668), .ZN(G15) );
  NOR2_X1 U740 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U741 ( .A(G116), .B(KEYINPUT115), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n672), .B(n671), .ZN(G18) );
  XNOR2_X1 U743 ( .A(G134), .B(n603), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n673), .B(KEYINPUT117), .ZN(G36) );
  NOR2_X1 U745 ( .A1(n674), .A2(KEYINPUT2), .ZN(n675) );
  XNOR2_X1 U746 ( .A(n675), .B(KEYINPUT77), .ZN(n677) );
  AND2_X1 U747 ( .A1(n677), .A2(n676), .ZN(n711) );
  NOR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U749 ( .A(KEYINPUT49), .B(n680), .Z(n681) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n683), .B(KEYINPUT118), .ZN(n687) );
  XNOR2_X1 U752 ( .A(KEYINPUT50), .B(n685), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U755 ( .A(KEYINPUT51), .B(n690), .Z(n691) );
  NAND2_X1 U756 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U757 ( .A(n693), .B(KEYINPUT119), .ZN(n706) );
  NOR2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U759 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U760 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U761 ( .A(n701), .B(KEYINPUT120), .ZN(n702) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U763 ( .A1(n694), .A2(n704), .ZN(n705) );
  NOR2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U765 ( .A(n707), .B(KEYINPUT52), .ZN(n708) );
  NOR2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U767 ( .A1(n694), .A2(n712), .ZN(n713) );
  XNOR2_X1 U768 ( .A(n713), .B(KEYINPUT121), .ZN(n714) );
  NAND2_X1 U769 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X2 U770 ( .A1(n716), .A2(G953), .ZN(n717) );
  XNOR2_X1 U771 ( .A(n717), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U772 ( .A1(n718), .A2(G469), .ZN(n724) );
  XOR2_X1 U773 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n720) );
  XNOR2_X1 U774 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n719) );
  XNOR2_X1 U775 ( .A(n720), .B(n719), .ZN(n721) );
  XOR2_X1 U776 ( .A(n722), .B(n721), .Z(n723) );
  XNOR2_X1 U777 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U778 ( .A1(n726), .A2(n725), .ZN(G54) );
  BUF_X1 U779 ( .A(n727), .Z(n728) );
  NAND2_X1 U780 ( .A1(n728), .A2(n743), .ZN(n732) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n729) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n729), .ZN(n730) );
  NAND2_X1 U783 ( .A1(n730), .A2(G898), .ZN(n731) );
  NAND2_X1 U784 ( .A1(n732), .A2(n731), .ZN(n738) );
  BUF_X1 U785 ( .A(n733), .Z(n734) );
  XOR2_X1 U786 ( .A(KEYINPUT126), .B(n734), .Z(n736) );
  NOR2_X1 U787 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U788 ( .A(n738), .B(n737), .ZN(G69) );
  XOR2_X1 U789 ( .A(n740), .B(n739), .Z(n745) );
  INV_X1 U790 ( .A(n745), .ZN(n742) );
  XNOR2_X1 U791 ( .A(n742), .B(n741), .ZN(n744) );
  NAND2_X1 U792 ( .A1(n744), .A2(n743), .ZN(n749) );
  XNOR2_X1 U793 ( .A(G227), .B(n745), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G953), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U797 ( .A(G137), .B(n750), .Z(G39) );
  XNOR2_X1 U798 ( .A(n751), .B(KEYINPUT116), .ZN(n752) );
  XNOR2_X1 U799 ( .A(n752), .B(KEYINPUT37), .ZN(n753) );
  XNOR2_X1 U800 ( .A(G125), .B(n753), .ZN(G27) );
  XNOR2_X1 U801 ( .A(G131), .B(KEYINPUT127), .ZN(n755) );
  XNOR2_X1 U802 ( .A(n755), .B(n754), .ZN(G33) );
endmodule

