//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT73), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT68), .B(G237), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT69), .A2(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT69), .A2(G953), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G210), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n191), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(new_n193), .A2(new_n194), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n198), .A2(G210), .A3(new_n192), .A4(new_n190), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n197), .A2(new_n201), .A3(new_n199), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G116), .ZN(new_n207));
  INV_X1    g021(.A(G116), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(KEYINPUT2), .B(G113), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n215), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n212), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  INV_X1    g035(.A(G134), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G137), .ZN(new_n223));
  AOI21_X1  g037(.A(G131), .B1(new_n222), .B2(G137), .ZN(new_n224));
  INV_X1    g038(.A(G137), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT11), .A3(G134), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n224), .A3(new_n229), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n222), .A2(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n223), .A2(new_n226), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G143), .ZN(new_n237));
  INV_X1    g051(.A(G143), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G128), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n225), .A2(G134), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(new_n248), .B2(new_n232), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n228), .B2(new_n230), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n251), .B(KEYINPUT1), .C1(new_n238), .C2(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G128), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n251), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n240), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT1), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n237), .A2(new_n239), .A3(new_n256), .A4(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n235), .A2(new_n246), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n205), .B1(new_n220), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n250), .A2(new_n258), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n261), .A2(KEYINPUT66), .B1(new_n235), .B2(new_n246), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n258), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT30), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n228), .A2(new_n230), .B1(G131), .B2(new_n233), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n261), .B1(new_n266), .B2(new_n245), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n219), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n260), .B1(new_n265), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n220), .B1(new_n259), .B2(KEYINPUT30), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n250), .A2(new_n258), .A3(new_n263), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n263), .B1(new_n250), .B2(new_n258), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n266), .A2(new_n245), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n273), .B1(new_n277), .B2(KEYINPUT30), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .A3(new_n260), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n272), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n261), .A2(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n235), .A2(new_n246), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n264), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n219), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n259), .A2(new_n220), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n219), .B1(new_n267), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT28), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n205), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n280), .A2(new_n281), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n281), .B1(new_n280), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n189), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(KEYINPUT32), .B(new_n189), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT75), .B(G902), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n278), .A2(new_n287), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n197), .A2(new_n201), .A3(new_n199), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n201), .B1(new_n197), .B2(new_n199), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n301), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n288), .A2(new_n292), .A3(new_n205), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n291), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n220), .B1(new_n259), .B2(KEYINPUT71), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n282), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT74), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n292), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n267), .A2(new_n219), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n287), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT28), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n318), .A2(new_n301), .A3(new_n205), .ZN(new_n319));
  OAI21_X1  g133(.A(G472), .B1(new_n308), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n298), .A2(new_n299), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G217), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n300), .B2(G234), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(KEYINPUT77), .A2(G125), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT77), .A2(G125), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OR3_X1    g141(.A1(new_n327), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT77), .A2(G125), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n330));
  NAND2_X1  g144(.A1(KEYINPUT77), .A2(G125), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n329), .A2(new_n330), .A3(G140), .A4(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G140), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n325), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT78), .B1(new_n335), .B2(G140), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n337), .A2(KEYINPUT79), .A3(KEYINPUT16), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT79), .B1(new_n337), .B2(KEYINPUT16), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n328), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n236), .ZN(new_n341));
  OAI211_X1 g155(.A(G146), .B(new_n328), .C1(new_n338), .C2(new_n339), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g157(.A(KEYINPUT24), .B(G110), .Z(new_n344));
  XNOR2_X1  g158(.A(G119), .B(G128), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(KEYINPUT76), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n206), .B2(G128), .ZN(new_n349));
  INV_X1    g163(.A(G128), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT23), .A3(G119), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n351), .C1(G119), .C2(new_n350), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(G110), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G125), .B(G140), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n236), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n352), .A2(G110), .B1(new_n345), .B2(new_n344), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n342), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n198), .A2(G221), .A3(G234), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT22), .B(G137), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n355), .A2(new_n359), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n362), .ZN(new_n364));
  INV_X1    g178(.A(new_n354), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n341), .B2(new_n342), .ZN(new_n366));
  INV_X1    g180(.A(new_n359), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n364), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n363), .A2(new_n368), .A3(new_n300), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n363), .A2(new_n368), .A3(KEYINPUT25), .A4(new_n300), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n324), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n363), .A2(new_n368), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n323), .A2(G902), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT80), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G469), .ZN(new_n379));
  INV_X1    g193(.A(new_n258), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G104), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G107), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n383), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(G104), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT3), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n389), .B1(new_n388), .B2(KEYINPUT3), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n381), .B(new_n387), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n385), .A2(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n394), .A3(KEYINPUT83), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n395), .B(G101), .C1(KEYINPUT83), .C2(new_n388), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n380), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT84), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n257), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n256), .B1(G143), .B2(new_n236), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n240), .B1(new_n401), .B2(new_n350), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n257), .A2(new_n399), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n393), .B(new_n396), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT12), .B1(new_n406), .B2(new_n235), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT12), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(new_n266), .C1(new_n398), .C2(new_n405), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n397), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT10), .A3(new_n258), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n387), .B1(new_n391), .B2(new_n392), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G101), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n393), .A2(KEYINPUT4), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT82), .B1(new_n386), .B2(new_n384), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n390), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n381), .B1(new_n418), .B2(new_n387), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n246), .B(new_n415), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT10), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n405), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n412), .A2(new_n420), .A3(new_n422), .A4(new_n266), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n198), .A2(G227), .ZN(new_n424));
  XOR2_X1   g238(.A(G110), .B(G140), .Z(new_n425));
  XOR2_X1   g239(.A(new_n424), .B(new_n425), .Z(new_n426));
  NAND2_X1  g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n410), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n412), .A2(new_n420), .A3(new_n422), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n235), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n430), .B2(new_n423), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n379), .B(new_n300), .C1(new_n428), .C2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n423), .B1(new_n407), .B2(new_n409), .ZN(new_n433));
  INV_X1    g247(.A(new_n426), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n430), .B1(new_n427), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT85), .B1(new_n423), .B2(new_n426), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n435), .B(G469), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(G469), .A2(G902), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n432), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT9), .B(G234), .ZN(new_n442));
  OAI21_X1  g256(.A(G221), .B1(new_n442), .B2(G902), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n443), .B(KEYINPUT81), .Z(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n445), .B(KEYINPUT91), .Z(new_n446));
  OR3_X1    g260(.A1(new_n242), .A2(new_n244), .A3(new_n327), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n255), .A2(new_n327), .A3(new_n257), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G224), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n450), .A2(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n449), .B(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n219), .B(new_n415), .C1(new_n416), .C2(new_n419), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n213), .B1(new_n207), .B2(new_n209), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT5), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G113), .B1(new_n207), .B2(KEYINPUT5), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(new_n218), .A3(new_n393), .A4(new_n396), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT6), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n453), .A2(new_n460), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n463), .B(KEYINPUT87), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(KEYINPUT6), .A3(new_n468), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n452), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G902), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT88), .B(KEYINPUT8), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n463), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT5), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n211), .B2(new_n214), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n218), .B1(new_n478), .B2(new_n457), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n397), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT89), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n457), .B1(KEYINPUT5), .B2(new_n212), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n217), .B2(new_n212), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n480), .A2(new_n481), .B1(new_n411), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n479), .A2(KEYINPUT89), .A3(new_n397), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n476), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n451), .A2(KEYINPUT7), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n449), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n448), .A2(KEYINPUT90), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n447), .A2(KEYINPUT90), .A3(new_n448), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n464), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n473), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n446), .B1(new_n472), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n464), .A2(new_n488), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n480), .A2(new_n481), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n411), .A2(new_n483), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n485), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n475), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n452), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n464), .A2(KEYINPUT6), .B1(new_n466), .B2(new_n468), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n503));
  AOI211_X1 g317(.A(new_n503), .B(new_n467), .C1(new_n453), .C2(new_n460), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n500), .A2(new_n505), .A3(new_n445), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n494), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G214), .B1(G237), .B2(G902), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n441), .A2(new_n444), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G478), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(KEYINPUT15), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n442), .A2(new_n322), .A3(G953), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n238), .A2(G128), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n350), .A2(G143), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n222), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n222), .B1(new_n514), .B2(new_n515), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n208), .A2(G122), .ZN(new_n519));
  INV_X1    g333(.A(G122), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G116), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(G107), .B1(new_n519), .B2(new_n522), .ZN(new_n524));
  OAI22_X1  g338(.A1(new_n517), .A2(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n521), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT94), .ZN(new_n529));
  AOI21_X1  g343(.A(G107), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n525), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n514), .A2(new_n515), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(G134), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n520), .A2(G116), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n382), .B1(new_n535), .B2(KEYINPUT14), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n534), .A2(new_n516), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n529), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT94), .B1(new_n519), .B2(new_n521), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n382), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT96), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n350), .B2(G143), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n238), .A2(KEYINPUT13), .A3(G128), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n515), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G134), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT95), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT95), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n550), .A3(G134), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n528), .A2(G107), .A3(new_n529), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n541), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n554), .A3(new_n516), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n513), .B1(new_n543), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n531), .B1(new_n525), .B2(new_n530), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n538), .A2(new_n541), .A3(KEYINPUT96), .ZN(new_n558));
  AND4_X1   g372(.A1(new_n555), .A2(new_n557), .A3(new_n558), .A4(new_n513), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n300), .B1(new_n556), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT97), .ZN(new_n561));
  INV_X1    g375(.A(new_n300), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n539), .A2(new_n540), .A3(new_n382), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n516), .B1(new_n563), .B2(new_n530), .ZN(new_n564));
  INV_X1    g378(.A(new_n551), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n550), .B1(new_n547), .B2(G134), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n557), .B(new_n558), .C1(new_n564), .C2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n513), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n555), .A2(new_n557), .A3(new_n558), .A4(new_n513), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT97), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n512), .B1(new_n561), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n511), .B1(new_n560), .B2(KEYINPUT97), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n575), .A2(KEYINPUT98), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n572), .A2(new_n573), .ZN(new_n579));
  AOI211_X1 g393(.A(KEYINPUT97), .B(new_n562), .C1(new_n570), .C2(new_n571), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n511), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n576), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT92), .B(G143), .ZN(new_n585));
  INV_X1    g399(.A(G214), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n195), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(KEYINPUT92), .A2(G143), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n198), .A2(G214), .A3(new_n192), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G131), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n587), .A2(new_n247), .A3(new_n589), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(KEYINPUT17), .A3(G131), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n341), .A2(new_n342), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(G113), .B(G122), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(new_n385), .ZN(new_n598));
  AND2_X1   g412(.A1(KEYINPUT18), .A2(G131), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n590), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n357), .B1(new_n337), .B2(new_n236), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n590), .A2(KEYINPUT93), .A3(new_n599), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT93), .B1(new_n590), .B2(new_n599), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n600), .B(new_n601), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n596), .A2(new_n598), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n598), .B1(new_n596), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n473), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G475), .ZN(new_n609));
  INV_X1    g423(.A(G952), .ZN(new_n610));
  AOI211_X1 g424(.A(G953), .B(new_n610), .C1(G234), .C2(G237), .ZN(new_n611));
  INV_X1    g425(.A(new_n198), .ZN(new_n612));
  NAND2_X1  g426(.A1(G234), .A2(G237), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n562), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT99), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT21), .B(G898), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT20), .ZN(new_n619));
  INV_X1    g433(.A(new_n598), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n591), .A2(new_n593), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT19), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n356), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n337), .B2(new_n622), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n624), .A2(G146), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n621), .A2(new_n342), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n601), .B1(new_n590), .B2(new_n599), .ZN(new_n627));
  INV_X1    g441(.A(new_n604), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n602), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n620), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n596), .A2(new_n598), .A3(new_n605), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(G475), .A2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n619), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n633), .ZN(new_n635));
  AOI211_X1 g449(.A(KEYINPUT20), .B(new_n635), .C1(new_n630), .C2(new_n631), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n609), .B(new_n618), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n509), .A2(new_n584), .A3(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n321), .A2(new_n378), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT100), .B(G101), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G3));
  OAI21_X1  g455(.A(new_n305), .B1(new_n267), .B2(new_n219), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n285), .A2(new_n268), .ZN(new_n643));
  AOI211_X1 g457(.A(new_n271), .B(new_n642), .C1(new_n643), .C2(new_n273), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT31), .B1(new_n278), .B2(new_n260), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n286), .A2(new_n287), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT28), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n305), .B1(new_n648), .B2(new_n311), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT72), .B1(new_n646), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n280), .A2(new_n281), .A3(new_n293), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n188), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n300), .B1(new_n294), .B2(new_n295), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n652), .B1(G472), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n441), .A2(new_n444), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(new_n377), .A3(new_n373), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n445), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n472), .A2(new_n493), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n445), .B1(new_n500), .B2(new_n505), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n508), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT101), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n658), .B1(new_n472), .B2(new_n493), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n506), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n665), .A3(new_n508), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n662), .A2(new_n618), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n609), .B1(new_n634), .B2(new_n636), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n572), .A2(G478), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n570), .A2(new_n571), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT33), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT33), .B1(new_n671), .B2(new_n672), .ZN(new_n674));
  OAI211_X1 g488(.A(G478), .B(new_n300), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n668), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n657), .A2(new_n667), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT34), .B(G104), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  OAI21_X1  g494(.A(KEYINPUT98), .B1(new_n575), .B2(new_n576), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n581), .A2(new_n582), .A3(new_n578), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR3_X1    g497(.A1(new_n637), .A2(new_n683), .A3(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n662), .A2(new_n666), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(KEYINPUT104), .B1(new_n637), .B2(new_n683), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n657), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT35), .B(G107), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G9));
  NAND2_X1  g505(.A1(new_n371), .A2(new_n372), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n323), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n355), .A2(new_n359), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n364), .A2(KEYINPUT36), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n376), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n638), .A2(new_n654), .A3(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  AOI22_X1  g515(.A1(new_n692), .A2(new_n323), .B1(new_n376), .B2(new_n696), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n685), .A2(new_n655), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT105), .B(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n611), .B1(new_n615), .B2(new_n704), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n683), .A2(new_n668), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n321), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  XOR2_X1   g522(.A(new_n507), .B(KEYINPUT38), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n584), .A2(new_n668), .ZN(new_n710));
  INV_X1    g524(.A(new_n508), .ZN(new_n711));
  NOR4_X1   g525(.A1(new_n709), .A2(new_n710), .A3(new_n698), .A4(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n302), .A2(new_n205), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n473), .B1(new_n316), .B2(new_n305), .ZN(new_n714));
  OAI21_X1  g528(.A(G472), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n298), .A2(new_n299), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n705), .B(KEYINPUT39), .Z(new_n717));
  NAND3_X1  g531(.A1(new_n441), .A2(new_n444), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n718), .A2(KEYINPUT40), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n712), .A2(new_n716), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G143), .ZN(G45));
  NOR2_X1   g536(.A1(new_n677), .A2(new_n705), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n703), .A2(new_n321), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT106), .B(G146), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G48));
  NOR2_X1   g540(.A1(new_n667), .A2(new_n677), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n300), .B1(new_n428), .B2(new_n431), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(G469), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n444), .A3(new_n432), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n727), .A2(new_n378), .A3(new_n321), .A4(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT41), .B(G113), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT107), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n732), .B(new_n734), .ZN(G15));
  NAND3_X1  g549(.A1(new_n321), .A2(new_n378), .A3(new_n731), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n688), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n208), .ZN(G18));
  AND3_X1   g552(.A1(new_n731), .A2(new_n662), .A3(new_n666), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n702), .A2(new_n584), .A3(new_n637), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n321), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G119), .ZN(G21));
  INV_X1    g556(.A(new_n667), .ZN(new_n743));
  INV_X1    g557(.A(new_n668), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n683), .A3(new_n730), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n318), .A2(new_n205), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n188), .B1(new_n746), .B2(new_n280), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n653), .B2(G472), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n745), .A3(new_n378), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n653), .A2(G472), .ZN(new_n752));
  INV_X1    g566(.A(new_n747), .ZN(new_n753));
  AND4_X1   g567(.A1(new_n751), .A2(new_n752), .A3(new_n698), .A4(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n751), .B1(new_n748), .B2(new_n698), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n723), .B(new_n739), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT109), .B(G125), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n756), .B(new_n757), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n298), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n296), .A2(KEYINPUT110), .A3(new_n297), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(new_n299), .A3(new_n320), .A4(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n677), .A2(new_n705), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n507), .A2(new_n711), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n655), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n762), .A2(new_n765), .A3(new_n378), .A4(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n321), .A2(new_n378), .A3(new_n723), .A4(new_n768), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n764), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  AND4_X1   g587(.A1(new_n378), .A2(new_n321), .A3(new_n706), .A4(new_n768), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(new_n222), .ZN(G36));
  NOR2_X1   g589(.A1(new_n654), .A2(new_n702), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n777));
  INV_X1    g591(.A(new_n676), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n777), .B1(new_n778), .B2(new_n668), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(KEYINPUT43), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n779), .B(KEYINPUT43), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(KEYINPUT44), .A3(new_n776), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n786), .A3(KEYINPUT113), .A4(new_n766), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n435), .B1(new_n437), .B2(new_n438), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n379), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n790), .B2(new_n789), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n440), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n788), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n792), .A2(KEYINPUT111), .A3(KEYINPUT46), .A4(new_n440), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n432), .A4(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(new_n444), .A3(new_n717), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n787), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n767), .B1(new_n782), .B2(new_n783), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT113), .B1(new_n801), .B2(new_n786), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NOR4_X1   g618(.A1(new_n321), .A2(new_n763), .A3(new_n378), .A4(new_n767), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n798), .A2(KEYINPUT47), .A3(new_n444), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT47), .B1(new_n798), .B2(new_n444), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  NAND2_X1  g624(.A1(new_n729), .A2(new_n432), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(KEYINPUT114), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT49), .Z(new_n813));
  INV_X1    g627(.A(new_n716), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n444), .A2(new_n508), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n378), .A2(new_n815), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n744), .A2(new_n816), .A3(new_n676), .A4(new_n709), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n813), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n731), .A2(new_n611), .A3(new_n766), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n785), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n762), .A2(new_n378), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND4_X1   g638(.A1(new_n378), .A2(new_n752), .A3(new_n611), .A4(new_n753), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n785), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n739), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n814), .A2(new_n378), .A3(new_n819), .ZN(new_n828));
  INV_X1    g642(.A(new_n677), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n610), .B(G953), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n824), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n822), .A2(new_n823), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n748), .A2(new_n698), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT108), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n748), .A2(new_n751), .A3(new_n698), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n668), .A2(new_n676), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n820), .A2(new_n838), .B1(new_n828), .B2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n709), .A2(new_n711), .A3(new_n731), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT50), .B1(new_n826), .B2(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(KEYINPUT50), .A2(new_n785), .A3(new_n825), .A4(new_n841), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n812), .A2(new_n444), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n807), .A2(new_n808), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n826), .A2(new_n766), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n844), .A2(new_n845), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n826), .A2(new_n841), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT50), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n843), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(KEYINPUT117), .A3(new_n840), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n834), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n834), .B(new_n840), .C1(new_n847), .C2(new_n849), .ZN(new_n859));
  OR2_X1    g673(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n856), .A2(KEYINPUT116), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n833), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n703), .B(new_n321), .C1(new_n706), .C2(new_n723), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n698), .A2(new_n655), .A3(new_n705), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n685), .A2(new_n710), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n716), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n756), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(KEYINPUT52), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n756), .A2(new_n865), .A3(new_n871), .A4(new_n868), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n763), .B1(new_n836), .B2(new_n837), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n575), .A2(new_n576), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n668), .A2(new_n705), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n321), .A2(new_n876), .A3(new_n698), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n768), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n774), .B1(new_n769), .B2(new_n771), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n507), .A2(new_n618), .A3(new_n508), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n654), .A2(new_n829), .A3(new_n656), .A4(new_n883), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n639), .A2(new_n749), .A3(new_n741), .A4(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n321), .A2(new_n378), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n684), .A2(new_n686), .A3(new_n687), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n886), .B(new_n731), .C1(new_n887), .C2(new_n727), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n882), .A2(new_n668), .A3(new_n876), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n656), .A2(new_n889), .A3(new_n296), .A4(new_n752), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT115), .B1(new_n699), .B2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n699), .A2(new_n890), .A3(KEYINPUT115), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n885), .A2(new_n888), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n881), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n874), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n732), .B1(new_n688), .B2(new_n736), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n699), .A2(KEYINPUT115), .A3(new_n890), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n891), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n885), .A3(new_n880), .A4(new_n879), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n873), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n864), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n874), .A2(new_n895), .A3(KEYINPUT53), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n901), .B1(new_n900), .B2(new_n873), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n905), .A3(KEYINPUT54), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n863), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n818), .B1(new_n907), .B2(new_n908), .ZN(G75));
  NOR2_X1   g723(.A1(new_n198), .A2(G952), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n904), .A2(new_n905), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n912), .A2(new_n562), .A3(new_n446), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n502), .A2(new_n504), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n452), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n505), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT55), .ZN(new_n917));
  OR2_X1    g731(.A1(new_n917), .A2(KEYINPUT56), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n911), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n912), .A2(new_n562), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n445), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n922), .B2(new_n917), .ZN(G51));
  XOR2_X1   g737(.A(new_n440), .B(KEYINPUT57), .Z(new_n924));
  NAND3_X1  g738(.A1(new_n903), .A2(new_n906), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n431), .B2(new_n428), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n921), .A2(new_n792), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n910), .B1(new_n926), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(new_n632), .ZN(new_n929));
  NAND2_X1  g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n921), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n911), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n921), .A2(new_n929), .A3(new_n930), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G60));
  OR2_X1    g748(.A1(new_n673), .A2(new_n674), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n510), .A2(new_n473), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n937), .B(new_n938), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n903), .A2(new_n906), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n903), .A2(KEYINPUT120), .A3(new_n906), .A4(new_n940), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n939), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n903), .A2(new_n906), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n910), .B1(new_n947), .B2(new_n936), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n945), .A2(new_n948), .ZN(G63));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT122), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n904), .B2(new_n905), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n696), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n911), .B1(new_n955), .B2(new_n374), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT61), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n956), .B2(new_n957), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(G66));
  NAND2_X1  g775(.A1(new_n894), .A2(new_n198), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT123), .Z(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n616), .B2(new_n450), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n914), .B1(G898), .B2(new_n198), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G69));
  AOI21_X1  g781(.A(new_n198), .B1(G227), .B2(G900), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n677), .B1(new_n668), .B2(new_n876), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n767), .A2(new_n718), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n886), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n973), .A2(new_n809), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n803), .A2(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n756), .A2(new_n865), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n721), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n612), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n643), .B1(new_n268), .B2(new_n267), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(new_n624), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n969), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(G900), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n984), .B2(new_n198), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n799), .A2(new_n821), .A3(new_n867), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n809), .A2(new_n880), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n976), .B1(new_n800), .B2(new_n802), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT126), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT126), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n990), .B(new_n976), .C1(new_n800), .C2(new_n802), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n987), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n985), .B1(new_n992), .B2(new_n198), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n968), .B1(new_n983), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n979), .A2(new_n803), .A3(new_n974), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n198), .ZN(new_n996));
  INV_X1    g810(.A(new_n982), .ZN(new_n997));
  AOI21_X1  g811(.A(KEYINPUT125), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n968), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n992), .A2(new_n198), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n998), .B(new_n999), .C1(new_n1000), .C2(new_n985), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n994), .A2(new_n1001), .ZN(G72));
  AND2_X1   g816(.A1(new_n302), .A2(new_n205), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n894), .B(new_n987), .C1(new_n989), .C2(new_n991), .ZN(new_n1004));
  NAND2_X1  g818(.A1(G472), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT63), .Z(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1003), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n894), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n979), .A2(new_n1009), .A3(new_n974), .A4(new_n803), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n1006), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n910), .B1(new_n1011), .B2(new_n713), .ZN(new_n1012));
  INV_X1    g826(.A(KEYINPUT127), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n302), .A2(new_n305), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1007), .B1(new_n1015), .B2(new_n270), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n912), .A2(new_n1013), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1013), .B1(new_n912), .B2(new_n1016), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1008), .B(new_n1012), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(G57));
endmodule


