//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT73), .B(G902), .Z(new_n188));
  INV_X1    g002(.A(KEYINPUT28), .ZN(new_n189));
  XOR2_X1   g003(.A(G116), .B(G119), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G113), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n194), .A2(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n196), .B(new_n201), .C1(new_n193), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G134), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G137), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  AND3_X1   g024(.A1(new_n208), .A2(KEYINPUT64), .A3(G137), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT64), .B1(new_n208), .B2(G137), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT11), .B1(new_n208), .B2(G137), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n206), .A3(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n205), .A2(new_n210), .A3(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(KEYINPUT0), .A2(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n202), .A2(new_n203), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n202), .A2(new_n203), .A3(new_n222), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n212), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n218), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G131), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n230), .B2(new_n219), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n192), .B1(new_n220), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n221), .A2(new_n222), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n199), .A2(new_n200), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n224), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND4_X1   g049(.A1(new_n214), .A2(new_n218), .A3(new_n227), .A4(new_n228), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n214), .B1(new_n213), .B2(new_n218), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n192), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n205), .A2(new_n210), .A3(new_n219), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n189), .B1(new_n232), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n189), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT72), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  INV_X1    g063(.A(G237), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n250), .A2(new_n251), .A3(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n249), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT29), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n188), .B1(new_n248), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT30), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n238), .A2(new_n259), .A3(new_n240), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(new_n238), .B2(new_n240), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n192), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n241), .ZN(new_n263));
  INV_X1    g077(.A(new_n255), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT29), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n242), .A2(new_n244), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n255), .B(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n258), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n258), .A3(new_n268), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n187), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n241), .A2(new_n255), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT67), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n241), .A2(new_n276), .A3(new_n255), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n262), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT31), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT68), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n281), .A3(KEYINPUT31), .ZN(new_n282));
  INV_X1    g096(.A(new_n267), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n242), .B2(new_n244), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT30), .B1(new_n220), .B2(new_n231), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n238), .A2(new_n259), .A3(new_n240), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n239), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n241), .A2(new_n276), .A3(new_n255), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT69), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n275), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n262), .A2(new_n275), .A3(new_n292), .A4(new_n277), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT69), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n273), .B1(new_n285), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT32), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n295), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(new_n280), .A3(new_n282), .A4(new_n284), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n273), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n272), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G125), .ZN(new_n305));
  INV_X1    g119(.A(G125), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G140), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n307), .A3(KEYINPUT16), .ZN(new_n308));
  OR3_X1    g122(.A1(new_n306), .A2(KEYINPUT16), .A3(G140), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G146), .ZN(new_n310));
  XNOR2_X1  g124(.A(G125), .B(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n194), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n197), .A2(G119), .ZN(new_n313));
  NAND2_X1  g127(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OR2_X1    g129(.A1(new_n197), .A2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g131(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n313), .B1(new_n318), .B2(new_n314), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n317), .A2(new_n319), .A3(G110), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n316), .A2(new_n313), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT24), .B(G110), .Z(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n310), .B(new_n312), .C1(new_n320), .C2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT75), .B1(new_n317), .B2(new_n319), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G110), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT75), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n322), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n308), .A2(G146), .A3(new_n309), .ZN(new_n330));
  AOI21_X1  g144(.A(G146), .B1(new_n308), .B2(new_n309), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n324), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G137), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n251), .A2(G221), .A3(G234), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n324), .B(new_n336), .C1(new_n328), .C2(new_n332), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n188), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n338), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  INV_X1    g159(.A(G217), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n188), .B2(G234), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n345), .B1(new_n344), .B2(new_n347), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n338), .A2(new_n339), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n347), .A2(G902), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n303), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT9), .B(G234), .ZN(new_n356));
  OAI21_X1  g170(.A(G221), .B1(new_n356), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G104), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G107), .ZN(new_n360));
  OR2_X1    g174(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n361));
  INV_X1    g175(.A(G107), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G104), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n359), .A2(G107), .ZN(new_n366));
  NAND2_X1  g180(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT78), .B1(new_n364), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  AND2_X1   g184(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n361), .B1(new_n363), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n366), .A2(new_n365), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n372), .A2(new_n373), .A3(new_n360), .A4(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n369), .A2(new_n370), .A3(new_n375), .A4(G101), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n235), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n369), .A2(G101), .A3(new_n375), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n364), .A2(new_n368), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n370), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n379), .A2(new_n382), .A3(KEYINPUT79), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT79), .B1(new_n379), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  AOI21_X1  g200(.A(G128), .B1(new_n202), .B2(new_n203), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n202), .A2(new_n203), .A3(G128), .ZN(new_n388));
  INV_X1    g202(.A(new_n193), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n390), .B2(new_n196), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n372), .A2(new_n381), .A3(new_n360), .A4(new_n374), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n363), .A2(new_n360), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(KEYINPUT80), .A3(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n205), .A2(KEYINPUT10), .A3(new_n392), .A4(new_n394), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n201), .B(new_n400), .C1(new_n193), .C2(new_n204), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n396), .A2(new_n399), .B1(new_n386), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n236), .A2(new_n237), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n385), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n404), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n205), .B1(new_n392), .B2(new_n394), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n401), .A2(new_n392), .A3(new_n394), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n406), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT12), .B(new_n406), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(G110), .B(G140), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n251), .A2(G227), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n379), .A2(new_n382), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT79), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n379), .A2(new_n382), .A3(KEYINPUT79), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n377), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n402), .A2(new_n386), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT80), .B1(new_n391), .B2(new_n395), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n397), .A2(new_n398), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n406), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n417), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n405), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n418), .A2(new_n430), .A3(G469), .ZN(new_n431));
  NAND2_X1  g245(.A1(G469), .A2(G902), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n385), .A2(new_n403), .A3(new_n404), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n404), .B1(new_n385), .B2(new_n403), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n417), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n405), .A2(new_n413), .A3(new_n429), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n188), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n358), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n235), .B2(new_n306), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n226), .A2(KEYINPUT83), .A3(G125), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT84), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n390), .A2(new_n306), .A3(new_n196), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n251), .A2(G224), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT85), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n452), .A2(new_n457), .A3(new_n453), .A4(new_n454), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n376), .A2(new_n192), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n383), .B2(new_n384), .ZN(new_n464));
  INV_X1    g278(.A(G113), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n466));
  INV_X1    g280(.A(G116), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(G119), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n465), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(new_n190), .B2(new_n466), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n190), .A2(new_n191), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n395), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n464), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT6), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n464), .A2(new_n473), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n474), .B(KEYINPUT82), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n462), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G902), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n474), .B(KEYINPUT8), .Z(new_n484));
  INV_X1    g298(.A(KEYINPUT5), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n469), .B1(new_n485), .B2(new_n190), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n471), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n484), .B1(new_n487), .B2(new_n395), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n470), .A2(new_n471), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n488), .B1(new_n395), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n448), .A2(new_n449), .A3(new_n454), .ZN(new_n491));
  OR2_X1    g305(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n492));
  NAND2_X1  g306(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n457), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n490), .B(new_n495), .C1(new_n460), .C2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n475), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n483), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n446), .B1(new_n482), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n475), .A2(KEYINPUT6), .B1(new_n477), .B2(new_n478), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n478), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n461), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n499), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n504), .A3(new_n445), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n444), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G475), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n311), .B(new_n194), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n250), .A2(new_n251), .A3(G214), .ZN(new_n509));
  NAND2_X1  g323(.A1(KEYINPUT87), .A2(G143), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(KEYINPUT87), .A2(G143), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(KEYINPUT87), .A2(G143), .ZN(new_n514));
  NOR2_X1   g328(.A1(G237), .A2(G953), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(G214), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT18), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n513), .B(new_n516), .C1(new_n517), .C2(new_n214), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n514), .A2(new_n510), .B1(new_n515), .B2(G214), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n509), .A2(new_n512), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(new_n517), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(G113), .B(G122), .Z(new_n525));
  XOR2_X1   g339(.A(KEYINPUT89), .B(G104), .Z(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT92), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n513), .A2(new_n214), .A3(new_n516), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n522), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n522), .A2(new_n530), .A3(KEYINPUT91), .A4(new_n531), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n330), .B2(new_n331), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n308), .A2(new_n309), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n194), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n310), .A3(KEYINPUT90), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n538), .B(new_n541), .C1(new_n531), .C2(new_n522), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n524), .B(new_n529), .C1(new_n536), .C2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(new_n483), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n524), .B1(new_n536), .B2(new_n542), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n528), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n507), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n527), .B1(new_n519), .B2(new_n523), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n311), .B(KEYINPUT19), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n330), .B1(new_n550), .B2(new_n194), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n551), .A2(new_n552), .B1(new_n522), .B2(new_n530), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n549), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n527), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n545), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  NOR2_X1   g372(.A1(G475), .A2(G902), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n548), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G478), .B1(KEYINPUT97), .B2(KEYINPUT15), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(KEYINPUT97), .B2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n197), .B2(G143), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n197), .A2(G143), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT93), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n198), .A2(G128), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n198), .A2(G128), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n570), .B(new_n571), .C1(new_n572), .C2(new_n566), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(KEYINPUT13), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G134), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT94), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n568), .B2(new_n572), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n197), .A2(G143), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(new_n579), .A3(KEYINPUT94), .ZN(new_n580));
  AOI21_X1  g394(.A(G134), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G116), .B(G122), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(new_n362), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n576), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G122), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G116), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT14), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n467), .A2(G122), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n586), .A2(G116), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n588), .B2(new_n587), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT96), .B1(new_n591), .B2(KEYINPUT14), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n592), .B(G107), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT95), .B1(new_n583), .B2(new_n362), .ZN(new_n597));
  AND4_X1   g411(.A1(KEYINPUT95), .A2(new_n587), .A3(new_n591), .A4(new_n362), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n578), .A2(G134), .A3(new_n580), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n596), .B(new_n599), .C1(new_n600), .C2(new_n581), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n585), .A2(new_n601), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n356), .A2(new_n346), .A3(G953), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n585), .A2(new_n601), .A3(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT98), .B1(new_n607), .B2(new_n188), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n585), .A2(new_n601), .A3(new_n603), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n603), .B1(new_n585), .B2(new_n601), .ZN(new_n610));
  OAI211_X1 g424(.A(KEYINPUT98), .B(new_n188), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n565), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n565), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n609), .A2(new_n610), .ZN(new_n615));
  INV_X1    g429(.A(new_n188), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n614), .B1(new_n617), .B2(KEYINPUT98), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(G952), .ZN(new_n620));
  AOI211_X1 g434(.A(G953), .B(new_n620), .C1(G234), .C2(G237), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n251), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT21), .B(G898), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n563), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n442), .A2(new_n506), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n355), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(G101), .ZN(G3));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n607), .B1(KEYINPUT99), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n630), .B1(new_n607), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n188), .A2(G478), .ZN(new_n633));
  OAI22_X1  g447(.A1(new_n632), .A2(new_n633), .B1(G478), .B2(new_n617), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n563), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(KEYINPUT100), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n563), .B2(new_n634), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n624), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n506), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n187), .B1(new_n300), .B2(new_n188), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n353), .A2(new_n644), .A3(new_n297), .A4(new_n442), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  AOI21_X1  g462(.A(new_n547), .B1(new_n613), .B2(new_n618), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n562), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n555), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n545), .A2(new_n556), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n653), .A3(new_n559), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT20), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n560), .A3(KEYINPUT101), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n651), .A3(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n641), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n645), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT102), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  INV_X1    g476(.A(new_n297), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n337), .A2(KEYINPUT36), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n333), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n333), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n351), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT103), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n348), .A2(new_n349), .A3(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n663), .A2(new_n643), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n626), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT104), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  INV_X1    g488(.A(G900), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n621), .B1(new_n622), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n649), .A2(new_n656), .A3(new_n651), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT105), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n482), .A2(new_n499), .A3(new_n446), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n445), .B1(new_n503), .B2(new_n504), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n443), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI211_X1 g496(.A(G469), .B(new_n616), .C1(new_n437), .C2(new_n438), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n357), .B1(new_n683), .B2(new_n433), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n265), .A2(new_n268), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT71), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n248), .A2(new_n256), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n688), .A3(new_n188), .A4(new_n271), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G472), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n300), .A2(new_n301), .A3(new_n273), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n301), .B1(new_n300), .B2(new_n273), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n669), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n679), .A2(new_n685), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n298), .A2(new_n302), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n669), .B1(new_n697), .B2(new_n690), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n685), .A4(new_n679), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G128), .ZN(G30));
  XOR2_X1   g516(.A(new_n676), .B(KEYINPUT39), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n442), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT108), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT40), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n500), .A2(new_n505), .ZN(new_n709));
  XOR2_X1   g523(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n267), .B1(new_n241), .B2(new_n232), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n275), .B2(new_n290), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n713), .B2(G902), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n691), .B2(new_n692), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n563), .A2(new_n619), .ZN(new_n717));
  NOR4_X1   g531(.A1(new_n716), .A2(new_n444), .A3(new_n694), .A4(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n707), .A2(new_n708), .A3(new_n711), .A4(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G143), .ZN(G45));
  NAND3_X1  g534(.A1(new_n563), .A2(new_n634), .A3(new_n677), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n685), .A2(new_n693), .A3(new_n694), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  INV_X1    g538(.A(new_n438), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n429), .B1(new_n428), .B2(new_n405), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n188), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n441), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n727), .A2(KEYINPUT109), .A3(G469), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n358), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n355), .A2(new_n642), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NAND3_X1  g549(.A1(new_n355), .A2(new_n658), .A3(new_n732), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  INV_X1    g551(.A(new_n732), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n682), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n625), .A3(new_n698), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT110), .B(G119), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G21));
  AOI22_X1  g556(.A1(new_n248), .A2(new_n283), .B1(KEYINPUT31), .B2(new_n278), .ZN(new_n743));
  AOI211_X1 g557(.A(G472), .B(G902), .C1(new_n743), .C2(new_n299), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n354), .A2(new_n643), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n682), .A2(new_n717), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n640), .A4(new_n732), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NOR3_X1   g562(.A1(new_n643), .A2(new_n744), .A3(new_n669), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n506), .A3(new_n732), .A4(new_n722), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n691), .B2(new_n692), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n298), .A2(KEYINPUT111), .A3(new_n302), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n690), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n500), .A2(new_n443), .A3(new_n505), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n756), .A2(new_n684), .A3(new_n757), .A4(new_n721), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n353), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n756), .A2(new_n684), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n693), .A2(new_n353), .A3(new_n760), .A4(new_n722), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n757), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  NAND3_X1  g578(.A1(new_n355), .A2(new_n679), .A3(new_n760), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G134), .ZN(G36));
  INV_X1    g580(.A(new_n563), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n634), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT43), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n768), .B1(KEYINPUT112), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g584(.A(KEYINPUT112), .B(KEYINPUT43), .Z(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n634), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n669), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(new_n663), .B2(new_n643), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n756), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n418), .B2(new_n430), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n440), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n418), .A2(KEYINPUT45), .A3(new_n430), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT46), .B1(new_n780), .B2(new_n432), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n683), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n432), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n358), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n703), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n776), .B(new_n786), .C1(new_n775), .C2(new_n774), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  XNOR2_X1  g602(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  MUX2_X1   g605(.A(new_n789), .B(new_n791), .S(new_n784), .Z(new_n792));
  NOR3_X1   g606(.A1(new_n756), .A2(new_n353), .A3(new_n721), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n303), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT114), .B(G140), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(G42));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n732), .A2(new_n444), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT120), .ZN(new_n799));
  INV_X1    g613(.A(new_n621), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n770), .B2(new_n772), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n745), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n799), .A2(new_n711), .A3(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT50), .Z(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n756), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n357), .B1(new_n730), .B2(new_n731), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n805), .B1(new_n792), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n353), .A2(new_n621), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n738), .A2(new_n715), .A3(new_n756), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT121), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n563), .A2(new_n634), .ZN(new_n811));
  INV_X1    g625(.A(new_n756), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n801), .A2(new_n732), .A3(new_n812), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n810), .A2(new_n811), .B1(new_n749), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n797), .B1(new_n804), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT122), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n804), .A2(new_n815), .A3(new_n797), .ZN(new_n818));
  INV_X1    g632(.A(new_n739), .ZN(new_n819));
  OAI211_X1 g633(.A(G952), .B(new_n251), .C1(new_n819), .C2(new_n802), .ZN(new_n820));
  INV_X1    g634(.A(new_n639), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n755), .A2(new_n353), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n813), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT48), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(KEYINPUT123), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g640(.A(KEYINPUT123), .B(KEYINPUT48), .Z(new_n827));
  OAI211_X1 g641(.A(new_n822), .B(new_n826), .C1(new_n824), .C2(new_n827), .ZN(new_n828));
  OR3_X1    g642(.A1(new_n817), .A2(new_n818), .A3(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n676), .B(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n669), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n684), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n746), .A2(new_n832), .A3(new_n715), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n723), .A2(new_n750), .A3(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n701), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(new_n701), .B2(new_n834), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT118), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n701), .A2(new_n834), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n701), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n619), .A2(new_n547), .A3(new_n676), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n651), .A3(new_n656), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n303), .A2(new_n669), .A3(new_n846), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n643), .A2(new_n669), .A3(new_n744), .A4(new_n721), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n760), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n763), .A2(new_n765), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n740), .A2(new_n733), .A3(new_n736), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n626), .B1(new_n355), .B2(new_n670), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT115), .B1(new_n641), .B2(new_n635), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n854));
  INV_X1    g668(.A(new_n635), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n506), .A2(new_n854), .A3(new_n640), .A4(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n853), .A2(new_n645), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n563), .B1(new_n613), .B2(new_n618), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n506), .A2(new_n640), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT116), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n506), .A2(new_n858), .A3(new_n861), .A4(new_n640), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n645), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n852), .A2(new_n857), .A3(new_n747), .A4(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n850), .A2(new_n851), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT53), .B1(new_n844), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n864), .A2(new_n851), .ZN(new_n867));
  INV_X1    g681(.A(new_n850), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n867), .B(new_n868), .C1(new_n835), .C2(new_n836), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT54), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n835), .A2(new_n836), .A3(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n841), .B1(new_n840), .B2(new_n842), .ZN(new_n874));
  OAI211_X1 g688(.A(KEYINPUT53), .B(new_n865), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n840), .A2(new_n842), .ZN(new_n877));
  AOI211_X1 g691(.A(KEYINPUT119), .B(KEYINPUT53), .C1(new_n877), .C2(new_n865), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n869), .B2(new_n870), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n875), .B(new_n876), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n872), .A2(new_n881), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n829), .A2(new_n882), .B1(G952), .B2(G953), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n354), .A2(new_n768), .A3(new_n444), .A4(new_n358), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n716), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n730), .A2(new_n731), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n711), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n886), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n883), .B1(new_n885), .B2(new_n889), .ZN(G75));
  NAND2_X1  g704(.A1(new_n869), .A2(new_n870), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT119), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n869), .A2(new_n879), .A3(new_n870), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n188), .B1(new_n894), .B2(new_n875), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n446), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n501), .A2(new_n502), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n462), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n503), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT55), .Z(new_n901));
  AND3_X1   g715(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n901), .B1(new_n896), .B2(new_n897), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n251), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(G51));
  XOR2_X1   g719(.A(new_n432), .B(KEYINPUT57), .Z(new_n906));
  AOI21_X1  g720(.A(new_n876), .B1(new_n894), .B2(new_n875), .ZN(new_n907));
  INV_X1    g721(.A(new_n881), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n439), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n895), .A2(new_n779), .A3(new_n778), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(G54));
  NAND3_X1  g726(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n913));
  INV_X1    g727(.A(new_n557), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n914), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n904), .ZN(G60));
  NAND2_X1  g731(.A1(G478), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT59), .Z(new_n919));
  NOR2_X1   g733(.A1(new_n632), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n907), .B2(new_n908), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n922));
  INV_X1    g736(.A(new_n904), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n920), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n875), .B1(new_n878), .B2(new_n880), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT54), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n925), .B1(new_n927), .B2(new_n881), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT124), .B1(new_n928), .B2(new_n904), .ZN(new_n929));
  INV_X1    g743(.A(new_n882), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n632), .B1(new_n930), .B2(new_n919), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n924), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n924), .A2(new_n929), .A3(KEYINPUT125), .A4(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G63));
  XNOR2_X1  g750(.A(KEYINPUT126), .B(KEYINPUT60), .ZN(new_n937));
  NAND2_X1  g751(.A1(G217), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n894), .B2(new_n875), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n665), .A3(new_n666), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n941), .B(new_n923), .C1(new_n350), .C2(new_n940), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT61), .Z(G66));
  INV_X1    g757(.A(G224), .ZN(new_n944));
  OAI21_X1  g758(.A(G953), .B1(new_n623), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n867), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n898), .B1(G898), .B2(new_n251), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G69));
  NAND3_X1  g762(.A1(new_n786), .A2(new_n746), .A3(new_n823), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n794), .A2(new_n787), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n723), .A2(new_n750), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n701), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n950), .A2(new_n763), .A3(new_n765), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(G953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n260), .A2(new_n261), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(new_n550), .Z(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n675), .B2(new_n251), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n719), .A2(new_n701), .A3(new_n951), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n858), .A2(new_n855), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n704), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n355), .A2(new_n812), .A3(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n794), .A2(new_n787), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n960), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n956), .B1(new_n966), .B2(new_n251), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n958), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n251), .B1(G227), .B2(G900), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(G72));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT63), .Z(new_n972));
  INV_X1    g786(.A(new_n867), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n972), .B1(new_n953), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n974), .A2(new_n241), .A3(new_n264), .A4(new_n262), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n966), .B2(new_n973), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n255), .A3(new_n263), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n977), .A3(new_n923), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n866), .A2(new_n871), .ZN(new_n979));
  INV_X1    g793(.A(new_n972), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n263), .A2(new_n264), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n278), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT127), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n978), .B1(new_n979), .B2(new_n983), .ZN(G57));
endmodule


