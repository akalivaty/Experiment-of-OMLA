//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n603, new_n604, new_n605, new_n607, new_n608, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  NOR2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT23), .ZN(new_n204));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT24), .ZN(new_n206));
  INV_X1    g005(.A(G183gat), .ZN(new_n207));
  INV_X1    g006(.A(G190gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT25), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n211), .B(new_n212), .C1(KEYINPUT24), .C2(new_n205), .ZN(new_n213));
  NOR3_X1   g012(.A1(new_n204), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n210), .A2(KEYINPUT64), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT26), .ZN(new_n217));
  OR3_X1    g016(.A1(new_n203), .A2(KEYINPUT66), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT66), .B1(new_n203), .B2(new_n217), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n217), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n212), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT65), .B1(new_n207), .B2(KEYINPUT27), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT27), .B(G183gat), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n208), .B(new_n222), .C1(new_n223), .C2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n223), .A2(KEYINPUT28), .A3(new_n208), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n205), .B(new_n221), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G127gat), .B(G134gat), .Z(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  XOR2_X1   g030(.A(G113gat), .B(G120gat), .Z(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n233), .B(new_n235), .Z(new_n236));
  NOR3_X1   g035(.A1(new_n229), .A2(KEYINPUT68), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n237), .B1(new_n236), .B2(new_n229), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT68), .B1(new_n229), .B2(new_n236), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT33), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G15gat), .B(G43gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT34), .B1(new_n240), .B2(new_n242), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT34), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n238), .A2(new_n249), .A3(new_n241), .A4(new_n239), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n248), .B(new_n250), .C1(new_n243), .C2(new_n246), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT32), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n254), .B1(new_n240), .B2(new_n242), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n252), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n255), .B1(new_n252), .B2(new_n253), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n202), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n261));
  XNOR2_X1  g060(.A(G78gat), .B(G106gat), .ZN(new_n262));
  INV_X1    g061(.A(G50gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT70), .B(G197gat), .ZN(new_n266));
  INV_X1    g065(.A(G204gat), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n266), .A2(new_n267), .ZN(new_n269));
  INV_X1    g068(.A(G211gat), .ZN(new_n270));
  INV_X1    g069(.A(G218gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI22_X1  g071(.A1(new_n268), .A2(new_n269), .B1(KEYINPUT22), .B2(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276));
  XOR2_X1   g075(.A(G141gat), .B(G148gat), .Z(new_n277));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(G155gat), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n280), .A2(G162gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT73), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n277), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT74), .B(G162gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n278), .B1(new_n289), .B2(G155gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n275), .A2(new_n276), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT82), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n291), .A2(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(new_n276), .ZN(new_n298));
  INV_X1    g097(.A(new_n275), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n295), .A2(KEYINPUT82), .ZN(new_n302));
  INV_X1    g101(.A(G228gat), .ZN(new_n303));
  INV_X1    g102(.A(G233gat), .ZN(new_n304));
  OAI22_X1  g103(.A1(new_n301), .A2(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n291), .A2(KEYINPUT3), .ZN(new_n306));
  NOR3_X1   g105(.A1(new_n306), .A2(new_n303), .A3(new_n304), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(new_n292), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G22gat), .ZN(new_n310));
  INV_X1    g109(.A(G22gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n305), .A2(new_n311), .A3(new_n308), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n265), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n265), .A3(new_n312), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n261), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(new_n261), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n317), .A2(new_n318), .A3(new_n313), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT69), .B(KEYINPUT36), .C1(new_n256), .C2(new_n257), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n260), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n316), .A2(new_n319), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(KEYINPUT35), .A3(new_n258), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n229), .A2(new_n276), .ZN(new_n326));
  INV_X1    g125(.A(G226gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n304), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n229), .A2(G226gat), .A3(G233gat), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n328), .A2(new_n275), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n275), .B1(new_n328), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G8gat), .B(G36gat), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT71), .ZN(new_n334));
  XOR2_X1   g133(.A(G64gat), .B(G92gat), .Z(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n332), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT72), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n332), .A2(new_n336), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n341), .B1(new_n338), .B2(new_n337), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT79), .B(KEYINPUT6), .Z(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349));
  OR3_X1    g148(.A1(new_n236), .A2(new_n349), .A3(new_n291), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n236), .B2(new_n291), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n297), .A2(new_n236), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n350), .B(new_n351), .C1(new_n306), .C2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT77), .ZN(new_n356));
  OR3_X1    g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT5), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n355), .B2(KEYINPUT5), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT5), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n236), .B(new_n291), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(new_n354), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n357), .A2(new_n358), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G1gat), .B(G29gat), .Z(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n348), .B1(new_n362), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n348), .A3(new_n367), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n347), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n362), .A2(new_n367), .ZN(new_n372));
  OR2_X1    g171(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(KEYINPUT80), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n347), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n345), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n325), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(new_n370), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n379), .B(new_n346), .C1(new_n380), .C2(new_n368), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n376), .ZN(new_n382));
  INV_X1    g181(.A(new_n332), .ZN(new_n383));
  OR2_X1    g182(.A1(new_n383), .A2(KEYINPUT37), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT38), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n336), .B1(new_n383), .B2(KEYINPUT37), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n337), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n353), .A2(new_n354), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n391), .B(KEYINPUT39), .C1(new_n354), .C2(new_n360), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n392), .B(new_n367), .C1(KEYINPUT39), .C2(new_n391), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT40), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n394), .ZN(new_n395));
  OAI22_X1  g194(.A1(new_n382), .A2(new_n390), .B1(new_n344), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n260), .A2(new_n321), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n398), .A3(new_n323), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT35), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n344), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n323), .A2(new_n258), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n378), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n263), .A2(G43gat), .ZN(new_n405));
  INV_X1    g204(.A(G43gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(G50gat), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT15), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT84), .B(G43gat), .Z(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n263), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n411), .A2(KEYINPUT85), .B1(new_n406), .B2(G50gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(G43gat), .ZN(new_n413));
  OR3_X1    g212(.A1(new_n413), .A2(KEYINPUT85), .A3(G50gat), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT15), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(G36gat), .ZN(new_n416));
  INV_X1    g215(.A(G29gat), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n416), .B1(new_n417), .B2(KEYINPUT14), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n419));
  MUX2_X1   g218(.A(new_n416), .B(new_n418), .S(new_n419), .Z(new_n420));
  OAI21_X1  g219(.A(new_n409), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G8gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G15gat), .B(G22gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT16), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(G1gat), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n422), .B1(new_n425), .B2(KEYINPUT87), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(G1gat), .B2(new_n423), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  OR2_X1    g227(.A1(new_n420), .A2(new_n409), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n411), .A2(KEYINPUT85), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(new_n407), .A3(new_n414), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT15), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n420), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n432), .B(new_n429), .C1(new_n436), .C2(new_n408), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n421), .A2(new_n432), .A3(KEYINPUT17), .A4(new_n429), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n428), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n431), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G229gat), .A2(G233gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(KEYINPUT18), .A3(new_n444), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n421), .A2(new_n429), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n442), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n430), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n444), .B(KEYINPUT13), .Z(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(KEYINPUT88), .A3(new_n452), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n448), .A3(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G113gat), .B(G141gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  XOR2_X1   g260(.A(G169gat), .B(G197gat), .Z(new_n462));
  XNOR2_X1  g261(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT12), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n447), .A2(new_n448), .A3(new_n457), .A4(new_n464), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n404), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT89), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n404), .A2(new_n471), .A3(new_n468), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT94), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT94), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n476), .A2(G99gat), .A3(G106gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n477), .A3(KEYINPUT8), .ZN(new_n478));
  OAI21_X1  g277(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n479));
  AND2_X1   g278(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n482));
  INV_X1    g281(.A(G85gat), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n482), .A2(new_n483), .A3(G92gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n478), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(G99gat), .B(G106gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n478), .B(new_n486), .C1(new_n484), .C2(new_n481), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n491), .B1(new_n439), .B2(new_n440), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(G190gat), .B(G218gat), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT41), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(new_n449), .B2(new_n490), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n493), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n494), .B1(new_n492), .B2(new_n499), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n497), .A2(KEYINPUT41), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n504), .B(KEYINPUT93), .Z(new_n505));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n501), .A2(new_n507), .A3(new_n502), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G57gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT90), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT90), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G57gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n516), .A3(G64gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n513), .A2(G64gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G71gat), .A2(G78gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(G71gat), .A2(G78gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT9), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G64gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(G57gat), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT9), .B1(new_n518), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n521), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n529), .A2(new_n522), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n520), .A2(new_n525), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n428), .B1(KEYINPUT21), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n533), .B2(new_n524), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT90), .B(G57gat), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n518), .B1(new_n535), .B2(G64gat), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n529), .B1(KEYINPUT9), .B2(new_n522), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT21), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XOR2_X1   g339(.A(G127gat), .B(G155gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n532), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT91), .ZN(new_n545));
  XOR2_X1   g344(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G183gat), .B(G211gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT92), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n547), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n543), .B(new_n550), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n512), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n554), .B(new_n555), .Z(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(G230gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n304), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n489), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n482), .A2(new_n483), .ZN(new_n562));
  NAND2_X1  g361(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(G92gat), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n479), .A2(new_n480), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n486), .B1(new_n566), .B2(new_n478), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n538), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n531), .A2(new_n488), .A3(new_n489), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n531), .A2(new_n488), .A3(KEYINPUT95), .A4(new_n489), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT10), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n569), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT10), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT10), .B1(new_n571), .B2(new_n572), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(new_n574), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n560), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n573), .A2(new_n560), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n557), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n582), .B(new_n556), .C1(new_n560), .C2(new_n573), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n553), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n473), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n375), .A2(new_n376), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g393(.A1(new_n473), .A2(new_n345), .A3(new_n588), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT42), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT97), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(new_n424), .ZN(new_n598));
  OR3_X1    g397(.A1(new_n595), .A2(G8gat), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(G8gat), .B1(new_n595), .B2(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n595), .A2(new_n596), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(G1325gat));
  INV_X1    g401(.A(new_n258), .ZN(new_n603));
  OR3_X1    g402(.A1(new_n589), .A2(G15gat), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(G15gat), .B1(new_n589), .B2(new_n398), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(G1326gat));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n320), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT43), .B(G22gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(G1327gat));
  INV_X1    g408(.A(new_n587), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n610), .A2(new_n511), .A3(new_n551), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n611), .B1(new_n470), .B2(new_n472), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n612), .A2(new_n417), .A3(new_n592), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT98), .B(KEYINPUT45), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n404), .A2(new_n616), .A3(new_n511), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n404), .A2(new_n616), .A3(KEYINPUT44), .A4(new_n511), .ZN(new_n620));
  INV_X1    g419(.A(new_n468), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n621), .A2(new_n552), .A3(new_n587), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n619), .A2(new_n592), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n417), .B1(new_n623), .B2(KEYINPUT100), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n624), .B1(KEYINPUT100), .B2(new_n623), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n615), .A2(new_n625), .ZN(G1328gat));
  NAND3_X1  g425(.A1(new_n612), .A2(new_n416), .A3(new_n345), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n627), .A2(KEYINPUT46), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(KEYINPUT46), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n619), .A2(new_n620), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n630), .A2(new_n345), .A3(new_n622), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n628), .B(new_n629), .C1(new_n416), .C2(new_n631), .ZN(G1329gat));
  AOI21_X1  g431(.A(new_n410), .B1(new_n612), .B2(new_n258), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n398), .A2(new_n413), .ZN(new_n634));
  AND4_X1   g433(.A1(new_n620), .A2(new_n619), .A3(new_n622), .A4(new_n634), .ZN(new_n635));
  OR3_X1    g434(.A1(new_n633), .A2(KEYINPUT47), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT47), .B1(new_n633), .B2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(G1330gat));
  INV_X1    g437(.A(KEYINPUT48), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n320), .A2(new_n263), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT101), .Z(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n612), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n619), .A2(new_n320), .A3(new_n620), .A4(new_n622), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT102), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(G50gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(KEYINPUT102), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n643), .A2(G50gat), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n612), .A2(new_n641), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n639), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(G1331gat));
  NAND2_X1  g450(.A1(new_n621), .A2(new_n587), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n553), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n404), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(new_n591), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n535), .ZN(G1332gat));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n404), .A2(KEYINPUT103), .A3(new_n653), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n344), .A2(KEYINPUT104), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n344), .A2(KEYINPUT104), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n662), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT105), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n658), .A2(new_n666), .A3(new_n659), .A4(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1333gat));
  NAND4_X1  g469(.A1(new_n658), .A2(G71gat), .A3(new_n397), .A4(new_n659), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n654), .A2(new_n603), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(G71gat), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT50), .ZN(G1334gat));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n320), .A3(new_n659), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g475(.A1(new_n652), .A2(new_n552), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n630), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(G85gat), .B1(new_n678), .B2(new_n591), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n468), .A2(new_n552), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n404), .A2(new_n511), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT51), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT51), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n404), .A2(new_n683), .A3(new_n511), .A4(new_n680), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n587), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n483), .A3(new_n592), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n679), .A2(new_n687), .ZN(G1336gat));
  NOR2_X1   g487(.A1(new_n662), .A2(G92gat), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT52), .ZN(new_n691));
  INV_X1    g490(.A(new_n662), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n619), .A2(new_n620), .A3(new_n692), .A4(new_n677), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G92gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n690), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n619), .A2(new_n345), .A3(new_n620), .A4(new_n677), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n686), .A2(new_n689), .B1(new_n696), .B2(G92gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n691), .B2(new_n697), .ZN(G1337gat));
  OAI21_X1  g497(.A(G99gat), .B1(new_n678), .B2(new_n398), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n603), .A2(G99gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n685), .B2(new_n700), .ZN(G1338gat));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n323), .A2(G106gat), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n685), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT53), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n619), .A2(new_n320), .A3(new_n620), .A4(new_n677), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G106gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n706), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n709), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT53), .B1(new_n711), .B2(new_n705), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(G1339gat));
  OR2_X1    g512(.A1(new_n580), .A2(new_n574), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n714), .A2(new_n559), .A3(new_n576), .A4(new_n578), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n582), .A2(new_n715), .A3(KEYINPUT54), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT54), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n717), .B(new_n560), .C1(new_n579), .C2(new_n581), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n557), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT107), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n718), .A2(new_n721), .A3(new_n557), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n716), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(new_n724), .A3(KEYINPUT55), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n582), .A2(new_n715), .A3(KEYINPUT54), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n718), .A2(new_n721), .A3(new_n557), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n721), .B1(new_n718), .B2(new_n557), .ZN(new_n728));
  OAI211_X1 g527(.A(KEYINPUT55), .B(new_n726), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n586), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n443), .A2(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n463), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n511), .A2(new_n467), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n731), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT109), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n731), .A2(new_n738), .A3(new_n741), .A4(new_n735), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n731), .A2(new_n468), .A3(new_n735), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n467), .A2(new_n587), .A3(new_n737), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT110), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n511), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n551), .B1(new_n743), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n588), .A2(new_n621), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n591), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n402), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n752), .A2(new_n692), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n468), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n587), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT111), .B(G120gat), .Z(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1341gat));
  NAND2_X1  g557(.A1(new_n753), .A2(new_n552), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G127gat), .ZN(G1342gat));
  NOR4_X1   g559(.A1(new_n752), .A2(G134gat), .A3(new_n345), .A4(new_n512), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT56), .ZN(new_n762));
  INV_X1    g561(.A(new_n753), .ZN(new_n763));
  OAI21_X1  g562(.A(G134gat), .B1(new_n763), .B2(new_n512), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1343gat));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767));
  AOI211_X1 g566(.A(new_n591), .B(new_n322), .C1(new_n748), .C2(new_n749), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n621), .A2(G141gat), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT115), .Z(new_n770));
  AND3_X1   g569(.A1(new_n768), .A2(new_n662), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n692), .A2(new_n591), .A3(new_n397), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n320), .A2(KEYINPUT57), .ZN(new_n773));
  XNOR2_X1  g572(.A(KEYINPUT112), .B(KEYINPUT55), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n732), .B1(new_n733), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n724), .B1(new_n723), .B2(KEYINPUT55), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT113), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n731), .A2(new_n780), .A3(new_n775), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n468), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n511), .B1(new_n782), .B2(new_n745), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n551), .B1(new_n783), .B2(new_n743), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n773), .B1(new_n784), .B2(new_n749), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n748), .A2(new_n749), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT57), .B1(new_n786), .B2(new_n320), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n468), .B(new_n772), .C1(new_n785), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G141gat), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n771), .B1(new_n789), .B2(KEYINPUT114), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n791), .A3(G141gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n767), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n771), .ZN(new_n794));
  XOR2_X1   g593(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n795));
  NAND3_X1  g594(.A1(new_n789), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n766), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n788), .A2(new_n791), .A3(G141gat), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n791), .B1(new_n788), .B2(G141gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n799), .A2(new_n800), .A3(new_n771), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT117), .B(new_n796), .C1(new_n801), .C2(new_n767), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n798), .A2(new_n802), .ZN(G1344gat));
  AND2_X1   g602(.A1(new_n768), .A2(new_n662), .ZN(new_n804));
  INV_X1    g603(.A(G148gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n804), .A2(new_n805), .A3(new_n587), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n772), .B1(new_n785), .B2(new_n787), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n807), .A2(new_n610), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n809), .A3(G148gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT118), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n808), .A2(new_n812), .A3(new_n809), .A4(G148gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n739), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n781), .A2(new_n468), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n780), .B1(new_n731), .B2(new_n775), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n745), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n815), .B1(new_n818), .B2(new_n512), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n749), .B1(new_n819), .B2(new_n552), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT57), .B1(new_n820), .B2(new_n320), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n786), .A2(KEYINPUT57), .A3(new_n320), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n772), .A2(new_n587), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n805), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT119), .B1(new_n824), .B2(new_n825), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n809), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n806), .B1(new_n814), .B2(new_n830), .ZN(G1345gat));
  OAI21_X1  g630(.A(G155gat), .B1(new_n807), .B2(new_n551), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n804), .A2(new_n280), .A3(new_n552), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1346gat));
  NOR3_X1   g633(.A1(new_n345), .A2(new_n289), .A3(new_n512), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n768), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT120), .Z(new_n837));
  OR2_X1    g636(.A1(new_n807), .A2(new_n512), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n289), .B1(new_n838), .B2(new_n839), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n837), .B1(new_n840), .B2(new_n841), .ZN(G1347gat));
  AOI21_X1  g641(.A(new_n592), .B1(new_n748), .B2(new_n749), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n751), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n345), .ZN(new_n845));
  INV_X1    g644(.A(G169gat), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(new_n621), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n692), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(KEYINPUT122), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n468), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n847), .B1(new_n850), .B2(new_n846), .ZN(G1348gat));
  INV_X1    g650(.A(G176gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n852), .A3(new_n587), .ZN(new_n853));
  OAI21_X1  g652(.A(G176gat), .B1(new_n845), .B2(new_n610), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1349gat));
  OAI21_X1  g654(.A(G183gat), .B1(new_n845), .B2(new_n551), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n552), .A2(new_n223), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n848), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g658(.A(G190gat), .B1(new_n845), .B2(new_n512), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT61), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n849), .A2(new_n208), .A3(new_n511), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(G1351gat));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n592), .A2(new_n344), .A3(new_n397), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(new_n745), .ZN(new_n867));
  INV_X1    g666(.A(new_n774), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n586), .B1(new_n723), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n730), .B2(new_n725), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n621), .B1(new_n870), .B2(new_n780), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n867), .B1(new_n871), .B2(new_n779), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n739), .B1(new_n872), .B2(new_n511), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n873), .A2(new_n551), .B1(new_n621), .B2(new_n588), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n866), .B1(new_n874), .B2(new_n323), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT123), .B1(new_n875), .B2(new_n822), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n821), .A2(new_n823), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n468), .B(new_n865), .C1(new_n876), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G197gat), .ZN(new_n880));
  INV_X1    g679(.A(new_n322), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n843), .A2(new_n881), .A3(new_n692), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(G197gat), .A3(new_n621), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n864), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g684(.A(KEYINPUT124), .B(new_n883), .C1(new_n879), .C2(G197gat), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n587), .A2(new_n267), .ZN(new_n888));
  OAI22_X1  g687(.A1(new_n882), .A2(new_n888), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n889));
  NAND2_X1  g688(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n889), .B(new_n890), .Z(new_n891));
  INV_X1    g690(.A(new_n865), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n875), .A2(KEYINPUT123), .A3(new_n822), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n877), .B1(new_n821), .B2(new_n823), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n610), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n891), .B(KEYINPUT126), .C1(new_n895), .C2(new_n267), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n267), .B1(new_n898), .B2(new_n587), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n889), .B(new_n890), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(G1353gat));
  OAI211_X1 g701(.A(new_n552), .B(new_n865), .C1(new_n821), .C2(new_n823), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT63), .B1(new_n903), .B2(G211gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n552), .A2(new_n270), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n904), .A2(new_n905), .B1(new_n882), .B2(new_n906), .ZN(G1354gat));
  INV_X1    g706(.A(KEYINPUT127), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n271), .B1(new_n898), .B2(new_n511), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n882), .A2(G218gat), .A3(new_n512), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n910), .ZN(new_n912));
  AOI211_X1 g711(.A(new_n512), .B(new_n892), .C1(new_n893), .C2(new_n894), .ZN(new_n913));
  OAI211_X1 g712(.A(KEYINPUT127), .B(new_n912), .C1(new_n913), .C2(new_n271), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n911), .A2(new_n914), .ZN(G1355gat));
endmodule


