//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:17 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND4_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT0), .A4(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n190), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(KEYINPUT11), .A3(G134), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G131), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(KEYINPUT65), .A3(G131), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n201), .A2(new_n199), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n208), .A2(KEYINPUT64), .A3(new_n209), .A4(new_n198), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n198), .A2(new_n201), .A3(new_n209), .A4(new_n199), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT64), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n195), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n211), .B(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n192), .A2(new_n217), .A3(G128), .ZN(new_n218));
  INV_X1    g032(.A(new_n199), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n197), .A2(G137), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G128), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n188), .B(new_n190), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n215), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT30), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT2), .B(G113), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G119), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n233), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n228), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n205), .A2(new_n206), .B1(new_n210), .B2(new_n213), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n195), .ZN(new_n241));
  INV_X1    g055(.A(new_n195), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n202), .A2(KEYINPUT65), .A3(G131), .ZN(new_n243));
  AOI21_X1  g057(.A(KEYINPUT65), .B1(new_n202), .B2(G131), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT66), .B(new_n242), .C1(new_n245), .C2(new_n216), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n225), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n227), .B(new_n238), .C1(new_n247), .C2(KEYINPUT30), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n207), .A2(new_n214), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n242), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n218), .A2(new_n223), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n214), .A2(new_n252), .A3(new_n221), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n238), .B(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n250), .A2(new_n253), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n248), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G237), .ZN(new_n261));
  AOI21_X1  g075(.A(G953), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n263), .B(KEYINPUT27), .Z(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT29), .B1(new_n257), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n215), .B2(new_n225), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n253), .B(new_n269), .C1(new_n240), .C2(new_n195), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n255), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT72), .ZN(new_n274));
  INV_X1    g088(.A(new_n238), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n256), .B1(new_n247), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT28), .ZN(new_n277));
  INV_X1    g091(.A(new_n266), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n279), .A3(new_n272), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n274), .A2(new_n277), .A3(new_n278), .A4(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n267), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n278), .A2(KEYINPUT29), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n238), .B(KEYINPUT67), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n215), .B2(new_n225), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n256), .A2(KEYINPUT73), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n226), .A2(new_n287), .A3(new_n255), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(KEYINPUT28), .A3(new_n288), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n274), .A2(new_n283), .A3(new_n280), .A4(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n290), .A2(KEYINPUT74), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(KEYINPUT74), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n282), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G472), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n256), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(new_n266), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n248), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n274), .A2(new_n277), .A3(new_n280), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n266), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n248), .A2(new_n298), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n248), .A2(new_n298), .A3(KEYINPUT69), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(KEYINPUT31), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n296), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI211_X1 g124(.A(KEYINPUT32), .B(new_n296), .C1(new_n302), .C2(new_n307), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n294), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G221), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT9), .B(G234), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT82), .Z(new_n318));
  INV_X1    g132(.A(G469), .ZN(new_n319));
  XNOR2_X1  g133(.A(G110), .B(G140), .ZN(new_n320));
  INV_X1    g134(.A(G227), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(G953), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n320), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G104), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n325), .B2(G107), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  INV_X1    g141(.A(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G104), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(G107), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G101), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n331), .A2(G101), .ZN(new_n334));
  INV_X1    g148(.A(G101), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n326), .A2(new_n329), .A3(new_n335), .A4(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT4), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n333), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n195), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G104), .B(G107), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT83), .B1(new_n341), .B2(new_n335), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n328), .A2(G104), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n330), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G101), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(new_n223), .A3(new_n218), .A4(new_n336), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n348), .A2(KEYINPUT84), .A3(KEYINPUT10), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT10), .B1(new_n348), .B2(KEYINPUT84), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT85), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n207), .B2(new_n214), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n355), .B(new_n340), .C1(new_n349), .C2(new_n350), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n324), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n240), .B(new_n340), .C1(new_n349), .C2(new_n350), .ZN(new_n358));
  INV_X1    g172(.A(new_n348), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n347), .A2(new_n336), .B1(new_n223), .B2(new_n218), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n249), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT12), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT12), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n249), .B(new_n363), .C1(new_n359), .C2(new_n360), .ZN(new_n364));
  AND4_X1   g178(.A1(new_n358), .A2(new_n362), .A3(new_n364), .A4(new_n324), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n319), .B(new_n316), .C1(new_n357), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT86), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n345), .B1(new_n344), .B2(G101), .ZN(new_n368));
  AOI211_X1 g182(.A(KEYINPUT83), .B(new_n335), .C1(new_n343), .C2(new_n330), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n336), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT84), .B1(new_n370), .B2(new_n251), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n348), .A2(KEYINPUT84), .A3(KEYINPUT10), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n355), .B1(new_n375), .B2(new_n340), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n339), .B(new_n353), .C1(new_n373), .C2(new_n374), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n323), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n358), .A2(new_n362), .A3(new_n364), .A4(new_n324), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n380), .A2(new_n381), .A3(new_n319), .A4(new_n316), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n367), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n358), .A2(new_n362), .A3(new_n364), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n323), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n354), .A2(new_n324), .A3(new_n356), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n319), .B1(new_n387), .B2(new_n316), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n318), .B1(new_n383), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G214), .B1(G237), .B2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(G210), .B1(G237), .B2(G902), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n195), .A2(G125), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(G125), .B1(new_n218), .B2(new_n223), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G953), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G224), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n397), .B(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n238), .B(new_n333), .C1(new_n334), .C2(new_n337), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT5), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n402), .B(G113), .C1(new_n403), .C2(new_n236), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n347), .A2(new_n404), .A3(new_n235), .A4(new_n336), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n401), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G110), .B(G122), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n409), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(KEYINPUT87), .A2(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n406), .A2(new_n408), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n399), .A2(KEYINPUT7), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n395), .B2(new_n396), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n394), .B(new_n417), .C1(new_n252), .C2(G125), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n407), .B(KEYINPUT8), .Z(new_n420));
  NAND2_X1  g234(.A1(new_n404), .A2(new_n235), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n370), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(new_n405), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(G902), .B1(new_n424), .B2(new_n410), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n393), .B1(new_n414), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n414), .A2(new_n425), .A3(new_n393), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n392), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n222), .A2(G143), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n430), .A2(KEYINPUT13), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(KEYINPUT13), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n431), .B(new_n432), .C1(G128), .C2(new_n189), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(G134), .ZN(new_n434));
  XNOR2_X1  g248(.A(G128), .B(G143), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n197), .ZN(new_n436));
  XNOR2_X1  g250(.A(G116), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(new_n328), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(new_n328), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT93), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n435), .B(new_n197), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT14), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n232), .A2(KEYINPUT14), .A3(G122), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(G107), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G217), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n314), .A2(new_n450), .A3(G953), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n451), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n439), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n452), .A2(KEYINPUT94), .A3(new_n316), .A4(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n456), .A2(KEYINPUT15), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n455), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT18), .A2(G131), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n260), .A2(G237), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n462));
  OAI211_X1 g276(.A(G214), .B(new_n398), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(new_n189), .ZN(new_n464));
  AOI21_X1  g278(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT88), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n189), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT88), .A3(new_n460), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT89), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n471), .B2(new_n460), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n469), .A2(KEYINPUT89), .A3(new_n470), .A4(new_n459), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G140), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G125), .ZN(new_n479));
  INV_X1    g293(.A(G125), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G140), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(new_n187), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n187), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT79), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(KEYINPUT79), .A3(new_n187), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n473), .A2(new_n477), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n469), .A2(new_n209), .A3(new_n470), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT90), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n471), .A2(G131), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT17), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT90), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n469), .A2(new_n495), .A3(new_n470), .A4(new_n209), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n479), .A2(new_n481), .A3(KEYINPUT16), .ZN(new_n498));
  OR3_X1    g312(.A1(new_n480), .A2(KEYINPUT16), .A3(G140), .ZN(new_n499));
  AOI21_X1  g313(.A(G146), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n499), .A3(G146), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n209), .B1(new_n469), .B2(new_n470), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(KEYINPUT17), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n325), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n490), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n490), .B2(new_n506), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n316), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT92), .B(G475), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G475), .A2(G902), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT91), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n516));
  INV_X1    g330(.A(new_n502), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n482), .B(KEYINPUT19), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(new_n187), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n490), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n508), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n490), .A2(new_n506), .A3(new_n508), .ZN(new_n524));
  AOI211_X1 g338(.A(KEYINPUT20), .B(new_n515), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT20), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n488), .B1(new_n468), .B2(new_n472), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n527), .A2(new_n477), .B1(new_n516), .B2(new_n519), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n524), .B1(new_n508), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n515), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n526), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n458), .B(new_n513), .C1(new_n525), .C2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G952), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G953), .ZN(new_n534));
  INV_X1    g348(.A(G234), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n258), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n316), .B(new_n398), .C1(G234), .C2(G237), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT21), .B(G898), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n532), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n390), .A2(new_n429), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT81), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n230), .A2(G128), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT75), .B1(new_n222), .B2(G119), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n230), .B2(G128), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT23), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT76), .B(G110), .C1(new_n547), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n222), .A2(G119), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n544), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT24), .B(G110), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n551), .B(new_n557), .C1(new_n517), .C2(new_n500), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n549), .A2(KEYINPUT23), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n548), .A3(new_n546), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n544), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT76), .B1(new_n561), .B2(G110), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT77), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n501), .A2(new_n502), .B1(new_n554), .B2(new_n556), .ZN(new_n564));
  INV_X1    g378(.A(new_n562), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT77), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n551), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G110), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n559), .A2(new_n560), .A3(new_n569), .A4(new_n544), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n553), .A2(new_n555), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT78), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n486), .A2(new_n487), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n502), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n313), .A2(new_n535), .A3(G953), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n568), .A2(new_n575), .A3(new_n579), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n316), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n581), .A2(KEYINPUT25), .A3(new_n316), .A4(new_n582), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n585), .A2(KEYINPUT80), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT80), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n583), .A2(new_n588), .A3(new_n584), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n450), .B1(G234), .B2(new_n316), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n543), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n585), .A2(KEYINPUT80), .A3(new_n586), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n593), .A2(KEYINPUT81), .A3(new_n590), .A4(new_n589), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n581), .A2(new_n582), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n590), .A2(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n592), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n312), .A2(new_n542), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  NAND2_X1  g416(.A1(new_n301), .A2(new_n266), .ZN(new_n603));
  INV_X1    g417(.A(new_n300), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n307), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n316), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n308), .B1(new_n606), .B2(G472), .ZN(new_n607));
  INV_X1    g421(.A(new_n540), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n429), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n513), .B1(new_n525), .B2(new_n531), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n452), .A2(new_n611), .A3(new_n454), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT95), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n452), .A2(KEYINPUT95), .A3(new_n611), .A4(new_n454), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n453), .B1(new_n449), .B2(KEYINPUT96), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n449), .A2(KEYINPUT96), .A3(new_n453), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT33), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n316), .A2(G478), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n452), .A2(new_n316), .A3(new_n454), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(G478), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n610), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n609), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n600), .A2(new_n607), .A3(new_n390), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  AOI21_X1  g441(.A(new_n508), .B1(new_n490), .B2(new_n520), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n530), .B1(new_n509), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT20), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n529), .A2(new_n526), .A3(new_n530), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n630), .A2(new_n631), .B1(new_n511), .B2(new_n512), .ZN(new_n632));
  INV_X1    g446(.A(new_n458), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n609), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n600), .A2(new_n607), .A3(new_n390), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n328), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NOR2_X1   g453(.A1(new_n580), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n576), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n597), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT98), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n592), .A2(new_n594), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n542), .A2(new_n607), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  AND3_X1   g461(.A1(new_n644), .A2(new_n390), .A3(new_n429), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n538), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n536), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n634), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n648), .A2(new_n312), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT99), .B(G128), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G30));
  NAND2_X1  g470(.A1(new_n605), .A2(new_n295), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT32), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n308), .A2(new_n309), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n305), .A2(new_n306), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n286), .A2(new_n266), .A3(new_n288), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n663), .B2(G902), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n632), .A2(new_n392), .A3(new_n458), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n592), .A3(new_n594), .A4(new_n643), .ZN(new_n666));
  AOI22_X1  g480(.A1(new_n660), .A2(new_n664), .B1(new_n666), .B2(KEYINPUT100), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n651), .B(KEYINPUT39), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n668), .B1(new_n390), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n388), .B1(new_n367), .B2(new_n382), .ZN(new_n671));
  INV_X1    g485(.A(new_n669), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n671), .A2(KEYINPUT40), .A3(new_n318), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n428), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n426), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n666), .A2(KEYINPUT100), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n667), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NAND3_X1  g494(.A1(new_n610), .A2(new_n622), .A3(new_n651), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n648), .A2(new_n312), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G146), .ZN(G48));
  AOI21_X1  g498(.A(G902), .B1(new_n378), .B2(new_n379), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT101), .B1(new_n685), .B2(new_n319), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n316), .B1(new_n357), .B2(new_n365), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n688), .A3(G469), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n317), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n383), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n686), .A2(new_n689), .B1(new_n367), .B2(new_n382), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT102), .B1(new_n695), .B2(new_n691), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n312), .A3(new_n600), .A4(new_n624), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  NAND4_X1  g514(.A1(new_n697), .A2(new_n312), .A3(new_n600), .A4(new_n635), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G116), .ZN(G18));
  OAI21_X1  g516(.A(new_n391), .B1(new_n674), .B2(new_n426), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n692), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n312), .A2(new_n541), .A3(new_n644), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NAND3_X1  g520(.A1(new_n274), .A2(new_n289), .A3(new_n280), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n266), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n307), .A2(new_n708), .A3(new_n604), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n295), .ZN(new_n710));
  INV_X1    g524(.A(G472), .ZN(new_n711));
  AOI21_X1  g525(.A(G902), .B1(new_n302), .B2(new_n307), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n599), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n632), .A2(new_n703), .A3(new_n458), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n608), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n697), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n606), .A2(G472), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n644), .A2(new_n720), .A3(new_n710), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n682), .A2(new_n691), .A3(new_n429), .A4(new_n695), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n692), .A2(new_n703), .A3(new_n681), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n606), .A2(G472), .B1(new_n295), .B2(new_n709), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(KEYINPUT103), .A3(new_n644), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  NOR2_X1   g542(.A1(new_n319), .A2(new_n316), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n367), .B2(new_n382), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n386), .A2(KEYINPUT104), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n354), .A2(new_n732), .A3(new_n324), .A4(new_n356), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n731), .A2(G469), .A3(new_n385), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT105), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n385), .A2(new_n733), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n736), .A2(new_n737), .A3(G469), .A4(new_n731), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n730), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n675), .A2(new_n391), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n317), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n740), .A2(new_n682), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n312), .A3(new_n600), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT42), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n209), .ZN(G33));
  AOI21_X1  g560(.A(new_n599), .B1(new_n660), .B2(new_n294), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n653), .A2(new_n740), .A3(new_n742), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n630), .A2(new_n631), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n622), .A2(new_n752), .A3(new_n513), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n632), .B(new_n622), .C1(new_n756), .C2(KEYINPUT43), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n644), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n751), .B1(new_n759), .B2(new_n607), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n720), .A2(new_n657), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(KEYINPUT44), .A3(new_n644), .A4(new_n758), .ZN(new_n762));
  INV_X1    g576(.A(new_n741), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n319), .B1(new_n387), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n385), .A4(new_n733), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n729), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n383), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n769), .B(new_n729), .C1(new_n765), .C2(new_n766), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n691), .B(new_n669), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n760), .A2(new_n762), .A3(new_n763), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  OAI21_X1  g588(.A(new_n691), .B1(new_n768), .B2(new_n770), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI211_X1 g591(.A(KEYINPUT47), .B(new_n691), .C1(new_n768), .C2(new_n770), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n599), .A2(new_n682), .A3(new_n763), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n780), .A2(new_n312), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  AND4_X1   g597(.A1(new_n698), .A2(new_n701), .A3(new_n705), .A4(new_n717), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT42), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n744), .B(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n601), .A2(new_n645), .A3(new_n625), .A4(new_n636), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT108), .B1(new_n532), .B2(new_n652), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n632), .A2(new_n790), .A3(new_n458), .A4(new_n651), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n390), .A2(new_n763), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n312), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n743), .A2(new_n725), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n795), .A2(new_n644), .B1(new_n747), .B2(new_n748), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n784), .A2(new_n786), .A3(new_n788), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT109), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n592), .A2(new_n594), .A3(new_n643), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n652), .A2(new_n317), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n429), .A2(new_n610), .A3(new_n633), .A4(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n740), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n664), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n658), .B2(new_n659), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n801), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n804), .A2(new_n740), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n644), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n664), .B1(new_n310), .B2(new_n311), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(KEYINPUT109), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n648), .B(new_n312), .C1(new_n653), .C2(new_n682), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n727), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT110), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n800), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n815), .A2(new_n816), .A3(new_n800), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n798), .B(new_n799), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n727), .A2(new_n814), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n804), .A2(new_n740), .ZN(new_n821));
  AND4_X1   g635(.A1(KEYINPUT109), .A2(new_n811), .A3(new_n821), .A4(new_n802), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT109), .B1(new_n810), .B2(new_n811), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT52), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n813), .A2(new_n800), .A3(new_n727), .A4(new_n814), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT53), .B1(new_n827), .B2(new_n797), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n811), .A2(new_n599), .ZN(new_n831));
  INV_X1    g645(.A(new_n692), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n763), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n536), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n835), .A2(new_n610), .A3(new_n622), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n758), .A2(new_n537), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  INV_X1    g652(.A(new_n721), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n838), .A2(KEYINPUT113), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(KEYINPUT112), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n837), .A2(new_n599), .A3(new_n713), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n391), .B1(KEYINPUT112), .B2(new_n845), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n832), .A2(new_n676), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n846), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n836), .A2(new_n844), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n695), .A2(new_n318), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n763), .B1(new_n779), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n850), .A2(new_n846), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n848), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n830), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n838), .A2(new_n747), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT48), .Z(new_n859));
  NAND2_X1  g673(.A1(new_n847), .A2(new_n704), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(new_n534), .C1(new_n835), .C2(new_n623), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n852), .A2(new_n830), .A3(new_n856), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n827), .A2(new_n797), .A3(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n784), .A2(new_n786), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n796), .A2(new_n788), .A3(KEYINPUT111), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT111), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n312), .A2(new_n792), .B1(new_n743), .B2(new_n725), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n749), .B1(new_n871), .B2(new_n802), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n870), .B1(new_n872), .B2(new_n787), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n868), .B(new_n874), .C1(new_n818), .C2(new_n817), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n866), .B1(KEYINPUT53), .B2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n829), .B(new_n865), .C1(new_n876), .C2(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n533), .A2(new_n398), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n676), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n880), .A2(new_n318), .A3(new_n392), .A4(new_n753), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n695), .B(KEYINPUT49), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n831), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT107), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n879), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT114), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n879), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n398), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n815), .A2(new_n816), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT52), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n815), .A2(new_n816), .A3(new_n800), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n867), .B1(new_n873), .B2(new_n869), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n799), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n897), .A2(new_n316), .A3(new_n866), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n898), .B2(G210), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n411), .A2(new_n413), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(new_n400), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n891), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n899), .B2(new_n903), .ZN(G51));
  XNOR2_X1  g719(.A(new_n729), .B(KEYINPUT57), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n897), .A2(new_n907), .A3(new_n866), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n875), .A2(KEYINPUT53), .ZN(new_n909));
  INV_X1    g723(.A(new_n866), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT54), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n906), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n380), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n898), .A2(new_n766), .A3(new_n765), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n890), .B1(new_n913), .B2(new_n914), .ZN(G54));
  AND2_X1   g729(.A1(KEYINPUT58), .A2(G475), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n876), .A2(G902), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n529), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n898), .A2(new_n529), .A3(new_n916), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n891), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT115), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT115), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n919), .A2(new_n920), .A3(new_n923), .A4(new_n891), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(G60));
  OAI21_X1  g739(.A(new_n907), .B1(new_n897), .B2(new_n866), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n926), .A2(new_n829), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  OAI21_X1  g743(.A(new_n619), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n619), .A2(new_n929), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n931), .B1(new_n908), .B2(new_n911), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT116), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n933), .A3(new_n891), .ZN(new_n934));
  INV_X1    g748(.A(new_n931), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n909), .A2(KEYINPUT54), .A3(new_n910), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n926), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT116), .B1(new_n937), .B2(new_n890), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n930), .A2(new_n934), .A3(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT60), .Z(new_n941));
  NAND4_X1  g755(.A1(new_n909), .A2(new_n910), .A3(new_n641), .A4(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n909), .A2(new_n910), .A3(new_n941), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n891), .B(new_n942), .C1(new_n943), .C2(new_n596), .ZN(new_n944));
  NAND2_X1  g758(.A1(KEYINPUT117), .A2(KEYINPUT61), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT117), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n876), .A2(new_n941), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n890), .B1(new_n950), .B2(new_n595), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n951), .A2(new_n946), .A3(new_n947), .A4(new_n942), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n949), .A2(new_n952), .ZN(G66));
  INV_X1    g767(.A(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n539), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n784), .A2(new_n788), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n900), .B1(G898), .B2(new_n398), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G69));
  OAI21_X1  g773(.A(new_n227), .B1(new_n247), .B2(KEYINPUT30), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n518), .ZN(new_n961));
  XOR2_X1   g775(.A(KEYINPUT118), .B(KEYINPUT119), .Z(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n773), .A2(new_n782), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n747), .A2(new_n715), .A3(new_n772), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n820), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n786), .A2(new_n967), .A3(new_n749), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n786), .B2(new_n749), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n398), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n321), .A2(G900), .A3(G953), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n963), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n741), .B1(new_n634), .B2(new_n623), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n747), .A2(new_n390), .A3(new_n669), .A4(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n773), .A2(new_n782), .A3(new_n976), .ZN(new_n977));
  AND3_X1   g791(.A1(new_n679), .A2(new_n727), .A3(new_n814), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n679), .A2(new_n727), .A3(new_n814), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n981), .A2(KEYINPUT120), .A3(KEYINPUT62), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT120), .B1(new_n981), .B2(KEYINPUT62), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n974), .B1(new_n984), .B2(G953), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n973), .B1(new_n963), .B2(new_n985), .ZN(G72));
  XNOR2_X1  g800(.A(KEYINPUT122), .B(KEYINPUT63), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n711), .A2(new_n316), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n956), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n990), .B1(new_n970), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n257), .B(KEYINPUT124), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n266), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n257), .A2(new_n266), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n661), .B1(KEYINPUT126), .B2(new_n997), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n989), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n819), .A2(new_n828), .A3(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n995), .A2(new_n891), .A3(new_n1001), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n980), .B(new_n956), .C1(new_n982), .C2(new_n983), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n990), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT123), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1003), .A2(KEYINPUT123), .A3(new_n990), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n993), .A2(new_n278), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  AND4_X1   g823(.A1(KEYINPUT125), .A2(new_n1006), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1008), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1011));
  AOI21_X1  g825(.A(KEYINPUT125), .B1(new_n1011), .B2(new_n1007), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1002), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(KEYINPUT127), .B(new_n1002), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(G57));
endmodule


