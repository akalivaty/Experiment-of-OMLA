

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797;

  INV_X1 U372 ( .A(n504), .ZN(n355) );
  XNOR2_X1 U373 ( .A(n649), .B(KEYINPUT33), .ZN(n723) );
  XNOR2_X1 U374 ( .A(KEYINPUT6), .B(n618), .ZN(n668) );
  INV_X1 U375 ( .A(n673), .ZN(n690) );
  XNOR2_X1 U376 ( .A(n617), .B(n369), .ZN(n406) );
  XNOR2_X1 U377 ( .A(n562), .B(G146), .ZN(n356) );
  XNOR2_X1 U378 ( .A(G113), .B(G143), .ZN(n593) );
  XNOR2_X1 U379 ( .A(G146), .B(G125), .ZN(n579) );
  NAND2_X2 U380 ( .A1(n477), .A2(n655), .ZN(n511) );
  AND2_X2 U381 ( .A1(n458), .A2(n465), .ZN(n464) );
  AND2_X4 U382 ( .A1(n354), .A2(n353), .ZN(n755) );
  INV_X1 U383 ( .A(n772), .ZN(n353) );
  XNOR2_X2 U384 ( .A(n505), .B(n355), .ZN(n354) );
  XNOR2_X1 U385 ( .A(n561), .B(n356), .ZN(n573) );
  XNOR2_X1 U386 ( .A(n361), .B(n616), .ZN(n696) );
  XNOR2_X1 U387 ( .A(n696), .B(n486), .ZN(n618) );
  NOR2_X2 U388 ( .A1(n685), .A2(n769), .ZN(n686) );
  XNOR2_X1 U389 ( .A(n485), .B(G107), .ZN(n604) );
  XNOR2_X2 U390 ( .A(n488), .B(G128), .ZN(n404) );
  XNOR2_X2 U391 ( .A(n521), .B(KEYINPUT32), .ZN(n793) );
  NOR2_X2 U392 ( .A1(n440), .A2(n373), .ZN(n521) );
  NOR2_X1 U393 ( .A1(n730), .A2(G902), .ZN(n617) );
  NOR2_X1 U394 ( .A1(n734), .A2(n746), .ZN(n663) );
  NAND2_X1 U395 ( .A1(n690), .A2(n691), .ZN(n687) );
  XNOR2_X1 U396 ( .A(n574), .B(G469), .ZN(n627) );
  XNOR2_X1 U397 ( .A(n661), .B(KEYINPUT31), .ZN(n746) );
  NOR2_X1 U398 ( .A1(n627), .A2(n687), .ZN(n662) );
  INV_X2 U399 ( .A(G143), .ZN(n488) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n595) );
  AND2_X1 U401 ( .A1(n458), .A2(n527), .ZN(n467) );
  BUF_X1 U402 ( .A(n796), .Z(n360) );
  NOR2_X1 U403 ( .A1(n745), .A2(n366), .ZN(n448) );
  NOR2_X1 U404 ( .A1(G902), .A2(n762), .ZN(n603) );
  INV_X2 U405 ( .A(G116), .ZN(n485) );
  INV_X2 U406 ( .A(G953), .ZN(n784) );
  INV_X1 U407 ( .A(KEYINPUT106), .ZN(n486) );
  NAND2_X1 U408 ( .A1(n357), .A2(n681), .ZN(n754) );
  NAND2_X1 U409 ( .A1(n359), .A2(n358), .ZN(n357) );
  INV_X1 U410 ( .A(n679), .ZN(n359) );
  INV_X1 U411 ( .A(n783), .ZN(n358) );
  NAND2_X1 U412 ( .A1(n386), .A2(n384), .ZN(n535) );
  XNOR2_X1 U413 ( .A(n499), .B(n498), .ZN(n698) );
  XNOR2_X1 U414 ( .A(n363), .B(KEYINPUT107), .ZN(n707) );
  XNOR2_X1 U415 ( .A(n603), .B(n602), .ZN(n419) );
  BUF_X1 U416 ( .A(n775), .Z(n405) );
  XNOR2_X1 U417 ( .A(n493), .B(n780), .ZN(n762) );
  OR2_X1 U418 ( .A1(n680), .A2(n437), .ZN(n681) );
  XNOR2_X1 U419 ( .A(n517), .B(n552), .ZN(n566) );
  INV_X1 U420 ( .A(G101), .ZN(n478) );
  XNOR2_X1 U421 ( .A(G113), .B(G101), .ZN(n551) );
  NOR2_X1 U422 ( .A1(n730), .A2(G902), .ZN(n361) );
  XOR2_X2 U423 ( .A(G122), .B(G104), .Z(n470) );
  XNOR2_X1 U424 ( .A(n520), .B(G110), .ZN(n482) );
  XNOR2_X1 U425 ( .A(n420), .B(n599), .ZN(n493) );
  BUF_X1 U426 ( .A(n604), .Z(n362) );
  XNOR2_X2 U427 ( .A(n643), .B(KEYINPUT19), .ZN(n477) );
  XNOR2_X1 U428 ( .A(n604), .B(n482), .ZN(n481) );
  XNOR2_X1 U429 ( .A(n519), .B(n566), .ZN(n775) );
  XNOR2_X1 U430 ( .A(n481), .B(n470), .ZN(n519) );
  INV_X1 U431 ( .A(KEYINPUT30), .ZN(n454) );
  INV_X1 U432 ( .A(KEYINPUT109), .ZN(n568) );
  XNOR2_X1 U433 ( .A(n586), .B(n529), .ZN(n673) );
  XNOR2_X1 U434 ( .A(n585), .B(n587), .ZN(n529) );
  NOR2_X1 U435 ( .A1(G902), .A2(n767), .ZN(n586) );
  XNOR2_X1 U436 ( .A(n409), .B(n407), .ZN(n608) );
  XNOR2_X1 U437 ( .A(KEYINPUT8), .B(KEYINPUT66), .ZN(n409) );
  NOR2_X1 U438 ( .A1(n408), .A2(G953), .ZN(n407) );
  INV_X1 U439 ( .A(G234), .ZN(n408) );
  XNOR2_X1 U440 ( .A(n421), .B(n423), .ZN(n420) );
  INV_X1 U441 ( .A(KEYINPUT39), .ZN(n490) );
  NAND2_X1 U442 ( .A1(KEYINPUT47), .A2(n398), .ZN(n397) );
  INV_X1 U443 ( .A(KEYINPUT69), .ZN(n398) );
  AND2_X1 U444 ( .A1(n392), .A2(n641), .ZN(n391) );
  INV_X1 U445 ( .A(KEYINPUT44), .ZN(n413) );
  XNOR2_X1 U446 ( .A(G131), .B(G140), .ZN(n597) );
  XNOR2_X1 U447 ( .A(G104), .B(G110), .ZN(n427) );
  INV_X1 U448 ( .A(KEYINPUT48), .ZN(n647) );
  XNOR2_X1 U449 ( .A(n489), .B(n380), .ZN(n442) );
  OR2_X1 U450 ( .A1(G237), .A2(G902), .ZN(n569) );
  AND2_X1 U451 ( .A1(n703), .A2(n454), .ZN(n451) );
  AND2_X1 U452 ( .A1(n673), .A2(n410), .ZN(n626) );
  NOR2_X1 U453 ( .A1(n411), .A2(n615), .ZN(n410) );
  XNOR2_X1 U454 ( .A(n627), .B(KEYINPUT1), .ZN(n688) );
  XOR2_X1 U455 ( .A(G478), .B(n611), .Z(n633) );
  NOR2_X1 U456 ( .A1(n764), .A2(G902), .ZN(n611) );
  INV_X1 U457 ( .A(KEYINPUT94), .ZN(n544) );
  BUF_X1 U458 ( .A(n696), .Z(n495) );
  XNOR2_X1 U459 ( .A(n506), .B(KEYINPUT103), .ZN(n606) );
  INV_X1 U460 ( .A(KEYINPUT9), .ZN(n506) );
  XNOR2_X1 U461 ( .A(n425), .B(n572), .ZN(n445) );
  INV_X1 U462 ( .A(KEYINPUT81), .ZN(n504) );
  INV_X1 U463 ( .A(n635), .ZN(n503) );
  INV_X1 U464 ( .A(KEYINPUT70), .ZN(n590) );
  INV_X1 U465 ( .A(KEYINPUT22), .ZN(n461) );
  INV_X1 U466 ( .A(G475), .ZN(n600) );
  XNOR2_X1 U467 ( .A(n581), .B(n582), .ZN(n767) );
  INV_X1 U468 ( .A(KEYINPUT125), .ZN(n484) );
  XNOR2_X1 U469 ( .A(n640), .B(KEYINPUT76), .ZN(n392) );
  NAND2_X1 U470 ( .A1(n367), .A2(n395), .ZN(n394) );
  OR2_X1 U471 ( .A1(n664), .A2(KEYINPUT69), .ZN(n395) );
  AND2_X1 U472 ( .A1(n742), .A2(n397), .ZN(n389) );
  XNOR2_X1 U473 ( .A(n702), .B(KEYINPUT77), .ZN(n664) );
  XNOR2_X1 U474 ( .A(n584), .B(n496), .ZN(n588) );
  XNOR2_X1 U475 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n496) );
  XNOR2_X1 U476 ( .A(n385), .B(n494), .ZN(n384) );
  INV_X1 U477 ( .A(KEYINPUT85), .ZN(n494) );
  XNOR2_X1 U478 ( .A(G137), .B(G134), .ZN(n562) );
  XNOR2_X1 U479 ( .A(n448), .B(n447), .ZN(n702) );
  INV_X1 U480 ( .A(KEYINPUT105), .ZN(n447) );
  XNOR2_X1 U481 ( .A(G116), .B(G131), .ZN(n563) );
  INV_X1 U482 ( .A(KEYINPUT16), .ZN(n520) );
  XNOR2_X1 U483 ( .A(n551), .B(n518), .ZN(n517) );
  INV_X1 U484 ( .A(KEYINPUT3), .ZN(n518) );
  XNOR2_X1 U485 ( .A(n470), .B(n422), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n596), .B(KEYINPUT100), .ZN(n422) );
  INV_X1 U487 ( .A(KEYINPUT99), .ZN(n596) );
  XNOR2_X1 U488 ( .A(n424), .B(n430), .ZN(n423) );
  INV_X1 U489 ( .A(KEYINPUT98), .ZN(n430) );
  XOR2_X1 U490 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n594) );
  INV_X1 U491 ( .A(KEYINPUT73), .ZN(n570) );
  XNOR2_X1 U492 ( .A(n426), .B(n374), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n597), .B(n427), .ZN(n426) );
  XNOR2_X1 U494 ( .A(n370), .B(n579), .ZN(n540) );
  XNOR2_X1 U495 ( .A(n539), .B(n538), .ZN(n537) );
  XNOR2_X1 U496 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n539) );
  XNOR2_X1 U497 ( .A(KEYINPUT89), .B(KEYINPUT87), .ZN(n538) );
  XNOR2_X1 U498 ( .A(n547), .B(KEYINPUT4), .ZN(n548) );
  INV_X1 U499 ( .A(KEYINPUT65), .ZN(n547) );
  AND2_X1 U500 ( .A1(n474), .A2(n492), .ZN(n473) );
  INV_X1 U501 ( .A(n795), .ZN(n492) );
  NAND2_X1 U502 ( .A1(G234), .A2(G237), .ZN(n556) );
  OR2_X1 U503 ( .A1(n703), .A2(n454), .ZN(n450) );
  INV_X1 U504 ( .A(n419), .ZN(n471) );
  XNOR2_X1 U505 ( .A(G128), .B(G110), .ZN(n528) );
  XNOR2_X1 U506 ( .A(G140), .B(KEYINPUT23), .ZN(n434) );
  XNOR2_X1 U507 ( .A(G119), .B(G137), .ZN(n577) );
  XOR2_X1 U508 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n757) );
  INV_X1 U509 ( .A(KEYINPUT28), .ZN(n487) );
  XNOR2_X1 U510 ( .A(n632), .B(n456), .ZN(n722) );
  INV_X1 U511 ( .A(KEYINPUT41), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n619), .B(KEYINPUT111), .ZN(n414) );
  INV_X1 U513 ( .A(KEYINPUT96), .ZN(n498) );
  NAND2_X1 U514 ( .A1(n660), .A2(n495), .ZN(n499) );
  XNOR2_X1 U515 ( .A(n613), .B(n612), .ZN(n745) );
  INV_X1 U516 ( .A(KEYINPUT104), .ZN(n612) );
  NAND2_X1 U517 ( .A1(n471), .A2(n633), .ZN(n613) );
  INV_X1 U518 ( .A(n495), .ZN(n542) );
  XNOR2_X1 U519 ( .A(n509), .B(n508), .ZN(n764) );
  XNOR2_X1 U520 ( .A(n607), .B(n368), .ZN(n508) );
  XNOR2_X1 U521 ( .A(n609), .B(n610), .ZN(n509) );
  NAND2_X1 U522 ( .A1(n388), .A2(G210), .ZN(n491) );
  XNOR2_X1 U523 ( .A(n457), .B(KEYINPUT40), .ZN(n794) );
  INV_X1 U524 ( .A(KEYINPUT114), .ZN(n479) );
  NAND2_X1 U525 ( .A1(n371), .A2(n503), .ZN(n502) );
  AND2_X1 U526 ( .A1(n500), .A2(n460), .ZN(n416) );
  BUF_X1 U527 ( .A(n745), .Z(n417) );
  AND2_X1 U528 ( .A1(n472), .A2(n419), .ZN(n366) );
  XNOR2_X1 U529 ( .A(n766), .B(n483), .ZN(n768) );
  INV_X1 U530 ( .A(KEYINPUT60), .ZN(n512) );
  XNOR2_X1 U531 ( .A(n433), .B(n381), .ZN(n432) );
  AND2_X1 U532 ( .A1(n472), .A2(n471), .ZN(n363) );
  AND2_X1 U533 ( .A1(n525), .A2(n583), .ZN(n364) );
  XNOR2_X1 U534 ( .A(KEYINPUT113), .B(n624), .ZN(n791) );
  INV_X1 U535 ( .A(KEYINPUT82), .ZN(n648) );
  AND2_X1 U536 ( .A1(n449), .A2(n473), .ZN(n365) );
  AND2_X1 U537 ( .A1(n390), .A2(n389), .ZN(n367) );
  XNOR2_X1 U538 ( .A(G134), .B(KEYINPUT7), .ZN(n368) );
  XNOR2_X1 U539 ( .A(n616), .B(n568), .ZN(n369) );
  AND2_X1 U540 ( .A1(G224), .A2(n784), .ZN(n370) );
  AND2_X1 U541 ( .A1(n419), .A2(n633), .ZN(n371) );
  AND2_X1 U542 ( .A1(n531), .A2(n648), .ZN(n372) );
  OR2_X1 U543 ( .A1(n500), .A2(n690), .ZN(n373) );
  XOR2_X1 U544 ( .A(n478), .B(G107), .Z(n374) );
  AND2_X1 U545 ( .A1(n626), .A2(n406), .ZN(n375) );
  BUF_X1 U546 ( .A(n688), .Z(n500) );
  AND2_X1 U547 ( .A1(n453), .A2(n450), .ZN(n376) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(KEYINPUT75), .ZN(n377) );
  XOR2_X1 U549 ( .A(n659), .B(KEYINPUT74), .Z(n378) );
  AND2_X1 U550 ( .A1(KEYINPUT69), .A2(n636), .ZN(n379) );
  XNOR2_X1 U551 ( .A(KEYINPUT46), .B(KEYINPUT83), .ZN(n380) );
  XOR2_X1 U552 ( .A(n753), .B(n752), .Z(n381) );
  XOR2_X1 U553 ( .A(n730), .B(KEYINPUT62), .Z(n382) );
  XOR2_X1 U554 ( .A(n684), .B(n683), .Z(n383) );
  NOR2_X1 U555 ( .A1(G952), .A2(n784), .ZN(n769) );
  INV_X1 U556 ( .A(n769), .ZN(n532) );
  NAND2_X1 U557 ( .A1(n792), .A2(KEYINPUT44), .ZN(n385) );
  XNOR2_X2 U558 ( .A(n462), .B(n378), .ZN(n792) );
  NAND2_X1 U559 ( .A1(n387), .A2(n675), .ZN(n386) );
  XNOR2_X1 U560 ( .A(n674), .B(n413), .ZN(n387) );
  NOR2_X2 U561 ( .A1(n793), .A2(n738), .ZN(n674) );
  NAND2_X1 U562 ( .A1(n388), .A2(G472), .ZN(n534) );
  NAND2_X1 U563 ( .A1(n388), .A2(G478), .ZN(n763) );
  NAND2_X1 U564 ( .A1(n388), .A2(G217), .ZN(n766) );
  NAND2_X1 U565 ( .A1(n388), .A2(G469), .ZN(n433) );
  NOR2_X4 U566 ( .A1(n439), .A2(n755), .ZN(n388) );
  NAND2_X1 U567 ( .A1(n664), .A2(n379), .ZN(n390) );
  AND2_X1 U568 ( .A1(n393), .A2(n391), .ZN(n396) );
  XNOR2_X1 U569 ( .A(n796), .B(KEYINPUT78), .ZN(n393) );
  XNOR2_X2 U570 ( .A(n480), .B(n479), .ZN(n796) );
  NAND2_X1 U571 ( .A1(n396), .A2(n394), .ZN(n507) );
  BUF_X1 U572 ( .A(n477), .Z(n399) );
  NOR2_X1 U573 ( .A1(n688), .A2(n687), .ZN(n660) );
  XNOR2_X1 U574 ( .A(n578), .B(n577), .ZN(n582) );
  XNOR2_X1 U575 ( .A(n401), .B(G146), .ZN(n400) );
  XNOR2_X1 U576 ( .A(n561), .B(n562), .ZN(n401) );
  XNOR2_X1 U577 ( .A(n534), .B(n382), .ZN(n533) );
  XNOR2_X1 U578 ( .A(n767), .B(n484), .ZN(n483) );
  NOR2_X1 U579 ( .A1(n475), .A2(n437), .ZN(n436) );
  NAND2_X1 U580 ( .A1(n436), .A2(n365), .ZN(n505) );
  INV_X1 U581 ( .A(n762), .ZN(n515) );
  BUF_X1 U582 ( .A(n667), .Z(n402) );
  BUF_X1 U583 ( .A(n682), .Z(n403) );
  XNOR2_X1 U584 ( .A(n444), .B(n647), .ZN(n476) );
  BUF_X1 U585 ( .A(n734), .Z(n415) );
  AND2_X1 U586 ( .A1(n412), .A2(n526), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n541), .B(KEYINPUT95), .ZN(n734) );
  XNOR2_X1 U588 ( .A(n658), .B(n377), .ZN(n463) );
  NAND2_X1 U589 ( .A1(n463), .A2(n371), .ZN(n462) );
  XNOR2_X1 U590 ( .A(n446), .B(n536), .ZN(n412) );
  NAND2_X1 U591 ( .A1(n671), .A2(n731), .ZN(n446) );
  INV_X1 U592 ( .A(n406), .ZN(n460) );
  NAND2_X1 U593 ( .A1(n406), .A2(n451), .ZN(n429) );
  NOR2_X1 U594 ( .A1(n406), .A2(n454), .ZN(n452) );
  INV_X1 U595 ( .A(n691), .ZN(n411) );
  OR2_X1 U596 ( .A1(n412), .A2(n526), .ZN(n525) );
  NAND2_X1 U597 ( .A1(n414), .A2(n366), .ZN(n642) );
  NAND2_X1 U598 ( .A1(n791), .A2(KEYINPUT82), .ZN(n474) );
  OR2_X2 U599 ( .A1(n756), .A2(n755), .ZN(n497) );
  NAND2_X1 U600 ( .A1(n431), .A2(n416), .ZN(n672) );
  NAND2_X1 U601 ( .A1(n608), .A2(G221), .ZN(n580) );
  INV_X1 U602 ( .A(n475), .ZN(n438) );
  XNOR2_X1 U603 ( .A(n418), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U604 ( .A1(n533), .A2(n532), .ZN(n418) );
  NAND2_X1 U605 ( .A1(n595), .A2(G214), .ZN(n424) );
  NOR2_X1 U606 ( .A1(n452), .A2(n428), .ZN(n501) );
  NAND2_X1 U607 ( .A1(n429), .A2(n376), .ZN(n428) );
  NAND2_X1 U608 ( .A1(n431), .A2(n459), .ZN(n440) );
  XNOR2_X2 U609 ( .A(n510), .B(n461), .ZN(n431) );
  NOR2_X1 U610 ( .A1(n432), .A2(n769), .ZN(G54) );
  XNOR2_X1 U611 ( .A(n434), .B(KEYINPUT24), .ZN(n435) );
  XNOR2_X1 U612 ( .A(n435), .B(n528), .ZN(n578) );
  NAND2_X1 U613 ( .A1(n438), .A2(n365), .ZN(n783) );
  INV_X1 U614 ( .A(KEYINPUT2), .ZN(n437) );
  INV_X1 U615 ( .A(n754), .ZN(n439) );
  NOR2_X1 U616 ( .A1(n440), .A2(n645), .ZN(n669) );
  AND2_X1 U617 ( .A1(n441), .A2(n750), .ZN(n443) );
  XNOR2_X1 U618 ( .A(n507), .B(n530), .ZN(n441) );
  NAND2_X1 U619 ( .A1(n443), .A2(n442), .ZN(n444) );
  XNOR2_X1 U620 ( .A(n445), .B(n400), .ZN(n751) );
  NAND2_X1 U621 ( .A1(n469), .A2(n468), .ZN(n679) );
  NAND2_X1 U622 ( .A1(n476), .A2(n372), .ZN(n449) );
  INV_X1 U623 ( .A(n615), .ZN(n453) );
  NAND2_X1 U624 ( .A1(n794), .A2(n797), .ZN(n489) );
  XNOR2_X1 U625 ( .A(n455), .B(KEYINPUT42), .ZN(n797) );
  NAND2_X1 U626 ( .A1(n722), .A2(n638), .ZN(n455) );
  NAND2_X1 U627 ( .A1(n625), .A2(n366), .ZN(n457) );
  XNOR2_X1 U628 ( .A(n592), .B(n490), .ZN(n625) );
  AND2_X1 U629 ( .A1(n458), .A2(n525), .ZN(n524) );
  NAND2_X1 U630 ( .A1(n522), .A2(n523), .ZN(n458) );
  INV_X1 U631 ( .A(n668), .ZN(n459) );
  NAND2_X1 U632 ( .A1(n464), .A2(n364), .ZN(n468) );
  AND2_X1 U633 ( .A1(n527), .A2(n678), .ZN(n465) );
  NAND2_X1 U634 ( .A1(n466), .A2(KEYINPUT80), .ZN(n469) );
  NAND2_X1 U635 ( .A1(n467), .A2(n364), .ZN(n466) );
  NAND2_X1 U636 ( .A1(n535), .A2(n676), .ZN(n527) );
  INV_X1 U637 ( .A(n633), .ZN(n472) );
  NOR2_X1 U638 ( .A1(n476), .A2(n648), .ZN(n475) );
  NAND2_X1 U639 ( .A1(n638), .A2(n399), .ZN(n639) );
  NOR2_X2 U640 ( .A1(n634), .A2(n502), .ZN(n480) );
  INV_X1 U641 ( .A(n791), .ZN(n531) );
  XNOR2_X1 U642 ( .A(n375), .B(n487), .ZN(n630) );
  NAND2_X1 U643 ( .A1(n761), .A2(n760), .ZN(n516) );
  XNOR2_X1 U644 ( .A(n545), .B(n544), .ZN(n543) );
  XNOR2_X2 U645 ( .A(n591), .B(n590), .ZN(n634) );
  XNOR2_X1 U646 ( .A(n491), .B(n383), .ZN(n685) );
  XNOR2_X1 U647 ( .A(n775), .B(n553), .ZN(n682) );
  NAND2_X1 U648 ( .A1(n497), .A2(n757), .ZN(n761) );
  XNOR2_X1 U649 ( .A(n516), .B(n515), .ZN(n514) );
  AND2_X2 U650 ( .A1(n501), .A2(n662), .ZN(n591) );
  NAND2_X1 U651 ( .A1(n667), .A2(n666), .ZN(n510) );
  XNOR2_X2 U652 ( .A(n511), .B(n657), .ZN(n667) );
  XNOR2_X1 U653 ( .A(n513), .B(n512), .ZN(G60) );
  NAND2_X1 U654 ( .A1(n514), .A2(n532), .ZN(n513) );
  INV_X1 U655 ( .A(n535), .ZN(n523) );
  NAND2_X1 U656 ( .A1(n524), .A2(n527), .ZN(n772) );
  INV_X1 U657 ( .A(n676), .ZN(n526) );
  XNOR2_X2 U658 ( .A(n404), .B(n548), .ZN(n561) );
  INV_X1 U659 ( .A(KEYINPUT68), .ZN(n530) );
  NAND2_X1 U660 ( .A1(n637), .A2(n703), .ZN(n643) );
  XNOR2_X1 U661 ( .A(n555), .B(n554), .ZN(n637) );
  INV_X1 U662 ( .A(KEYINPUT108), .ZN(n536) );
  XNOR2_X1 U663 ( .A(n540), .B(n537), .ZN(n550) );
  NAND2_X1 U664 ( .A1(n543), .A2(n542), .ZN(n541) );
  NAND2_X1 U665 ( .A1(n667), .A2(n662), .ZN(n545) );
  XNOR2_X1 U666 ( .A(n550), .B(n549), .ZN(n553) );
  AND2_X1 U667 ( .A1(n595), .A2(G210), .ZN(n546) );
  INV_X1 U668 ( .A(KEYINPUT80), .ZN(n678) );
  XNOR2_X1 U669 ( .A(n564), .B(n546), .ZN(n565) );
  XNOR2_X1 U670 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U671 ( .A(n566), .B(n565), .ZN(n567) );
  INV_X1 U672 ( .A(KEYINPUT86), .ZN(n656) );
  XNOR2_X1 U673 ( .A(n573), .B(n567), .ZN(n730) );
  XNOR2_X1 U674 ( .A(n656), .B(KEYINPUT0), .ZN(n657) );
  XNOR2_X1 U675 ( .A(n601), .B(n600), .ZN(n602) );
  INV_X1 U676 ( .A(KEYINPUT35), .ZN(n659) );
  INV_X1 U677 ( .A(n500), .ZN(n645) );
  XNOR2_X1 U678 ( .A(n729), .B(n728), .ZN(G75) );
  XOR2_X1 U679 ( .A(G902), .B(KEYINPUT15), .Z(n583) );
  INV_X1 U680 ( .A(n561), .ZN(n549) );
  XOR2_X1 U681 ( .A(KEYINPUT88), .B(G119), .Z(n552) );
  NOR2_X1 U682 ( .A1(n583), .A2(n682), .ZN(n555) );
  NAND2_X1 U683 ( .A1(G210), .A2(n569), .ZN(n554) );
  INV_X1 U684 ( .A(n637), .ZN(n635) );
  XOR2_X1 U685 ( .A(KEYINPUT38), .B(n635), .Z(n631) );
  XNOR2_X1 U686 ( .A(n556), .B(KEYINPUT14), .ZN(n557) );
  NAND2_X1 U687 ( .A1(G952), .A2(n557), .ZN(n715) );
  NOR2_X1 U688 ( .A1(G953), .A2(n715), .ZN(n653) );
  NAND2_X1 U689 ( .A1(G902), .A2(n557), .ZN(n651) );
  OR2_X1 U690 ( .A1(n784), .A2(n651), .ZN(n558) );
  XNOR2_X1 U691 ( .A(KEYINPUT110), .B(n558), .ZN(n559) );
  NOR2_X1 U692 ( .A1(G900), .A2(n559), .ZN(n560) );
  NOR2_X1 U693 ( .A1(n653), .A2(n560), .ZN(n615) );
  XNOR2_X1 U694 ( .A(n563), .B(KEYINPUT5), .ZN(n564) );
  XNOR2_X1 U695 ( .A(G472), .B(KEYINPUT67), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G214), .A2(n569), .ZN(n703) );
  NAND2_X1 U697 ( .A1(G227), .A2(n784), .ZN(n571) );
  NOR2_X1 U698 ( .A1(n751), .A2(G902), .ZN(n574) );
  XOR2_X1 U699 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n576) );
  XNOR2_X1 U700 ( .A(KEYINPUT25), .B(KEYINPUT93), .ZN(n575) );
  XNOR2_X1 U701 ( .A(n576), .B(n575), .ZN(n587) );
  XNOR2_X1 U702 ( .A(KEYINPUT10), .B(n579), .ZN(n598) );
  XNOR2_X1 U703 ( .A(n580), .B(n598), .ZN(n581) );
  INV_X1 U704 ( .A(n583), .ZN(n680) );
  NAND2_X1 U705 ( .A1(n680), .A2(G234), .ZN(n584) );
  NAND2_X1 U706 ( .A1(G217), .A2(n588), .ZN(n585) );
  NAND2_X1 U707 ( .A1(n588), .A2(G221), .ZN(n589) );
  XOR2_X1 U708 ( .A(KEYINPUT21), .B(n589), .Z(n691) );
  NOR2_X1 U709 ( .A1(n634), .A2(n631), .ZN(n592) );
  XNOR2_X1 U710 ( .A(n594), .B(n593), .ZN(n599) );
  XNOR2_X1 U711 ( .A(n598), .B(n597), .ZN(n780) );
  XNOR2_X1 U712 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n601) );
  XNOR2_X1 U713 ( .A(n362), .B(n404), .ZN(n610) );
  XNOR2_X1 U714 ( .A(G122), .B(KEYINPUT102), .ZN(n605) );
  XNOR2_X1 U715 ( .A(n606), .B(n605), .ZN(n607) );
  NAND2_X1 U716 ( .A1(G217), .A2(n608), .ZN(n609) );
  AND2_X1 U717 ( .A1(n625), .A2(n417), .ZN(n614) );
  XNOR2_X1 U718 ( .A(n614), .B(KEYINPUT116), .ZN(n795) );
  NAND2_X1 U719 ( .A1(n626), .A2(n668), .ZN(n619) );
  NOR2_X1 U720 ( .A1(n645), .A2(n642), .ZN(n620) );
  NAND2_X1 U721 ( .A1(n620), .A2(n703), .ZN(n622) );
  XNOR2_X1 U722 ( .A(KEYINPUT112), .B(KEYINPUT43), .ZN(n621) );
  XNOR2_X1 U723 ( .A(n622), .B(n621), .ZN(n623) );
  NAND2_X1 U724 ( .A1(n623), .A2(n635), .ZN(n624) );
  INV_X1 U725 ( .A(n627), .ZN(n628) );
  XNOR2_X1 U726 ( .A(n628), .B(KEYINPUT115), .ZN(n629) );
  NOR2_X1 U727 ( .A1(n630), .A2(n629), .ZN(n638) );
  INV_X1 U728 ( .A(n631), .ZN(n704) );
  NAND2_X1 U729 ( .A1(n704), .A2(n703), .ZN(n701) );
  NOR2_X1 U730 ( .A1(n707), .A2(n701), .ZN(n632) );
  INV_X1 U731 ( .A(KEYINPUT47), .ZN(n636) );
  INV_X1 U732 ( .A(n639), .ZN(n742) );
  NAND2_X1 U733 ( .A1(n639), .A2(KEYINPUT47), .ZN(n640) );
  NAND2_X1 U734 ( .A1(n702), .A2(KEYINPUT47), .ZN(n641) );
  NOR2_X1 U735 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U736 ( .A(n644), .B(KEYINPUT36), .ZN(n646) );
  NAND2_X1 U737 ( .A1(n646), .A2(n645), .ZN(n750) );
  NAND2_X1 U738 ( .A1(n668), .A2(n660), .ZN(n649) );
  NOR2_X1 U739 ( .A1(G898), .A2(n784), .ZN(n650) );
  XOR2_X1 U740 ( .A(KEYINPUT90), .B(n650), .Z(n777) );
  NOR2_X1 U741 ( .A1(n777), .A2(n651), .ZN(n652) );
  NOR2_X1 U742 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U743 ( .A(KEYINPUT91), .B(n654), .ZN(n655) );
  NAND2_X1 U744 ( .A1(n723), .A2(n402), .ZN(n658) );
  NAND2_X1 U745 ( .A1(n698), .A2(n402), .ZN(n661) );
  XNOR2_X1 U746 ( .A(n663), .B(KEYINPUT97), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(n671) );
  NOR2_X1 U748 ( .A1(n707), .A2(n411), .ZN(n666) );
  XNOR2_X1 U749 ( .A(KEYINPUT84), .B(n669), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n670), .A2(n690), .ZN(n731) );
  NOR2_X1 U751 ( .A1(n690), .A2(n672), .ZN(n738) );
  NAND2_X1 U752 ( .A1(n674), .A2(n792), .ZN(n675) );
  XOR2_X1 U753 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n676) );
  XNOR2_X1 U754 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n684) );
  XNOR2_X1 U755 ( .A(n403), .B(KEYINPUT122), .ZN(n683) );
  XNOR2_X1 U756 ( .A(n686), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U757 ( .A1(n500), .A2(n687), .ZN(n689) );
  XNOR2_X1 U758 ( .A(n689), .B(KEYINPUT50), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U760 ( .A(n692), .B(KEYINPUT49), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U762 ( .A1(n495), .A2(n695), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U764 ( .A(n699), .B(KEYINPUT51), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n700), .A2(n722), .ZN(n712) );
  NOR2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n709) );
  NOR2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U768 ( .A(n705), .B(KEYINPUT120), .ZN(n706) );
  NOR2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n723), .A2(n710), .ZN(n711) );
  NAND2_X1 U772 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U773 ( .A(KEYINPUT52), .B(n713), .Z(n714) );
  NOR2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n721) );
  AND2_X1 U775 ( .A1(n783), .A2(n437), .ZN(n716) );
  XNOR2_X1 U776 ( .A(n716), .B(KEYINPUT79), .ZN(n718) );
  NAND2_X1 U777 ( .A1(n772), .A2(n437), .ZN(n717) );
  NAND2_X1 U778 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n719), .A2(n755), .ZN(n720) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n726) );
  AND2_X1 U781 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U782 ( .A1(n724), .A2(G953), .ZN(n725) );
  AND2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n729) );
  INV_X1 U784 ( .A(KEYINPUT121), .ZN(n727) );
  XNOR2_X1 U785 ( .A(n727), .B(KEYINPUT53), .ZN(n728) );
  XNOR2_X1 U786 ( .A(G101), .B(n731), .ZN(G3) );
  XOR2_X1 U787 ( .A(G104), .B(KEYINPUT117), .Z(n733) );
  NAND2_X1 U788 ( .A1(n415), .A2(n366), .ZN(n732) );
  XNOR2_X1 U789 ( .A(n733), .B(n732), .ZN(G6) );
  XOR2_X1 U790 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n736) );
  NAND2_X1 U791 ( .A1(n415), .A2(n417), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U793 ( .A(G107), .B(n737), .ZN(G9) );
  XOR2_X1 U794 ( .A(G110), .B(n738), .Z(G12) );
  XOR2_X1 U795 ( .A(KEYINPUT29), .B(KEYINPUT118), .Z(n740) );
  NAND2_X1 U796 ( .A1(n742), .A2(n417), .ZN(n739) );
  XNOR2_X1 U797 ( .A(n740), .B(n739), .ZN(n741) );
  XNOR2_X1 U798 ( .A(G128), .B(n741), .ZN(G30) );
  NAND2_X1 U799 ( .A1(n742), .A2(n366), .ZN(n743) );
  XNOR2_X1 U800 ( .A(n743), .B(G146), .ZN(G48) );
  NAND2_X1 U801 ( .A1(n746), .A2(n366), .ZN(n744) );
  XNOR2_X1 U802 ( .A(n744), .B(G113), .ZN(G15) );
  XOR2_X1 U803 ( .A(G116), .B(KEYINPUT119), .Z(n748) );
  NAND2_X1 U804 ( .A1(n746), .A2(n417), .ZN(n747) );
  XNOR2_X1 U805 ( .A(n748), .B(n747), .ZN(G18) );
  XOR2_X1 U806 ( .A(G125), .B(KEYINPUT37), .Z(n749) );
  XNOR2_X1 U807 ( .A(n750), .B(n749), .ZN(G27) );
  XOR2_X1 U808 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n753) );
  XNOR2_X1 U809 ( .A(n751), .B(KEYINPUT123), .ZN(n752) );
  NAND2_X1 U810 ( .A1(n754), .A2(G475), .ZN(n756) );
  NOR2_X1 U811 ( .A1(n756), .A2(n755), .ZN(n759) );
  INV_X1 U812 ( .A(n757), .ZN(n758) );
  NAND2_X1 U813 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U814 ( .A(n764), .B(n763), .ZN(n765) );
  NOR2_X1 U815 ( .A1(n769), .A2(n765), .ZN(G63) );
  NOR2_X1 U816 ( .A1(n769), .A2(n768), .ZN(G66) );
  NAND2_X1 U817 ( .A1(G953), .A2(G224), .ZN(n770) );
  XNOR2_X1 U818 ( .A(KEYINPUT61), .B(n770), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(G898), .ZN(n774) );
  OR2_X1 U820 ( .A1(n772), .A2(G953), .ZN(n773) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n779) );
  XNOR2_X1 U822 ( .A(n405), .B(KEYINPUT126), .ZN(n776) );
  NAND2_X1 U823 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U824 ( .A(n779), .B(n778), .Z(G69) );
  XNOR2_X1 U825 ( .A(n780), .B(KEYINPUT127), .ZN(n782) );
  XOR2_X1 U826 ( .A(n401), .B(n782), .Z(n786) );
  XNOR2_X1 U827 ( .A(n786), .B(n783), .ZN(n785) );
  NAND2_X1 U828 ( .A1(n785), .A2(n784), .ZN(n790) );
  XNOR2_X1 U829 ( .A(G227), .B(n786), .ZN(n787) );
  NAND2_X1 U830 ( .A1(n787), .A2(G900), .ZN(n788) );
  NAND2_X1 U831 ( .A1(n788), .A2(G953), .ZN(n789) );
  NAND2_X1 U832 ( .A1(n790), .A2(n789), .ZN(G72) );
  XOR2_X1 U833 ( .A(G140), .B(n791), .Z(G42) );
  XOR2_X1 U834 ( .A(n792), .B(G122), .Z(G24) );
  XOR2_X1 U835 ( .A(n793), .B(G119), .Z(G21) );
  XNOR2_X1 U836 ( .A(G131), .B(n794), .ZN(G33) );
  XOR2_X1 U837 ( .A(G134), .B(n795), .Z(G36) );
  XNOR2_X1 U838 ( .A(n360), .B(G143), .ZN(G45) );
  XNOR2_X1 U839 ( .A(G137), .B(n797), .ZN(G39) );
endmodule

