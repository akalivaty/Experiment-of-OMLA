

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XNOR2_X2 U555 ( .A(KEYINPUT97), .B(n746), .ZN(n794) );
  XNOR2_X1 U556 ( .A(n769), .B(n768), .ZN(n777) );
  XNOR2_X1 U557 ( .A(n758), .B(KEYINPUT102), .ZN(n770) );
  NOR2_X2 U558 ( .A1(n781), .A2(n779), .ZN(n780) );
  NAND2_X1 U559 ( .A1(n757), .A2(n756), .ZN(n758) );
  OR2_X2 U560 ( .A1(n858), .A2(n725), .ZN(n724) );
  XNOR2_X1 U561 ( .A(n528), .B(n527), .ZN(n627) );
  INV_X1 U562 ( .A(KEYINPUT32), .ZN(n768) );
  NOR2_X1 U563 ( .A1(G1966), .A2(n759), .ZN(n775) );
  BUF_X1 U564 ( .A(n627), .Z(n903) );
  INV_X1 U565 ( .A(KEYINPUT93), .ZN(n529) );
  NAND2_X1 U566 ( .A1(n627), .A2(G138), .ZN(n530) );
  XOR2_X1 U567 ( .A(n780), .B(KEYINPUT106), .Z(n520) );
  AND2_X1 U568 ( .A1(n799), .A2(n798), .ZN(n521) );
  AND2_X1 U569 ( .A1(n523), .A2(n831), .ZN(n522) );
  AND2_X1 U570 ( .A1(n829), .A2(n828), .ZN(n523) );
  NOR2_X1 U571 ( .A1(n786), .A2(n785), .ZN(n524) );
  XNOR2_X1 U572 ( .A(KEYINPUT101), .B(KEYINPUT31), .ZN(n525) );
  XOR2_X1 U573 ( .A(KEYINPUT28), .B(n735), .Z(n526) );
  OR2_X1 U574 ( .A1(n715), .A2(n745), .ZN(n717) );
  INV_X1 U575 ( .A(n771), .ZN(n747) );
  NAND2_X1 U576 ( .A1(n747), .A2(G8), .ZN(n748) );
  OR2_X1 U577 ( .A1(n775), .A2(n748), .ZN(n749) );
  XNOR2_X1 U578 ( .A(KEYINPUT99), .B(KEYINPUT29), .ZN(n737) );
  INV_X1 U579 ( .A(n745), .ZN(n739) );
  INV_X1 U580 ( .A(n739), .ZN(n760) );
  INV_X1 U581 ( .A(KEYINPUT96), .ZN(n711) );
  BUF_X1 U582 ( .A(n759), .Z(n785) );
  NAND2_X1 U583 ( .A1(n745), .A2(G8), .ZN(n746) );
  INV_X1 U584 ( .A(KEYINPUT17), .ZN(n527) );
  AND2_X1 U585 ( .A1(n533), .A2(G2104), .ZN(n567) );
  NOR2_X1 U586 ( .A1(n648), .A2(G651), .ZN(n673) );
  BUF_X1 U587 ( .A(n567), .Z(n904) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n538), .Z(n672) );
  XNOR2_X1 U589 ( .A(n530), .B(n529), .ZN(n532) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n909) );
  NAND2_X1 U591 ( .A1(n909), .A2(G114), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n537) );
  INV_X2 U593 ( .A(G2105), .ZN(n533) );
  NAND2_X1 U594 ( .A1(G102), .A2(n904), .ZN(n535) );
  NOR2_X4 U595 ( .A1(G2104), .A2(n533), .ZN(n907) );
  NAND2_X1 U596 ( .A1(G126), .A2(n907), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X2 U598 ( .A1(n537), .A2(n536), .ZN(G164) );
  INV_X1 U599 ( .A(G651), .ZN(n541) );
  NOR2_X1 U600 ( .A1(G543), .A2(n541), .ZN(n538) );
  NAND2_X1 U601 ( .A1(G65), .A2(n672), .ZN(n540) );
  XOR2_X1 U602 ( .A(KEYINPUT0), .B(G543), .Z(n648) );
  NAND2_X1 U603 ( .A1(G53), .A2(n673), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n546) );
  NOR2_X1 U605 ( .A1(G543), .A2(G651), .ZN(n666) );
  NAND2_X1 U606 ( .A1(G91), .A2(n666), .ZN(n544) );
  OR2_X1 U607 ( .A1(n541), .A2(n648), .ZN(n542) );
  XOR2_X1 U608 ( .A(KEYINPUT68), .B(n542), .Z(n668) );
  NAND2_X1 U609 ( .A1(G78), .A2(n668), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(G299) );
  NAND2_X1 U612 ( .A1(G64), .A2(n672), .ZN(n548) );
  NAND2_X1 U613 ( .A1(G52), .A2(n673), .ZN(n547) );
  NAND2_X1 U614 ( .A1(n548), .A2(n547), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n666), .A2(G90), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT70), .ZN(n551) );
  NAND2_X1 U617 ( .A1(G77), .A2(n668), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT71), .B(n552), .ZN(n553) );
  XNOR2_X1 U620 ( .A(KEYINPUT9), .B(n553), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(G171) );
  XOR2_X1 U622 ( .A(G2443), .B(G2446), .Z(n557) );
  XNOR2_X1 U623 ( .A(G2427), .B(G2451), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n563) );
  XOR2_X1 U625 ( .A(G2430), .B(G2454), .Z(n559) );
  XNOR2_X1 U626 ( .A(G1341), .B(G1348), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U628 ( .A(G2435), .B(G2438), .Z(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U630 ( .A(n563), .B(n562), .Z(n564) );
  AND2_X1 U631 ( .A1(G14), .A2(n564), .ZN(G401) );
  AND2_X1 U632 ( .A1(G137), .A2(n627), .ZN(n566) );
  AND2_X1 U633 ( .A1(G125), .A2(n907), .ZN(n565) );
  NOR2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n573) );
  INV_X1 U635 ( .A(KEYINPUT23), .ZN(n569) );
  AND2_X2 U636 ( .A1(G101), .A2(n567), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n571) );
  AND2_X1 U638 ( .A1(n909), .A2(G113), .ZN(n570) );
  NOR2_X1 U639 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n575) );
  INV_X1 U641 ( .A(KEYINPUT66), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n710) );
  BUF_X1 U643 ( .A(n710), .Z(G160) );
  AND2_X1 U644 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U645 ( .A(G108), .ZN(G238) );
  INV_X1 U646 ( .A(G120), .ZN(G236) );
  INV_X1 U647 ( .A(G69), .ZN(G235) );
  INV_X1 U648 ( .A(G132), .ZN(G219) );
  INV_X1 U649 ( .A(G82), .ZN(G220) );
  NAND2_X1 U650 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U651 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U652 ( .A(G223), .ZN(n848) );
  NAND2_X1 U653 ( .A1(n848), .A2(G567), .ZN(n577) );
  XOR2_X1 U654 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  XNOR2_X1 U655 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n583) );
  NAND2_X1 U656 ( .A1(G81), .A2(n666), .ZN(n578) );
  XNOR2_X1 U657 ( .A(n578), .B(KEYINPUT12), .ZN(n579) );
  XNOR2_X1 U658 ( .A(n579), .B(KEYINPUT72), .ZN(n581) );
  NAND2_X1 U659 ( .A1(G68), .A2(n668), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U661 ( .A(n583), .B(n582), .ZN(n586) );
  NAND2_X1 U662 ( .A1(n672), .A2(G56), .ZN(n584) );
  XOR2_X1 U663 ( .A(KEYINPUT14), .B(n584), .Z(n585) );
  NOR2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n673), .A2(G43), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n1009) );
  INV_X1 U667 ( .A(n1009), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n589), .A2(G860), .ZN(G153) );
  INV_X1 U669 ( .A(G171), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n599) );
  NAND2_X1 U671 ( .A1(G92), .A2(n666), .ZN(n591) );
  NAND2_X1 U672 ( .A1(G66), .A2(n672), .ZN(n590) );
  NAND2_X1 U673 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U674 ( .A(KEYINPUT74), .B(n592), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n673), .A2(G54), .ZN(n594) );
  NAND2_X1 U676 ( .A1(G79), .A2(n668), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U678 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U679 ( .A(KEYINPUT15), .B(n597), .Z(n858) );
  INV_X1 U680 ( .A(n858), .ZN(n1012) );
  INV_X1 U681 ( .A(G868), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n1012), .A2(n612), .ZN(n598) );
  NAND2_X1 U683 ( .A1(n599), .A2(n598), .ZN(G284) );
  NAND2_X1 U684 ( .A1(G63), .A2(n672), .ZN(n601) );
  NAND2_X1 U685 ( .A1(G51), .A2(n673), .ZN(n600) );
  NAND2_X1 U686 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U687 ( .A(KEYINPUT6), .B(n602), .Z(n610) );
  NAND2_X1 U688 ( .A1(n668), .A2(G76), .ZN(n606) );
  XOR2_X1 U689 ( .A(KEYINPUT75), .B(KEYINPUT4), .Z(n604) );
  NAND2_X1 U690 ( .A1(G89), .A2(n666), .ZN(n603) );
  XNOR2_X1 U691 ( .A(n604), .B(n603), .ZN(n605) );
  NAND2_X1 U692 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U693 ( .A(n607), .B(KEYINPUT76), .ZN(n608) );
  XNOR2_X1 U694 ( .A(KEYINPUT5), .B(n608), .ZN(n609) );
  NAND2_X1 U695 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U696 ( .A(KEYINPUT7), .B(n611), .ZN(G168) );
  XOR2_X1 U697 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U698 ( .A1(G286), .A2(n612), .ZN(n614) );
  NOR2_X1 U699 ( .A1(G868), .A2(G299), .ZN(n613) );
  NOR2_X1 U700 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U701 ( .A(KEYINPUT77), .B(n615), .Z(G297) );
  INV_X1 U702 ( .A(G559), .ZN(n616) );
  NOR2_X1 U703 ( .A1(G860), .A2(n616), .ZN(n617) );
  XNOR2_X1 U704 ( .A(n617), .B(KEYINPUT78), .ZN(n618) );
  NOR2_X1 U705 ( .A1(n1012), .A2(n618), .ZN(n619) );
  XNOR2_X1 U706 ( .A(n619), .B(KEYINPUT79), .ZN(n620) );
  XNOR2_X1 U707 ( .A(n620), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U708 ( .A1(G868), .A2(n1009), .ZN(n623) );
  NAND2_X1 U709 ( .A1(n858), .A2(G868), .ZN(n621) );
  NOR2_X1 U710 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U711 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U712 ( .A1(G123), .A2(n907), .ZN(n624) );
  XNOR2_X1 U713 ( .A(n624), .B(KEYINPUT18), .ZN(n626) );
  NAND2_X1 U714 ( .A1(n909), .A2(G111), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n626), .A2(n625), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G135), .A2(n903), .ZN(n629) );
  NAND2_X1 U717 ( .A1(G99), .A2(n904), .ZN(n628) );
  NAND2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U719 ( .A1(n631), .A2(n630), .ZN(n962) );
  XNOR2_X1 U720 ( .A(n962), .B(G2096), .ZN(n632) );
  XNOR2_X1 U721 ( .A(n632), .B(KEYINPUT80), .ZN(n634) );
  INV_X1 U722 ( .A(G2100), .ZN(n633) );
  NAND2_X1 U723 ( .A1(n634), .A2(n633), .ZN(G156) );
  NAND2_X1 U724 ( .A1(n858), .A2(G559), .ZN(n688) );
  XNOR2_X1 U725 ( .A(n1009), .B(n688), .ZN(n635) );
  NOR2_X1 U726 ( .A1(n635), .A2(G860), .ZN(n644) );
  NAND2_X1 U727 ( .A1(G80), .A2(n668), .ZN(n636) );
  XOR2_X1 U728 ( .A(KEYINPUT81), .B(n636), .Z(n638) );
  NAND2_X1 U729 ( .A1(n666), .A2(G93), .ZN(n637) );
  NAND2_X1 U730 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U731 ( .A(KEYINPUT82), .B(n639), .ZN(n643) );
  NAND2_X1 U732 ( .A1(G67), .A2(n672), .ZN(n641) );
  NAND2_X1 U733 ( .A1(G55), .A2(n673), .ZN(n640) );
  NAND2_X1 U734 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U735 ( .A1(n643), .A2(n642), .ZN(n681) );
  XNOR2_X1 U736 ( .A(n644), .B(n681), .ZN(G145) );
  NAND2_X1 U737 ( .A1(G49), .A2(n673), .ZN(n646) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n645) );
  NAND2_X1 U739 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U740 ( .A1(n672), .A2(n647), .ZN(n650) );
  NAND2_X1 U741 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U742 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U743 ( .A1(n668), .A2(G73), .ZN(n651) );
  XNOR2_X1 U744 ( .A(n651), .B(KEYINPUT2), .ZN(n658) );
  NAND2_X1 U745 ( .A1(G86), .A2(n666), .ZN(n653) );
  NAND2_X1 U746 ( .A1(G48), .A2(n673), .ZN(n652) );
  NAND2_X1 U747 ( .A1(n653), .A2(n652), .ZN(n656) );
  NAND2_X1 U748 ( .A1(G61), .A2(n672), .ZN(n654) );
  XNOR2_X1 U749 ( .A(KEYINPUT83), .B(n654), .ZN(n655) );
  NOR2_X1 U750 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U751 ( .A1(n658), .A2(n657), .ZN(G305) );
  NAND2_X1 U752 ( .A1(G88), .A2(n666), .ZN(n660) );
  NAND2_X1 U753 ( .A1(G75), .A2(n668), .ZN(n659) );
  NAND2_X1 U754 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U755 ( .A(KEYINPUT84), .B(n661), .Z(n665) );
  NAND2_X1 U756 ( .A1(G62), .A2(n672), .ZN(n663) );
  NAND2_X1 U757 ( .A1(G50), .A2(n673), .ZN(n662) );
  AND2_X1 U758 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U759 ( .A1(n665), .A2(n664), .ZN(G303) );
  INV_X1 U760 ( .A(G303), .ZN(G166) );
  NAND2_X1 U761 ( .A1(n666), .A2(G85), .ZN(n667) );
  XOR2_X1 U762 ( .A(KEYINPUT67), .B(n667), .Z(n670) );
  NAND2_X1 U763 ( .A1(G72), .A2(n668), .ZN(n669) );
  NAND2_X1 U764 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U765 ( .A(KEYINPUT69), .B(n671), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G60), .A2(n672), .ZN(n675) );
  NAND2_X1 U767 ( .A1(G47), .A2(n673), .ZN(n674) );
  AND2_X1 U768 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U769 ( .A1(n677), .A2(n676), .ZN(G290) );
  NOR2_X1 U770 ( .A1(G868), .A2(n681), .ZN(n678) );
  XNOR2_X1 U771 ( .A(n678), .B(KEYINPUT87), .ZN(n691) );
  XNOR2_X1 U772 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n680) );
  XNOR2_X1 U773 ( .A(G288), .B(KEYINPUT86), .ZN(n679) );
  XNOR2_X1 U774 ( .A(n680), .B(n679), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n681), .B(n1009), .ZN(n682) );
  XNOR2_X1 U776 ( .A(n682), .B(G305), .ZN(n683) );
  XNOR2_X1 U777 ( .A(n684), .B(n683), .ZN(n686) );
  XNOR2_X1 U778 ( .A(G299), .B(G166), .ZN(n685) );
  XNOR2_X1 U779 ( .A(n686), .B(n685), .ZN(n687) );
  XNOR2_X1 U780 ( .A(n687), .B(G290), .ZN(n854) );
  XNOR2_X1 U781 ( .A(n854), .B(n688), .ZN(n689) );
  NAND2_X1 U782 ( .A1(G868), .A2(n689), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(G295) );
  NAND2_X1 U784 ( .A1(G2084), .A2(G2078), .ZN(n692) );
  XOR2_X1 U785 ( .A(KEYINPUT20), .B(n692), .Z(n693) );
  NAND2_X1 U786 ( .A1(n693), .A2(G2090), .ZN(n694) );
  XNOR2_X1 U787 ( .A(n694), .B(KEYINPUT88), .ZN(n695) );
  XNOR2_X1 U788 ( .A(KEYINPUT21), .B(n695), .ZN(n696) );
  NAND2_X1 U789 ( .A1(G2072), .A2(n696), .ZN(G158) );
  XOR2_X1 U790 ( .A(KEYINPUT89), .B(G44), .Z(n697) );
  XNOR2_X1 U791 ( .A(KEYINPUT3), .B(n697), .ZN(G218) );
  NOR2_X1 U792 ( .A1(G220), .A2(G219), .ZN(n698) );
  XOR2_X1 U793 ( .A(KEYINPUT22), .B(n698), .Z(n699) );
  NOR2_X1 U794 ( .A1(G218), .A2(n699), .ZN(n700) );
  NAND2_X1 U795 ( .A1(G96), .A2(n700), .ZN(n852) );
  NAND2_X1 U796 ( .A1(n852), .A2(G2106), .ZN(n706) );
  NOR2_X1 U797 ( .A1(G235), .A2(G236), .ZN(n701) );
  XNOR2_X1 U798 ( .A(KEYINPUT90), .B(n701), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n702), .A2(G57), .ZN(n703) );
  NOR2_X1 U800 ( .A1(n703), .A2(G238), .ZN(n704) );
  XNOR2_X1 U801 ( .A(n704), .B(KEYINPUT91), .ZN(n853) );
  NAND2_X1 U802 ( .A1(n853), .A2(G567), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n927) );
  NAND2_X1 U804 ( .A1(G661), .A2(G483), .ZN(n707) );
  NOR2_X1 U805 ( .A1(n927), .A2(n707), .ZN(n851) );
  NAND2_X1 U806 ( .A1(G36), .A2(n851), .ZN(n708) );
  XNOR2_X1 U807 ( .A(n708), .B(KEYINPUT92), .ZN(G176) );
  INV_X1 U808 ( .A(G2067), .ZN(n715) );
  NOR2_X1 U809 ( .A1(G164), .A2(G1384), .ZN(n709) );
  XNOR2_X1 U810 ( .A(n709), .B(KEYINPUT65), .ZN(n802) );
  AND2_X2 U811 ( .A1(n710), .A2(G40), .ZN(n801) );
  XNOR2_X1 U812 ( .A(n801), .B(n711), .ZN(n712) );
  NOR2_X2 U813 ( .A1(n802), .A2(n712), .ZN(n714) );
  INV_X1 U814 ( .A(KEYINPUT64), .ZN(n713) );
  XNOR2_X2 U815 ( .A(n714), .B(n713), .ZN(n745) );
  NAND2_X1 U816 ( .A1(n745), .A2(G1348), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U818 ( .A(n718), .B(KEYINPUT98), .Z(n725) );
  AND2_X1 U819 ( .A1(n739), .A2(G1996), .ZN(n719) );
  XOR2_X1 U820 ( .A(n719), .B(KEYINPUT26), .Z(n722) );
  AND2_X1 U821 ( .A1(n760), .A2(G1341), .ZN(n720) );
  NOR2_X1 U822 ( .A1(n720), .A2(n1009), .ZN(n721) );
  AND2_X1 U823 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U824 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U825 ( .A1(n725), .A2(n858), .ZN(n726) );
  NAND2_X1 U826 ( .A1(n727), .A2(n726), .ZN(n733) );
  INV_X1 U827 ( .A(KEYINPUT27), .ZN(n729) );
  NAND2_X1 U828 ( .A1(G2072), .A2(n739), .ZN(n728) );
  XNOR2_X1 U829 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U830 ( .A1(n760), .A2(G1956), .ZN(n730) );
  NAND2_X1 U831 ( .A1(n731), .A2(n730), .ZN(n734) );
  NOR2_X1 U832 ( .A1(n734), .A2(G299), .ZN(n732) );
  NOR2_X1 U833 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U834 ( .A1(G299), .A2(n734), .ZN(n735) );
  NOR2_X1 U835 ( .A1(n736), .A2(n526), .ZN(n738) );
  XNOR2_X1 U836 ( .A(n738), .B(n737), .ZN(n743) );
  XOR2_X1 U837 ( .A(G2078), .B(KEYINPUT25), .Z(n991) );
  NAND2_X1 U838 ( .A1(n991), .A2(n739), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n760), .A2(G1961), .ZN(n740) );
  NAND2_X1 U840 ( .A1(n741), .A2(n740), .ZN(n751) );
  NOR2_X1 U841 ( .A1(G301), .A2(n751), .ZN(n742) );
  NOR2_X1 U842 ( .A1(n743), .A2(n742), .ZN(n744) );
  INV_X1 U843 ( .A(n744), .ZN(n757) );
  INV_X1 U844 ( .A(n794), .ZN(n759) );
  NOR2_X1 U845 ( .A1(n760), .A2(G2084), .ZN(n771) );
  XNOR2_X1 U846 ( .A(n749), .B(KEYINPUT30), .ZN(n750) );
  NOR2_X1 U847 ( .A1(G168), .A2(n750), .ZN(n754) );
  NAND2_X1 U848 ( .A1(G301), .A2(n751), .ZN(n752) );
  XOR2_X1 U849 ( .A(KEYINPUT100), .B(n752), .Z(n753) );
  NOR2_X1 U850 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U851 ( .A(n755), .B(n525), .ZN(n756) );
  NAND2_X1 U852 ( .A1(n770), .A2(G286), .ZN(n765) );
  NOR2_X1 U853 ( .A1(G1971), .A2(n785), .ZN(n762) );
  NOR2_X1 U854 ( .A1(n760), .A2(G2090), .ZN(n761) );
  NOR2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U856 ( .A1(n763), .A2(G303), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U858 ( .A(n766), .B(KEYINPUT104), .ZN(n767) );
  NAND2_X1 U859 ( .A1(n767), .A2(G8), .ZN(n769) );
  XOR2_X1 U860 ( .A(n770), .B(KEYINPUT103), .Z(n773) );
  NAND2_X1 U861 ( .A1(n771), .A2(G8), .ZN(n772) );
  NAND2_X1 U862 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X2 U864 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U865 ( .A1(G166), .A2(G8), .ZN(n778) );
  NOR2_X1 U866 ( .A1(G2090), .A2(n778), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n520), .A2(n785), .ZN(n800) );
  INV_X1 U868 ( .A(n781), .ZN(n783) );
  NOR2_X1 U869 ( .A1(G1976), .A2(G288), .ZN(n787) );
  NOR2_X1 U870 ( .A1(G1971), .A2(G303), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n787), .A2(n782), .ZN(n1016) );
  NAND2_X1 U872 ( .A1(n783), .A2(n1016), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G288), .A2(G1976), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT105), .B(n784), .Z(n1019) );
  INV_X1 U875 ( .A(n1019), .ZN(n786) );
  AND2_X1 U876 ( .A1(n787), .A2(KEYINPUT33), .ZN(n788) );
  AND2_X1 U877 ( .A1(n788), .A2(n794), .ZN(n789) );
  XNOR2_X1 U878 ( .A(G1981), .B(G305), .ZN(n1022) );
  NOR2_X1 U879 ( .A1(n789), .A2(n1022), .ZN(n792) );
  AND2_X1 U880 ( .A1(n524), .A2(n792), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n799) );
  AND2_X1 U882 ( .A1(n792), .A2(KEYINPUT33), .ZN(n797) );
  NOR2_X1 U883 ( .A1(G1981), .A2(G305), .ZN(n793) );
  XNOR2_X1 U884 ( .A(n793), .B(KEYINPUT24), .ZN(n795) );
  AND2_X1 U885 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n800), .A2(n521), .ZN(n832) );
  NAND2_X1 U888 ( .A1(n802), .A2(n801), .ZN(n830) );
  XNOR2_X1 U889 ( .A(KEYINPUT37), .B(G2067), .ZN(n841) );
  NAND2_X1 U890 ( .A1(G140), .A2(n903), .ZN(n804) );
  NAND2_X1 U891 ( .A1(G104), .A2(n904), .ZN(n803) );
  NAND2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U893 ( .A(KEYINPUT34), .B(n805), .ZN(n810) );
  NAND2_X1 U894 ( .A1(G116), .A2(n909), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G128), .A2(n907), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U897 ( .A(n808), .B(KEYINPUT35), .Z(n809) );
  NOR2_X1 U898 ( .A1(n810), .A2(n809), .ZN(n811) );
  XOR2_X1 U899 ( .A(KEYINPUT36), .B(n811), .Z(n812) );
  XOR2_X1 U900 ( .A(KEYINPUT94), .B(n812), .Z(n918) );
  OR2_X1 U901 ( .A1(n841), .A2(n918), .ZN(n953) );
  NOR2_X1 U902 ( .A1(n830), .A2(n953), .ZN(n839) );
  INV_X1 U903 ( .A(n839), .ZN(n829) );
  NAND2_X1 U904 ( .A1(G131), .A2(n903), .ZN(n814) );
  NAND2_X1 U905 ( .A1(G95), .A2(n904), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n814), .A2(n813), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G107), .A2(n909), .ZN(n816) );
  NAND2_X1 U908 ( .A1(G119), .A2(n907), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n895) );
  INV_X1 U911 ( .A(G1991), .ZN(n985) );
  NOR2_X1 U912 ( .A1(n895), .A2(n985), .ZN(n827) );
  NAND2_X1 U913 ( .A1(G141), .A2(n903), .ZN(n820) );
  NAND2_X1 U914 ( .A1(G129), .A2(n907), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n904), .A2(G105), .ZN(n821) );
  XOR2_X1 U917 ( .A(KEYINPUT38), .B(n821), .Z(n822) );
  NOR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U919 ( .A1(n909), .A2(G117), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n915) );
  AND2_X1 U921 ( .A1(G1996), .A2(n915), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n970) );
  NOR2_X1 U923 ( .A1(n970), .A2(n830), .ZN(n835) );
  XNOR2_X1 U924 ( .A(KEYINPUT95), .B(n835), .ZN(n828) );
  XNOR2_X1 U925 ( .A(G1986), .B(G290), .ZN(n1014) );
  INV_X1 U926 ( .A(n830), .ZN(n843) );
  NAND2_X1 U927 ( .A1(n1014), .A2(n843), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n832), .A2(n522), .ZN(n846) );
  NOR2_X1 U929 ( .A1(G1996), .A2(n915), .ZN(n967) );
  AND2_X1 U930 ( .A1(n985), .A2(n895), .ZN(n963) );
  NOR2_X1 U931 ( .A1(G1986), .A2(G290), .ZN(n833) );
  NOR2_X1 U932 ( .A1(n963), .A2(n833), .ZN(n834) );
  NOR2_X1 U933 ( .A1(n835), .A2(n834), .ZN(n836) );
  NOR2_X1 U934 ( .A1(n967), .A2(n836), .ZN(n837) );
  XOR2_X1 U935 ( .A(KEYINPUT39), .B(n837), .Z(n838) );
  NOR2_X1 U936 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n840), .B(KEYINPUT107), .ZN(n842) );
  NAND2_X1 U938 ( .A1(n918), .A2(n841), .ZN(n954) );
  NAND2_X1 U939 ( .A1(n842), .A2(n954), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n844), .A2(n843), .ZN(n845) );
  NAND2_X1 U941 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n847), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U943 ( .A1(G2106), .A2(n848), .ZN(G217) );
  AND2_X1 U944 ( .A1(G15), .A2(G2), .ZN(n849) );
  NAND2_X1 U945 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U946 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U947 ( .A1(n851), .A2(n850), .ZN(G188) );
  XOR2_X1 U948 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  INV_X1 U950 ( .A(G57), .ZN(G237) );
  NOR2_X1 U951 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  XOR2_X1 U953 ( .A(KEYINPUT114), .B(n854), .Z(n856) );
  XNOR2_X1 U954 ( .A(G171), .B(G286), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  NOR2_X1 U957 ( .A1(G37), .A2(n859), .ZN(G397) );
  XNOR2_X1 U958 ( .A(G1961), .B(KEYINPUT41), .ZN(n869) );
  XOR2_X1 U959 ( .A(G1981), .B(G1971), .Z(n861) );
  XNOR2_X1 U960 ( .A(G1986), .B(G1966), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U962 ( .A(G1976), .B(G1956), .Z(n863) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(n865), .B(n864), .Z(n867) );
  XNOR2_X1 U966 ( .A(G2474), .B(KEYINPUT110), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(G229) );
  XOR2_X1 U969 ( .A(KEYINPUT109), .B(G2078), .Z(n871) );
  XNOR2_X1 U970 ( .A(G2067), .B(G2072), .ZN(n870) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U972 ( .A(n872), .B(G2096), .Z(n874) );
  XNOR2_X1 U973 ( .A(G2084), .B(G2090), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U975 ( .A(G2678), .B(KEYINPUT43), .Z(n876) );
  XNOR2_X1 U976 ( .A(KEYINPUT42), .B(G2100), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(n878), .B(n877), .Z(G227) );
  NAND2_X1 U979 ( .A1(G124), .A2(n907), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n879), .B(KEYINPUT44), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G112), .A2(n909), .ZN(n880) );
  XOR2_X1 U982 ( .A(KEYINPUT111), .B(n880), .Z(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U984 ( .A1(G136), .A2(n903), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G100), .A2(n904), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U987 ( .A1(n886), .A2(n885), .ZN(G162) );
  NAND2_X1 U988 ( .A1(G118), .A2(n909), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G130), .A2(n907), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U991 ( .A1(n904), .A2(G106), .ZN(n889) );
  XNOR2_X1 U992 ( .A(n889), .B(KEYINPUT112), .ZN(n891) );
  NAND2_X1 U993 ( .A1(G142), .A2(n903), .ZN(n890) );
  NAND2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U995 ( .A(KEYINPUT45), .B(n892), .Z(n893) );
  NOR2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n899) );
  XNOR2_X1 U997 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n897) );
  XNOR2_X1 U998 ( .A(G160), .B(n895), .ZN(n896) );
  XNOR2_X1 U999 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U1000 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U1001 ( .A(G164), .B(n962), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1003 ( .A(n902), .B(G162), .Z(n917) );
  NAND2_X1 U1004 ( .A1(G139), .A2(n903), .ZN(n906) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n904), .ZN(n905) );
  NAND2_X1 U1006 ( .A1(n906), .A2(n905), .ZN(n914) );
  NAND2_X1 U1007 ( .A1(n907), .A2(G127), .ZN(n908) );
  XOR2_X1 U1008 ( .A(KEYINPUT113), .B(n908), .Z(n911) );
  NAND2_X1 U1009 ( .A1(n909), .A2(G115), .ZN(n910) );
  NAND2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1011 ( .A(KEYINPUT47), .B(n912), .Z(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n955) );
  XOR2_X1 U1013 ( .A(n915), .B(n955), .Z(n916) );
  XNOR2_X1 U1014 ( .A(n917), .B(n916), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(n919), .B(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n920), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G397), .A2(n922), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(G401), .A2(n927), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(KEYINPUT115), .B(n923), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G395), .A2(n924), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(n927), .ZN(G319) );
  XNOR2_X1 U1026 ( .A(G1341), .B(G19), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(G6), .B(G1981), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n935) );
  XOR2_X1 U1029 ( .A(KEYINPUT126), .B(G4), .Z(n931) );
  XNOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .ZN(n930) );
  XNOR2_X1 U1031 ( .A(n931), .B(n930), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(G1956), .B(G20), .ZN(n932) );
  NOR2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n936), .B(KEYINPUT60), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(G1971), .B(G22), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(G23), .B(G1976), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n940) );
  XOR2_X1 U1039 ( .A(G1986), .B(G24), .Z(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(KEYINPUT58), .B(n941), .ZN(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G21), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(G5), .B(G1961), .ZN(n944) );
  NOR2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(n948), .B(KEYINPUT61), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(KEYINPUT127), .B(n949), .ZN(n951) );
  INV_X1 U1049 ( .A(G16), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1051 ( .A1(n952), .A2(G11), .ZN(n982) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n961) );
  XOR2_X1 U1053 ( .A(G2072), .B(n955), .Z(n957) );
  XOR2_X1 U1054 ( .A(G164), .B(G2078), .Z(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1056 ( .A(KEYINPUT116), .B(n958), .Z(n959) );
  XNOR2_X1 U1057 ( .A(KEYINPUT50), .B(n959), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n974) );
  XNOR2_X1 U1059 ( .A(G2084), .B(G160), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n972) );
  XOR2_X1 U1062 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1064 ( .A(KEYINPUT51), .B(n968), .Z(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(KEYINPUT52), .B(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n976) );
  XNOR2_X1 U1070 ( .A(n977), .B(n976), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(KEYINPUT55), .A2(n978), .ZN(n980) );
  INV_X1 U1072 ( .A(G29), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n1008) );
  XNOR2_X1 U1075 ( .A(KEYINPUT54), .B(G34), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT121), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G2084), .B(n984), .ZN(n1002) );
  XNOR2_X1 U1078 ( .A(G2090), .B(G35), .ZN(n1000) );
  XNOR2_X1 U1079 ( .A(G25), .B(n985), .ZN(n986) );
  NAND2_X1 U1080 ( .A1(n986), .A2(G28), .ZN(n997) );
  XOR2_X1 U1081 ( .A(G2067), .B(G26), .Z(n987) );
  XNOR2_X1 U1082 ( .A(KEYINPUT119), .B(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(G33), .B(G2072), .ZN(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(KEYINPUT120), .B(n990), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(G1996), .B(G32), .ZN(n993) );
  XNOR2_X1 U1087 ( .A(n991), .B(G27), .ZN(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT53), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(n1003), .B(KEYINPUT122), .ZN(n1004) );
  XOR2_X1 U1095 ( .A(KEYINPUT55), .B(n1004), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(G29), .B(KEYINPUT123), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1035) );
  XOR2_X1 U1099 ( .A(G16), .B(KEYINPUT56), .Z(n1033) );
  XOR2_X1 U1100 ( .A(n1009), .B(G1341), .Z(n1011) );
  XNOR2_X1 U1101 ( .A(G171), .B(G1961), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1031) );
  XNOR2_X1 U1103 ( .A(G1348), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1029) );
  NAND2_X1 U1105 ( .A1(G1971), .A2(G303), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(G1956), .B(G299), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XOR2_X1 U1110 ( .A(G168), .B(G1966), .Z(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(KEYINPUT125), .B(n1023), .Z(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(n1025), .B(n1024), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1036), .ZN(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

