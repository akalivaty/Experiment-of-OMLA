//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G87), .A2(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G58), .ZN(new_n206));
  INV_X1    g0006(.A(G232), .ZN(new_n207));
  OAI21_X1  g0007(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AND2_X1   g0008(.A1(G107), .A2(G264), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G77), .A2(G244), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(KEYINPUT66), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n208), .B(new_n209), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G97), .A2(G257), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n216), .B(new_n217), .C1(new_n215), .C2(new_n214), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT1), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(KEYINPUT65), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT65), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n224), .A2(G1), .A3(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OR3_X1    g0031(.A1(new_n219), .A2(KEYINPUT64), .A3(G13), .ZN(new_n232));
  OAI21_X1  g0032(.A(KEYINPUT64), .B1(new_n219), .B2(G13), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n234), .B(G250), .C1(G257), .C2(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT0), .ZN(new_n236));
  NAND3_X1  g0036(.A1(new_n221), .A2(new_n231), .A3(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n213), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT67), .Z(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n207), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT2), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n245), .B(G226), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n242), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n206), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT68), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n252), .B(new_n255), .Z(G351));
  AND3_X1   g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n226), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT7), .B1(new_n262), .B2(new_n227), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(G68), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G159), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G58), .A2(G68), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n227), .B1(new_n202), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n270), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  AND3_X1   g0079(.A1(new_n279), .A2(KEYINPUT80), .A3(KEYINPUT16), .ZN(new_n280));
  AOI21_X1  g0080(.A(KEYINPUT16), .B1(new_n279), .B2(KEYINPUT80), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n259), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n257), .B1(new_n223), .B2(new_n225), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G1), .B2(new_n227), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n285), .ZN(new_n288));
  INV_X1    g0088(.A(G13), .ZN(new_n289));
  NOR3_X1   g0089(.A1(new_n289), .A2(new_n227), .A3(G1), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n282), .A2(new_n287), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n266), .A2(new_n267), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G226), .A3(G1698), .ZN(new_n296));
  INV_X1    g0096(.A(G1698), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(G223), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G87), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n296), .B(new_n298), .C1(new_n265), .C2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G1), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G41), .B2(G45), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT69), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  OAI211_X1 g0106(.A(G1), .B(G13), .C1(new_n265), .C2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(G274), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n304), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G232), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n302), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n311), .A2(G179), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n294), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT18), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n313), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT16), .ZN(new_n319));
  INV_X1    g0119(.A(G68), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n266), .A2(new_n227), .A3(new_n267), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT7), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n323), .B2(new_n268), .ZN(new_n324));
  NOR3_X1   g0124(.A1(new_n324), .A2(new_n274), .A3(new_n277), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT80), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n279), .A2(KEYINPUT80), .A3(KEYINPUT16), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n286), .B1(new_n329), .B2(new_n259), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n318), .B1(new_n330), .B2(new_n293), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT18), .A3(new_n314), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n311), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n311), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n330), .A2(new_n293), .A3(new_n333), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT17), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n283), .B1(new_n327), .B2(new_n328), .ZN(new_n339));
  NOR4_X1   g0139(.A1(new_n339), .A2(new_n286), .A3(new_n335), .A4(new_n292), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT17), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n333), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n317), .A2(new_n332), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n295), .A2(G238), .A3(G1698), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n295), .A2(G232), .A3(new_n297), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n262), .A2(G107), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT71), .A4(new_n346), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n301), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n309), .A2(G244), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n308), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n312), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n288), .A2(new_n271), .B1(G20), .B2(G77), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n227), .A2(G33), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT15), .B(G87), .Z(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n355), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n259), .ZN(new_n360));
  INV_X1    g0160(.A(G77), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n290), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT72), .ZN(new_n363));
  INV_X1    g0163(.A(new_n284), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT73), .B1(new_n364), .B2(G77), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT73), .ZN(new_n366));
  NOR3_X1   g0166(.A1(new_n284), .A2(new_n366), .A3(new_n361), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n360), .B(new_n363), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G179), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n351), .A2(new_n369), .A3(new_n308), .A4(new_n352), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n354), .B(new_n368), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n368), .B1(G200), .B2(new_n353), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n334), .B2(new_n353), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(G223), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n379));
  OAI211_X1 g0179(.A(G222), .B(new_n297), .C1(new_n260), .C2(new_n261), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n266), .A2(G77), .A3(new_n267), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT70), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n379), .A2(new_n380), .A3(KEYINPUT70), .A4(new_n381), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(new_n301), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n309), .A2(G226), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n308), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n388), .A2(new_n312), .ZN(new_n389));
  INV_X1    g0189(.A(G150), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n285), .A2(new_n356), .B1(new_n390), .B2(new_n272), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n227), .B1(new_n201), .B2(new_n251), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n259), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n290), .A2(new_n251), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(new_n251), .C2(new_n284), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n388), .B2(G179), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n343), .A2(new_n378), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n290), .A2(new_n320), .ZN(new_n399));
  NAND2_X1  g0199(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n400));
  OR2_X1    g0200(.A1(KEYINPUT78), .A2(KEYINPUT12), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n402), .B(KEYINPUT79), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(KEYINPUT12), .B2(new_n399), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n364), .A2(G68), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n272), .A2(new_n251), .B1(new_n356), .B2(new_n361), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n227), .A2(G68), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n259), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g0208(.A(new_n408), .B(KEYINPUT11), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n295), .A2(G226), .A3(new_n297), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n295), .A2(G232), .A3(G1698), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n301), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n309), .A2(G238), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n416), .A2(new_n308), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n415), .A2(new_n301), .B1(G238), .B2(new_n309), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n308), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G200), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT77), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT76), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(new_n426), .A3(new_n422), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n421), .B1(new_n420), .B2(new_n308), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n425), .B1(new_n430), .B2(G190), .ZN(new_n431));
  AOI211_X1 g0231(.A(KEYINPUT77), .B(new_n334), .C1(new_n427), .C2(new_n429), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n411), .B(new_n424), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n423), .A2(G169), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n423), .A2(new_n436), .A3(G169), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n369), .B1(new_n427), .B2(new_n429), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n410), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n388), .A2(G200), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT9), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n395), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n386), .A2(G190), .A3(new_n308), .A4(new_n387), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n395), .A2(new_n442), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n441), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT10), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n388), .A2(G200), .B1(new_n442), .B2(new_n395), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT10), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n443), .A4(new_n444), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n433), .A2(new_n440), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n377), .B1(new_n374), .B2(new_n376), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n398), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  OR2_X1    g0255(.A1(KEYINPUT81), .A2(G97), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT81), .A2(G97), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n227), .B(new_n455), .C1(new_n458), .C2(G33), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n227), .A2(G116), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT85), .B1(new_n259), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT85), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n283), .A2(new_n463), .A3(new_n460), .ZN(new_n464));
  OAI211_X1 g0264(.A(KEYINPUT20), .B(new_n459), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT86), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n459), .B1(new_n462), .B2(new_n464), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT20), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n259), .A2(KEYINPUT85), .A3(new_n461), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n463), .B1(new_n283), .B2(new_n460), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(KEYINPUT86), .A3(KEYINPUT20), .A4(new_n459), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n467), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n291), .A2(G116), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n303), .A2(G33), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n283), .A2(new_n291), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(G116), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT5), .B(G41), .ZN(new_n482));
  INV_X1    g0282(.A(G45), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G1), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n482), .A2(new_n307), .A3(G274), .A4(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n487));
  OAI211_X1 g0287(.A(G257), .B(new_n297), .C1(new_n260), .C2(new_n261), .ZN(new_n488));
  INV_X1    g0288(.A(G303), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n487), .B(new_n488), .C1(new_n489), .C2(new_n295), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n490), .B2(new_n301), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n484), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(G270), .A3(new_n307), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n494), .A2(KEYINPUT84), .A3(G270), .A4(new_n307), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n312), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n481), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n481), .A2(KEYINPUT21), .A3(new_n500), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n491), .A2(new_n499), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n369), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n481), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n505), .A2(new_n334), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(G200), .B2(new_n505), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(new_n475), .A3(new_n480), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n503), .A2(new_n504), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(G20), .B1(new_n266), .B2(new_n267), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT22), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n299), .B1(G33), .B2(G116), .ZN(new_n516));
  OR2_X1    g0316(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n513), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(KEYINPUT88), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G116), .ZN(new_n520));
  AOI21_X1  g0320(.A(G20), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n518), .B1(new_n521), .B2(new_n515), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n227), .A2(G107), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT23), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n523), .B1(new_n522), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n259), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n479), .A2(G107), .ZN(new_n529));
  INV_X1    g0329(.A(G107), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n290), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g0331(.A(new_n531), .B(KEYINPUT25), .Z(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G257), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n534));
  OAI211_X1 g0334(.A(G250), .B(new_n297), .C1(new_n260), .C2(new_n261), .ZN(new_n535));
  INV_X1    g0335(.A(G294), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n535), .C1(new_n265), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n301), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n494), .A2(G264), .A3(new_n307), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n538), .A2(new_n485), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n312), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n538), .A2(new_n539), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n369), .A3(new_n485), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n533), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n295), .A2(G244), .A3(G1698), .ZN(new_n545));
  OAI211_X1 g0345(.A(G238), .B(new_n297), .C1(new_n260), .C2(new_n261), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n520), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n301), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n484), .A2(G274), .ZN(new_n549));
  INV_X1    g0349(.A(new_n484), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n307), .A2(new_n550), .A3(G250), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G200), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n548), .A2(G190), .A3(new_n549), .A4(new_n551), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n291), .A2(new_n357), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n458), .A2(new_n299), .A3(new_n530), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n227), .B1(new_n414), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n513), .A2(G68), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n458), .B2(new_n356), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n555), .B1(new_n562), .B2(new_n259), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n478), .A2(new_n299), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n553), .A2(new_n554), .A3(new_n563), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n259), .ZN(new_n567));
  INV_X1    g0367(.A(new_n555), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n479), .A2(new_n357), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n552), .A2(new_n312), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n548), .A2(new_n369), .A3(new_n549), .A4(new_n551), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(G200), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n540), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n538), .A2(new_n539), .A3(new_n334), .A4(new_n485), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n528), .A2(new_n529), .A3(new_n578), .A4(new_n532), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n544), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n291), .A2(G97), .ZN(new_n581));
  INV_X1    g0381(.A(G97), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n478), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(G107), .B1(new_n263), .B2(new_n269), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n456), .A2(KEYINPUT6), .A3(new_n530), .A4(new_n457), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT6), .ZN(new_n586));
  AND2_X1   g0386(.A1(G97), .A2(G107), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n227), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n272), .A2(new_n361), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n584), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI211_X1 g0394(.A(new_n581), .B(new_n583), .C1(new_n594), .C2(new_n259), .ZN(new_n595));
  OAI211_X1 g0395(.A(G244), .B(new_n297), .C1(new_n260), .C2(new_n261), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT4), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n295), .A2(KEYINPUT4), .A3(G244), .A4(new_n297), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n295), .A2(G250), .A3(G1698), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n455), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n301), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n494), .A2(G257), .A3(new_n307), .ZN(new_n603));
  AOI21_X1  g0403(.A(KEYINPUT82), .B1(new_n603), .B2(new_n485), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n485), .A3(KEYINPUT82), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n602), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G200), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n603), .A2(new_n485), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT82), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n605), .B1(new_n601), .B2(new_n301), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G190), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n595), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n581), .B1(new_n594), .B2(new_n259), .ZN(new_n617));
  INV_X1    g0417(.A(new_n583), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n617), .A2(new_n618), .B1(new_n612), .B2(new_n369), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n607), .A2(new_n312), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n595), .A2(new_n608), .A3(new_n613), .A4(KEYINPUT83), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n616), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n580), .A2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n454), .A2(new_n512), .A3(new_n624), .ZN(G372));
  INV_X1    g0425(.A(new_n397), .ZN(new_n626));
  INV_X1    g0426(.A(new_n433), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n440), .B1(new_n627), .B2(new_n374), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n338), .A2(new_n342), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT18), .B1(new_n331), .B2(new_n314), .ZN(new_n631));
  AND4_X1   g0431(.A1(KEYINPUT18), .A2(new_n294), .A3(new_n313), .A4(new_n314), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n447), .A2(KEYINPUT91), .A3(new_n450), .ZN(new_n634));
  AOI21_X1  g0434(.A(KEYINPUT91), .B1(new_n447), .B2(new_n450), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n626), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT89), .ZN(new_n639));
  INV_X1    g0439(.A(new_n549), .ZN(new_n640));
  INV_X1    g0440(.A(new_n551), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n640), .B(new_n641), .C1(new_n547), .C2(new_n301), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n639), .B1(new_n642), .B2(new_n575), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n555), .B(new_n564), .C1(new_n259), .C2(new_n562), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n552), .A2(KEYINPUT89), .A3(G200), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n554), .A4(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n573), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n638), .B1(new_n647), .B2(new_n621), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n619), .A2(new_n566), .A3(new_n573), .A4(new_n620), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT90), .B1(new_n649), .B2(new_n638), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n612), .A2(new_n369), .ZN(new_n652));
  INV_X1    g0452(.A(new_n581), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n530), .B1(new_n323), .B2(new_n268), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n654), .A2(new_n590), .A3(new_n592), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n653), .B(new_n618), .C1(new_n655), .C2(new_n283), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n620), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n574), .A2(new_n651), .A3(KEYINPUT26), .A4(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n648), .A2(new_n650), .A3(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n503), .A2(new_n504), .A3(new_n507), .A4(new_n544), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n611), .A2(new_n605), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n575), .B1(new_n661), .B2(new_n602), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n656), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT83), .B1(new_n663), .B2(new_n613), .ZN(new_n664));
  AND4_X1   g0464(.A1(KEYINPUT83), .A2(new_n595), .A3(new_n608), .A4(new_n613), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n579), .A2(new_n573), .A3(new_n646), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(new_n667), .A3(new_n621), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n573), .B(new_n659), .C1(new_n660), .C2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n454), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n637), .A2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(G330), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n289), .A2(G20), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n303), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n481), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n512), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n481), .A3(new_n679), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n672), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n533), .A2(new_n679), .ZN(new_n689));
  INV_X1    g0489(.A(new_n579), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n544), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n544), .A2(new_n679), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT93), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT93), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n688), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n679), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n682), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n694), .B2(new_n696), .ZN(new_n701));
  INV_X1    g0501(.A(new_n692), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n234), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n458), .A2(new_n299), .A3(new_n530), .A4(new_n212), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n229), .B2(new_n707), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  INV_X1    g0512(.A(new_n573), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n579), .A2(new_n573), .A3(new_n646), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n623), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n503), .A2(new_n504), .A3(new_n507), .A4(new_n544), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n679), .B1(new_n717), .B2(new_n659), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n647), .A2(new_n638), .A3(new_n621), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n649), .A2(new_n638), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n717), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n721), .B1(new_n726), .B2(new_n699), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n512), .A2(new_n624), .A3(new_n699), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n506), .A2(new_n612), .A3(new_n642), .A4(new_n542), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n607), .A2(new_n505), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(new_n369), .A3(new_n552), .A4(new_n540), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n505), .A2(new_n552), .A3(new_n369), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(KEYINPUT30), .A3(new_n612), .A4(new_n542), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n731), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT31), .B1(new_n736), .B2(new_n679), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n672), .B1(new_n728), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n720), .A2(new_n727), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n712), .B1(new_n742), .B2(G1), .ZN(G364));
  NOR2_X1   g0543(.A1(new_n705), .A2(new_n295), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n230), .A2(new_n483), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n744), .B(new_n745), .C1(new_n252), .C2(new_n483), .ZN(new_n746));
  INV_X1    g0546(.A(G355), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n234), .A2(new_n295), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT96), .Z(new_n749));
  OAI221_X1 g0549(.A(new_n746), .B1(G116), .B2(new_n234), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n226), .B1(G20), .B2(new_n312), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g0556(.A1(new_n289), .A2(new_n483), .A3(G20), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT95), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(G1), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n706), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n751), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n227), .A2(new_n575), .A3(G179), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G190), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n334), .A2(G179), .A3(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n227), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n489), .B1(new_n766), .B2(new_n536), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n227), .A2(new_n369), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(G190), .A3(new_n575), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n295), .B1(new_n770), .B2(G322), .ZN(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n227), .A2(G190), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(G179), .A3(new_n575), .ZN(new_n774));
  INV_X1    g0574(.A(G329), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n773), .A2(new_n369), .A3(new_n575), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n771), .B1(new_n772), .B2(new_n774), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n768), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n767), .B(new_n777), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n763), .A2(new_n334), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT97), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT97), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n778), .A2(new_n334), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT99), .B(G326), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n781), .B1(new_n782), .B2(new_n786), .C1(new_n788), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n786), .ZN(new_n792));
  INV_X1    g0592(.A(new_n766), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G97), .ZN(new_n794));
  INV_X1    g0594(.A(new_n779), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n794), .B1(new_n795), .B2(new_n320), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n792), .A2(G107), .B1(new_n796), .B2(KEYINPUT98), .ZN(new_n797));
  OR3_X1    g0597(.A1(new_n776), .A2(KEYINPUT32), .A3(new_n273), .ZN(new_n798));
  OAI21_X1  g0598(.A(KEYINPUT32), .B1(new_n776), .B2(new_n273), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(new_n788), .C2(new_n251), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n764), .A2(new_n299), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n295), .B1(new_n774), .B2(new_n361), .C1(new_n769), .C2(new_n206), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n797), .B(new_n803), .C1(KEYINPUT98), .C2(new_n796), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n756), .B(new_n761), .C1(new_n762), .C2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT100), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(KEYINPUT100), .ZN(new_n808));
  INV_X1    g0608(.A(new_n754), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n807), .B(new_n808), .C1(new_n684), .C2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n688), .ZN(new_n811));
  INV_X1    g0611(.A(new_n761), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n685), .A2(new_n672), .A3(new_n687), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT101), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(G396));
  NAND2_X1  g0617(.A1(new_n792), .A2(G87), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n772), .B2(new_n776), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT102), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n262), .B1(new_n774), .B2(new_n212), .C1(new_n769), .C2(new_n536), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n794), .B1(new_n530), .B2(new_n764), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(G303), .C2(new_n787), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(new_n782), .C2(new_n795), .ZN(new_n824));
  INV_X1    g0624(.A(new_n774), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n787), .A2(G137), .B1(new_n825), .B2(G159), .ZN(new_n826));
  INV_X1    g0626(.A(G143), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n826), .B1(new_n827), .B2(new_n769), .C1(new_n390), .C2(new_n795), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT34), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n776), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G132), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n828), .A2(new_n829), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n295), .B1(new_n766), .B2(new_n206), .C1(new_n251), .C2(new_n764), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n792), .B2(G68), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n830), .A2(new_n832), .A3(new_n833), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n762), .B1(new_n824), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n751), .A2(new_n752), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n361), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n374), .A2(new_n679), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n368), .A2(new_n679), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n376), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n840), .B1(new_n374), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n839), .B(new_n761), .C1(new_n753), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n843), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n719), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n669), .A2(new_n699), .A3(new_n843), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n741), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g0651(.A1(new_n851), .A2(KEYINPUT104), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n761), .B1(new_n851), .B2(KEYINPUT104), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT103), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n849), .B2(new_n850), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  NOR3_X1   g0656(.A1(new_n849), .A2(new_n854), .A3(new_n850), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n844), .B1(new_n856), .B2(new_n857), .ZN(G384));
  NAND2_X1  g0658(.A1(new_n585), .A2(new_n589), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n212), .B1(new_n859), .B2(KEYINPUT35), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n860), .B(new_n228), .C1(KEYINPUT35), .C2(new_n859), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT36), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n276), .A2(G77), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n229), .A2(new_n863), .B1(G50), .B2(new_n320), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(G1), .A3(new_n289), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT105), .Z(new_n867));
  INV_X1    g0667(.A(KEYINPUT108), .ZN(new_n868));
  NOR4_X1   g0668(.A1(new_n511), .A2(new_n580), .A3(new_n623), .A4(new_n679), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n736), .A2(new_n679), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT31), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n737), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n869), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n410), .A2(new_n679), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n875), .B1(new_n433), .B2(new_n440), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n433), .A2(new_n440), .A3(new_n875), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n728), .A2(new_n740), .A3(KEYINPUT108), .ZN(new_n880));
  AND4_X1   g0680(.A1(new_n843), .A2(new_n874), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n341), .B1(new_n340), .B2(new_n333), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n282), .A2(new_n287), .A3(new_n336), .A4(new_n293), .ZN(new_n883));
  INV_X1    g0683(.A(new_n333), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n883), .A2(KEYINPUT17), .A3(new_n884), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n631), .A2(new_n632), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n677), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n294), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n315), .A2(new_n337), .A3(new_n888), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT106), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n294), .A2(new_n893), .A3(new_n887), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n294), .B2(new_n887), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n315), .B(new_n337), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n892), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n890), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n881), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n888), .A2(KEYINPUT106), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n294), .A2(new_n893), .A3(new_n887), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n315), .A2(new_n337), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI22_X1  g0712(.A1(new_n906), .A2(new_n912), .B1(new_n343), .B2(new_n910), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n899), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n905), .B1(new_n914), .B2(new_n901), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n903), .A2(new_n904), .B1(new_n915), .B2(new_n881), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n874), .A2(new_n880), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n454), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G330), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n914), .A2(new_n921), .A3(new_n901), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n890), .A2(new_n897), .A3(KEYINPUT38), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n890), .B2(new_n897), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT39), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n440), .A2(new_n679), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n332), .A2(new_n317), .A3(new_n677), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n433), .A2(new_n440), .A3(new_n875), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n931), .A2(new_n876), .ZN(new_n932));
  INV_X1    g0732(.A(new_n840), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n932), .B1(new_n847), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n902), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n454), .B1(new_n720), .B2(new_n727), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n637), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n920), .B(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n673), .A2(new_n303), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n867), .B1(new_n940), .B2(new_n941), .ZN(G367));
  OAI211_X1 g0742(.A(new_n666), .B(new_n621), .C1(new_n595), .C2(new_n699), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n657), .A2(new_n679), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n701), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT42), .Z(new_n947));
  XOR2_X1   g0747(.A(new_n945), .B(KEYINPUT109), .Z(new_n948));
  OAI21_X1  g0748(.A(new_n621), .B1(new_n948), .B2(new_n544), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n699), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n644), .A2(new_n699), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n713), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n647), .B2(new_n952), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n698), .A2(new_n948), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n960), .B1(new_n961), .B2(new_n959), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n706), .B(KEYINPUT41), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n688), .B(KEYINPUT111), .Z(new_n967));
  XNOR2_X1  g0767(.A(new_n697), .B(new_n700), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n811), .B2(KEYINPUT111), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n970), .A2(new_n742), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n703), .A2(new_n945), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT45), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n945), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n701), .B2(new_n702), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT44), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n698), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n971), .B1(new_n967), .B2(new_n969), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT112), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n986), .A2(new_n987), .A3(new_n742), .ZN(new_n988));
  INV_X1    g0788(.A(new_n698), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n982), .A2(new_n983), .A3(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n974), .A2(new_n985), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n966), .B1(new_n991), .B2(new_n742), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n964), .B1(new_n992), .B2(new_n760), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G294), .A2(new_n779), .B1(new_n787), .B2(G311), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n786), .B2(new_n458), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n262), .B1(new_n769), .B2(new_n489), .ZN(new_n996));
  INV_X1    g0796(.A(new_n764), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT46), .B1(new_n997), .B2(G116), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(G317), .C2(new_n831), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n782), .C2(new_n774), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n995), .B(new_n1001), .C1(G107), .C2(new_n793), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n792), .A2(G77), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n206), .B2(new_n764), .C1(new_n827), .C2(new_n788), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n779), .A2(G159), .B1(new_n825), .B2(G50), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT113), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n766), .A2(new_n320), .ZN(new_n1007));
  INV_X1    g0807(.A(G137), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n295), .B1(new_n776), .B2(new_n1008), .C1(new_n769), .C2(new_n390), .ZN(new_n1009));
  NOR4_X1   g0809(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT115), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1011), .B(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n812), .B1(new_n1014), .B2(new_n751), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n744), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n755), .B1(new_n234), .B2(new_n358), .C1(new_n241), .C2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(new_n809), .C2(new_n954), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n993), .A2(new_n1018), .ZN(G387));
  OR2_X1    g0819(.A1(new_n986), .A2(new_n742), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n986), .A2(new_n987), .A3(new_n742), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n987), .B1(new_n986), .B2(new_n742), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1020), .B(new_n706), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n787), .A2(G322), .B1(new_n825), .B2(G303), .ZN(new_n1024));
  INV_X1    g0824(.A(G317), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1024), .B1(new_n772), .B2(new_n795), .C1(new_n1025), .C2(new_n769), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT48), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n782), .B2(new_n766), .C1(new_n536), .C2(new_n764), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT49), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n295), .B1(new_n792), .B2(G116), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1029), .B(new_n1030), .C1(new_n776), .C2(new_n790), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n774), .A2(new_n320), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n262), .B1(new_n770), .B2(G50), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n788), .A2(new_n273), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT116), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1033), .B1(new_n390), .B2(new_n776), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1035), .B2(new_n1034), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n357), .A2(new_n793), .B1(new_n779), .B2(new_n288), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n792), .A2(G97), .B1(G77), .B2(new_n997), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1031), .B1(new_n1032), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n285), .A2(G50), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT50), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(G68), .A2(G77), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1043), .A2(new_n483), .A3(new_n1044), .A4(new_n709), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n744), .B(new_n1045), .C1(new_n246), .C2(new_n483), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(G107), .B2(new_n234), .C1(new_n709), .C2(new_n749), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1041), .A2(new_n751), .B1(new_n755), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n761), .C1(new_n697), .C2(new_n809), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n986), .B2(new_n760), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1023), .A2(new_n1051), .ZN(G393));
  XNOR2_X1  g0852(.A(new_n982), .B(new_n989), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n991), .A3(new_n706), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n760), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n948), .A2(new_n754), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n788), .A2(new_n1025), .B1(new_n772), .B2(new_n769), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n792), .A2(G107), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n779), .A2(G303), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n262), .B1(new_n774), .B2(new_n536), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n764), .A2(new_n782), .B1(new_n766), .B2(new_n212), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1063), .B(new_n1064), .C1(G322), .C2(new_n831), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n766), .A2(new_n361), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n295), .B1(new_n776), .B2(new_n827), .C1(new_n285), .C2(new_n774), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(G68), .C2(new_n997), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n818), .C1(new_n251), .C2(new_n795), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G150), .A2(new_n787), .B1(new_n770), .B2(G159), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT51), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1066), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n812), .B1(new_n1073), .B2(new_n751), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n744), .A2(new_n255), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n755), .C1(new_n234), .C2(new_n458), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT117), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1058), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1055), .A2(new_n1057), .A3(new_n1078), .ZN(G390));
  NAND3_X1  g0879(.A1(new_n917), .A2(G330), .A3(new_n454), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n937), .A2(new_n1080), .A3(new_n637), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n840), .B1(new_n718), .B2(new_n843), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n850), .A2(new_n845), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1084), .A2(new_n879), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n874), .A2(new_n879), .A3(new_n880), .A4(new_n843), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n672), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1084), .A2(new_n879), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n874), .A2(new_n880), .A3(G330), .A4(new_n843), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n932), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n726), .A2(new_n699), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n842), .A2(new_n374), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n840), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1089), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1081), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(KEYINPUT118), .B1(new_n934), .B2(new_n928), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT118), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1099), .B(new_n927), .C1(new_n1082), .C2(new_n932), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1098), .A2(new_n1100), .A3(new_n925), .A4(new_n922), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n910), .A2(new_n911), .A3(new_n907), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n910), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1102), .A2(new_n1103), .B1(new_n886), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n901), .B1(new_n1105), .B2(KEYINPUT38), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n927), .B(new_n1106), .C1(new_n1094), .C2(new_n932), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1101), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1087), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1089), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1101), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1097), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1101), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1087), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1096), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1113), .A2(new_n1116), .A3(new_n706), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n760), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n262), .B1(new_n774), .B2(new_n458), .C1(new_n769), .C2(new_n212), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n801), .A2(new_n1067), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(new_n530), .B2(new_n795), .ZN(new_n1122));
  AOI211_X1 g0922(.A(new_n1120), .B(new_n1122), .C1(G294), .C2(new_n831), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1123), .B1(new_n320), .B2(new_n786), .C1(new_n782), .C2(new_n788), .ZN(new_n1124));
  INV_X1    g0924(.A(G125), .ZN(new_n1125));
  XOR2_X1   g0925(.A(KEYINPUT54), .B(G143), .Z(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n295), .B1(new_n1125), .B2(new_n776), .C1(new_n1127), .C2(new_n774), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n795), .A2(new_n1008), .B1(new_n273), .B2(new_n766), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(G132), .C2(new_n770), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1130), .B1(new_n251), .B2(new_n786), .C1(new_n1131), .C2(new_n788), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n997), .A2(G150), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT53), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1124), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1135), .A2(new_n751), .B1(new_n285), .B2(new_n838), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n761), .B(new_n1136), .C1(new_n926), .C2(new_n753), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1117), .A2(new_n1119), .A3(new_n1137), .ZN(G378));
  INV_X1    g0938(.A(KEYINPUT56), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT91), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n451), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n447), .A2(KEYINPUT91), .A3(new_n450), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n397), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n395), .A2(new_n887), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT55), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1141), .A2(new_n397), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1147), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1139), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1144), .B1(new_n636), .B2(new_n397), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1148), .ZN(new_n1153));
  OAI21_X1  g0953(.A(KEYINPUT55), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(KEYINPUT56), .A3(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1151), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT120), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n752), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n838), .A2(new_n251), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n788), .A2(new_n1125), .B1(new_n764), .B2(new_n1127), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n779), .A2(G132), .B1(new_n825), .B2(G137), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1131), .B2(new_n769), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(G150), .C2(new_n793), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT59), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G41), .B1(new_n792), .B2(G159), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G33), .B1(new_n831), .B2(G124), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n795), .A2(new_n582), .B1(new_n320), .B2(new_n766), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G107), .A2(new_n770), .B1(new_n831), .B2(G283), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n358), .B2(new_n774), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G116), .C2(new_n787), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n792), .A2(G58), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n306), .B(new_n262), .C1(new_n764), .C2(new_n361), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT119), .Z(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT58), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n251), .B1(new_n260), .B2(G41), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1169), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n812), .B1(new_n1180), .B2(new_n751), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1160), .A2(new_n1161), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n929), .A2(new_n930), .A3(new_n935), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1149), .A2(new_n1150), .A3(new_n1139), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT56), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n916), .B2(G330), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n923), .A2(new_n924), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n904), .B1(new_n1189), .B2(new_n1086), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n874), .A2(new_n843), .A3(new_n880), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1191), .A2(new_n1106), .A3(KEYINPUT40), .A4(new_n879), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(G330), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT120), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1151), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1193), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1184), .B1(new_n1188), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n916), .A2(new_n1159), .A3(G330), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1187), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1193), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n936), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1183), .B1(new_n1204), .B2(new_n760), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1081), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1116), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n707), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1116), .B2(new_n1207), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT121), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1199), .A2(new_n1213), .A3(new_n1203), .ZN(new_n1214));
  OAI211_X1 g1014(.A(KEYINPUT121), .B(new_n1184), .C1(new_n1188), .C2(new_n1198), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1206), .B1(new_n1211), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(G375));
  NAND2_X1  g1018(.A1(new_n932), .A2(new_n752), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n262), .B1(new_n774), .B2(new_n530), .C1(new_n769), .C2(new_n782), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G303), .B2(new_n831), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n357), .A2(new_n793), .B1(new_n779), .B2(G116), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n787), .A2(G294), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1003), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n764), .A2(new_n582), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n779), .A2(new_n1126), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n295), .B1(new_n769), .B2(new_n1008), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G150), .B2(new_n825), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G50), .A2(new_n793), .B1(new_n787), .B2(G132), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1174), .A2(new_n1226), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n764), .A2(new_n273), .B1(new_n776), .B2(new_n1131), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT122), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1224), .A2(new_n1225), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1233), .A2(new_n751), .B1(new_n320), .B2(new_n838), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1219), .A2(new_n761), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1088), .A2(new_n1095), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(new_n760), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1088), .A2(new_n1081), .A3(new_n1095), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n965), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1239), .B2(new_n1096), .ZN(G381));
  XNOR2_X1  g1040(.A(new_n1217), .B(KEYINPUT123), .ZN(new_n1241));
  INV_X1    g1041(.A(G378), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G384), .A2(G381), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT124), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1023), .A2(new_n816), .A3(new_n1051), .ZN(new_n1246));
  OR3_X1    g1046(.A1(G387), .A2(G390), .A3(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1245), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(G407));
  NAND3_X1  g1050(.A1(new_n1241), .A2(new_n678), .A3(new_n1242), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(G407), .A2(G213), .A3(new_n1251), .ZN(G409));
  NAND2_X1  g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1246), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1253), .A2(KEYINPUT126), .A3(new_n1246), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1256), .A2(KEYINPUT127), .A3(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n993), .A2(new_n1018), .A3(G390), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1257), .B2(new_n1256), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G390), .B1(new_n993), .B2(new_n1018), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1261), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1263), .A2(KEYINPUT127), .A3(new_n1264), .A4(new_n1259), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n678), .A2(G213), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1199), .A2(new_n1203), .B1(new_n1116), .B2(new_n1207), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n706), .B1(new_n1269), .B2(KEYINPUT57), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1271));
  OAI211_X1 g1071(.A(G378), .B(new_n1205), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1200), .A2(new_n936), .A3(new_n1202), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n936), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1081), .B1(new_n1118), .B2(new_n1236), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1210), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1216), .A3(new_n706), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1280), .A2(KEYINPUT125), .A3(G378), .A4(new_n1205), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1274), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1214), .A2(new_n760), .A3(new_n1215), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1182), .C1(new_n966), .C2(new_n1209), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1284), .A2(new_n1242), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1268), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n707), .B1(new_n1238), .B2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1288), .B(new_n1097), .C1(new_n1287), .C2(new_n1238), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(G384), .A3(new_n1237), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G384), .B1(new_n1289), .B2(new_n1237), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1286), .A2(KEYINPUT63), .A3(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT63), .ZN(new_n1295));
  AOI21_X1  g1095(.A(KEYINPUT125), .B1(new_n1217), .B2(G378), .ZN(new_n1296));
  AND4_X1   g1096(.A1(KEYINPUT125), .A2(new_n1280), .A3(G378), .A4(new_n1205), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1285), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1267), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1293), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(G2897), .A3(new_n1268), .ZN(new_n1301));
  INV_X1    g1101(.A(G2897), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1293), .B1(new_n1302), .B2(new_n1267), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1295), .B1(new_n1299), .B2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1266), .B(new_n1294), .C1(new_n1306), .C2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1286), .B2(new_n1304), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1286), .B2(new_n1293), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1274), .A2(new_n1281), .B1(new_n1242), .B2(new_n1284), .ZN(new_n1313));
  NOR4_X1   g1113(.A1(new_n1313), .A2(KEYINPUT62), .A3(new_n1268), .A4(new_n1300), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1310), .A2(new_n1312), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1262), .A2(new_n1265), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1308), .B1(new_n1315), .B2(new_n1316), .ZN(G405));
  OAI21_X1  g1117(.A(new_n1282), .B1(G378), .B2(new_n1217), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1293), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1318), .A2(new_n1293), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1320), .A2(new_n1316), .A3(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1321), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1323), .A2(new_n1319), .B1(new_n1262), .B2(new_n1265), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1322), .A2(new_n1324), .ZN(G402));
endmodule


