//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT64), .B1(new_n196), .B2(new_n192), .ZN(new_n197));
  AND4_X1   g011(.A1(KEYINPUT64), .A2(new_n188), .A3(new_n190), .A4(new_n192), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI211_X1 g015(.A(KEYINPUT68), .B(new_n195), .C1(new_n197), .C2(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT66), .B(G137), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  AOI21_X1  g020(.A(KEYINPUT11), .B1(new_n206), .B2(G134), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G137), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n203), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n191), .A2(KEYINPUT1), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n219), .A2(new_n187), .A3(G143), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT67), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n187), .A2(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n223), .B(new_n224), .C1(new_n196), .C2(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n217), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n204), .A2(G134), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n208), .A2(G137), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n213), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(KEYINPUT30), .A3(new_n231), .ZN(new_n232));
  OR2_X1    g046(.A1(KEYINPUT2), .A2(G113), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT2), .A2(G113), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G116), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OR2_X1    g054(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n240), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n195), .C1(new_n197), .C2(new_n198), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n199), .A2(KEYINPUT65), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n214), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n231), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n232), .B(new_n244), .C1(new_n249), .C2(KEYINPUT30), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n243), .B(KEYINPUT69), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n215), .A3(new_n231), .ZN(new_n252));
  INV_X1    g066(.A(G237), .ZN(new_n253));
  INV_X1    g067(.A(G953), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G210), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n255), .B(KEYINPUT27), .Z(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT26), .ZN(new_n257));
  INV_X1    g071(.A(G101), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n250), .A2(new_n252), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT31), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT31), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n250), .A2(new_n262), .A3(new_n252), .A4(new_n259), .ZN(new_n263));
  INV_X1    g077(.A(new_n259), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n231), .A2(new_n248), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n244), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n265), .B1(new_n267), .B2(new_n252), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n252), .A2(new_n265), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n264), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n261), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(G472), .A2(G902), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT32), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n268), .A2(new_n270), .A3(new_n264), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n259), .B1(new_n250), .B2(new_n252), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n276), .A2(new_n277), .A3(KEYINPUT29), .ZN(new_n278));
  INV_X1    g092(.A(new_n252), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n251), .B1(new_n215), .B2(new_n231), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT28), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n281), .A2(KEYINPUT29), .A3(new_n259), .A4(new_n269), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(G472), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n272), .A2(KEYINPUT32), .A3(new_n273), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n275), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G217), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n288), .B1(G234), .B2(new_n283), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G125), .B(G140), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT16), .ZN(new_n292));
  INV_X1    g106(.A(G140), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G125), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(KEYINPUT16), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(new_n187), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n236), .A2(G128), .ZN(new_n297));
  OR2_X1    g111(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n236), .A2(G128), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G110), .ZN(new_n302));
  INV_X1    g116(.A(new_n299), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(new_n297), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT24), .B(G110), .Z(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n296), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n291), .A2(new_n187), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n308), .B(KEYINPUT70), .Z(new_n309));
  OR2_X1    g123(.A1(new_n295), .A2(new_n187), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n301), .A2(G110), .B1(new_n304), .B2(new_n305), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n254), .A2(G221), .A3(G234), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT22), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(G137), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n307), .B2(new_n312), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(KEYINPUT25), .B1(new_n320), .B2(new_n283), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(KEYINPUT25), .A3(new_n283), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n290), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n289), .A2(G902), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n324), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n287), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT71), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n331));
  INV_X1    g145(.A(G125), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n226), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n226), .B2(new_n332), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT79), .B(G224), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n254), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n199), .A2(G125), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n335), .A2(KEYINPUT7), .A3(new_n337), .A4(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G122), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(KEYINPUT8), .Z(new_n341));
  INV_X1    g155(.A(G107), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT73), .B1(new_n342), .B2(G104), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT73), .ZN(new_n344));
  INV_X1    g158(.A(G104), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(G107), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n345), .B2(G107), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n342), .A2(KEYINPUT3), .A3(G104), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n351), .A3(new_n258), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n342), .A2(G104), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n345), .A2(G107), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT5), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n357), .B(G113), .C1(KEYINPUT5), .C2(new_n237), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n241), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n241), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n352), .A2(new_n355), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n341), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n196), .A2(new_n219), .A3(G128), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n189), .A2(G146), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n216), .B1(new_n365), .B2(new_n222), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n224), .B1(new_n366), .B2(new_n223), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n218), .A2(KEYINPUT67), .A3(new_n220), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n332), .B(new_n364), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT78), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n226), .A2(new_n331), .A3(new_n332), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n338), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n337), .A2(KEYINPUT7), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n363), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n339), .A2(new_n374), .A3(KEYINPUT80), .ZN(new_n375));
  AOI21_X1  g189(.A(KEYINPUT80), .B1(new_n339), .B2(new_n374), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n347), .A2(new_n351), .A3(new_n258), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT74), .A2(G101), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(new_n347), .B2(new_n351), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT4), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n379), .A2(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n244), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n359), .ZN(new_n384));
  INV_X1    g198(.A(new_n340), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n375), .A2(new_n376), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n330), .B1(new_n387), .B2(G902), .ZN(new_n388));
  INV_X1    g202(.A(new_n386), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n385), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(KEYINPUT6), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n372), .B(new_n337), .Z(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n393), .A3(new_n385), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n376), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n339), .A2(new_n374), .A3(KEYINPUT80), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n389), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(KEYINPUT81), .A3(new_n283), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n388), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G210), .B1(G237), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n388), .A2(new_n399), .A3(new_n401), .A4(new_n395), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G475), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(new_n345), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n253), .A2(new_n254), .A3(G214), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(G143), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n410), .A2(new_n212), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n212), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n413));
  OR3_X1    g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n410), .B(new_n212), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n413), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n291), .B(KEYINPUT19), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n187), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n414), .A2(new_n416), .A3(new_n310), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n309), .B1(new_n187), .B2(new_n291), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT18), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n421), .A2(new_n212), .A3(KEYINPUT82), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n410), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n408), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n295), .B(G146), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n412), .A2(KEYINPUT17), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(KEYINPUT17), .C2(new_n415), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n408), .B(KEYINPUT84), .Z(new_n429));
  AND3_X1   g243(.A1(new_n428), .A2(new_n424), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n406), .B(new_n283), .C1(new_n425), .C2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n408), .B1(new_n428), .B2(new_n424), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n283), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G475), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n431), .A2(new_n432), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OR2_X1    g252(.A1(KEYINPUT87), .A2(G952), .ZN(new_n439));
  NAND2_X1  g253(.A1(KEYINPUT87), .A2(G952), .ZN(new_n440));
  AOI21_X1  g254(.A(G953), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G234), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n253), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(G898), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT88), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI211_X1 g261(.A(new_n283), .B(new_n254), .C1(G234), .C2(G237), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XOR2_X1   g263(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(G128), .A3(new_n189), .ZN(new_n451));
  XNOR2_X1  g265(.A(G128), .B(G143), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n451), .B(G134), .C1(new_n453), .C2(new_n450), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n208), .ZN(new_n455));
  INV_X1    g269(.A(G122), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G116), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n238), .A2(G122), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT85), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(new_n342), .ZN(new_n464));
  AOI21_X1  g278(.A(G107), .B1(new_n460), .B2(new_n462), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n454), .B(new_n455), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n465), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n452), .B(new_n208), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n458), .A2(KEYINPUT14), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n457), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n458), .A2(KEYINPUT14), .ZN(new_n471));
  OAI21_X1  g285(.A(G107), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n468), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT9), .B(G234), .Z(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n476), .A2(new_n288), .A3(G953), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n466), .A2(new_n473), .A3(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n283), .ZN(new_n482));
  INV_X1    g296(.A(G478), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT15), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n482), .B(new_n484), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n438), .A2(new_n449), .A3(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n405), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT71), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n327), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n203), .A2(new_n382), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n364), .A2(new_n366), .A3(new_n223), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n356), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT10), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n214), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n356), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n490), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT75), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n226), .A2(new_n361), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n203), .A2(new_n382), .B1(new_n500), .B2(KEYINPUT10), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(KEYINPUT75), .A3(new_n495), .A4(new_n494), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n492), .B1(new_n227), .B2(new_n356), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(new_n214), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT12), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G110), .B(G140), .ZN(new_n508));
  INV_X1    g322(.A(G227), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(G953), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n508), .B(new_n510), .Z(new_n511));
  NAND3_X1  g325(.A1(new_n503), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT76), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n501), .A2(new_n494), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n214), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n503), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n511), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n503), .A2(new_n507), .A3(new_n519), .A4(new_n511), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G469), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n283), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n511), .B1(new_n503), .B2(new_n507), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G469), .ZN(new_n527));
  NAND2_X1  g341(.A1(G469), .A2(G902), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n523), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G214), .B1(G237), .B2(G902), .ZN(new_n530));
  XOR2_X1   g344(.A(new_n530), .B(KEYINPUT77), .Z(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G221), .B1(new_n476), .B2(G902), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT72), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n529), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n329), .A2(new_n487), .A3(new_n489), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT89), .B(G101), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(G3));
  AND2_X1   g353(.A1(new_n529), .A2(new_n535), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n272), .A2(new_n283), .ZN(new_n541));
  NAND2_X1  g355(.A1(KEYINPUT90), .A2(G472), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n540), .A2(new_n326), .A3(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n449), .A2(new_n531), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n403), .A2(new_n546), .A3(new_n404), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n404), .A2(new_n546), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n550));
  AOI21_X1  g364(.A(G478), .B1(new_n481), .B2(new_n283), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT93), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT33), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT92), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n553), .A2(KEYINPUT92), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n481), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n479), .A2(KEYINPUT92), .A3(new_n553), .A4(new_n480), .ZN(new_n557));
  AOI211_X1 g371(.A(new_n483), .B(G902), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT94), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n551), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n557), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(G478), .A3(new_n283), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n550), .B1(new_n559), .B2(new_n565), .ZN(new_n566));
  AND4_X1   g380(.A1(new_n544), .A2(new_n545), .A3(new_n549), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT34), .B(G104), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(G6));
  INV_X1    g383(.A(new_n544), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n550), .A2(new_n485), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n549), .A2(new_n571), .A3(new_n545), .A4(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n547), .A2(new_n548), .A3(new_n545), .A4(new_n573), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT95), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n570), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT35), .B(G107), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G9));
  INV_X1    g393(.A(new_n323), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n289), .B1(new_n580), .B2(new_n321), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n317), .A2(KEYINPUT36), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n313), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n325), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n543), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n543), .A2(KEYINPUT96), .A3(new_n585), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n588), .A2(new_n487), .A3(new_n536), .A4(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT97), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT37), .B(G110), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G12));
  INV_X1    g407(.A(G900), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n448), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n443), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n596), .B(KEYINPUT98), .Z(new_n597));
  NOR2_X1   g411(.A1(new_n572), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n585), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n549), .A2(new_n287), .A3(new_n600), .A4(new_n536), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G128), .ZN(G30));
  AND3_X1   g416(.A1(new_n438), .A2(new_n532), .A3(new_n485), .ZN(new_n603));
  INV_X1    g417(.A(new_n584), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n324), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g420(.A(new_n606), .B(KEYINPUT100), .Z(new_n607));
  XOR2_X1   g421(.A(new_n597), .B(KEYINPUT39), .Z(new_n608));
  NAND2_X1  g422(.A1(new_n540), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT40), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n250), .A2(new_n252), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n264), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n279), .A2(new_n280), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n283), .B1(new_n613), .B2(new_n259), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n275), .A2(new_n286), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT99), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n405), .B(new_n619), .ZN(new_n620));
  OR4_X1    g434(.A1(new_n607), .A2(new_n610), .A3(new_n618), .A4(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G143), .ZN(G45));
  NOR2_X1   g436(.A1(new_n605), .A2(new_n597), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n566), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n549), .A2(new_n287), .A3(new_n536), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G146), .ZN(G48));
  AOI21_X1  g441(.A(new_n522), .B1(new_n521), .B2(new_n283), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n535), .A3(new_n523), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n327), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n549), .A2(new_n631), .A3(new_n545), .A4(new_n566), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT41), .B(G113), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G15));
  INV_X1    g448(.A(new_n631), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n574), .B2(new_n576), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT101), .B(G116), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G18));
  INV_X1    g452(.A(new_n523), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n628), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n547), .A2(new_n640), .A3(new_n548), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n287), .A2(new_n486), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n534), .A2(new_n531), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n641), .A2(new_n642), .A3(new_n585), .A4(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G119), .ZN(G21));
  AND3_X1   g459(.A1(new_n547), .A2(new_n548), .A3(new_n603), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n541), .A2(G472), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n281), .A2(new_n269), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n261), .B(new_n263), .C1(new_n648), .C2(new_n259), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n273), .B(KEYINPUT102), .Z(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n326), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n449), .ZN(new_n654));
  INV_X1    g468(.A(new_n630), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n646), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G122), .ZN(G24));
  NOR3_X1   g471(.A1(new_n647), .A2(new_n605), .A3(new_n651), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n559), .A2(new_n565), .ZN(new_n659));
  INV_X1    g473(.A(new_n597), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n438), .A3(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n641), .A2(new_n643), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G125), .ZN(G27));
  NAND3_X1  g479(.A1(new_n403), .A2(new_n532), .A3(new_n404), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(KEYINPUT103), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n403), .A2(new_n668), .A3(new_n532), .A4(new_n404), .ZN(new_n669));
  AND2_X1   g483(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n286), .A2(KEYINPUT104), .ZN(new_n671));
  INV_X1    g485(.A(new_n286), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n274), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n285), .B(new_n671), .C1(new_n673), .C2(KEYINPUT104), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n326), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n670), .A2(new_n675), .A3(new_n540), .A4(new_n662), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n328), .A2(new_n667), .A3(new_n540), .A4(new_n669), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n661), .A2(KEYINPUT42), .ZN(new_n679));
  AOI22_X1  g493(.A1(new_n676), .A2(KEYINPUT42), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G131), .ZN(G33));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n678), .B2(new_n598), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n677), .A2(KEYINPUT105), .A3(new_n572), .A4(new_n597), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G134), .ZN(G36));
  NAND2_X1  g500(.A1(new_n659), .A2(new_n550), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT43), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n688), .A2(new_n543), .A3(new_n605), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n670), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT106), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n526), .B(KEYINPUT45), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT46), .B1(new_n696), .B2(new_n528), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n639), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(KEYINPUT46), .A3(new_n528), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n535), .A3(new_n608), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n692), .A2(new_n703), .A3(new_n670), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n694), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT107), .B(G137), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G39));
  NAND2_X1  g521(.A1(new_n700), .A2(new_n535), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT47), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n287), .A2(new_n661), .A3(new_n326), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n670), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT108), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n293), .ZN(G42));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n536), .A2(new_n287), .A3(new_n548), .A4(new_n547), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n547), .A2(new_n548), .A3(new_n640), .A4(new_n643), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n658), .A2(new_n662), .ZN(new_n718));
  OAI22_X1  g532(.A1(new_n716), .A2(new_n599), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n716), .A2(new_n624), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT110), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n605), .A2(new_n723), .A3(new_n660), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT109), .B1(new_n585), .B2(new_n597), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n529), .A4(new_n535), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n646), .A2(new_n722), .A3(new_n616), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n547), .A2(new_n548), .A3(new_n603), .A4(new_n616), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT110), .B1(new_n729), .B2(new_n726), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n721), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n601), .A2(new_n664), .A3(new_n626), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n728), .A2(new_n730), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT52), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n644), .A2(new_n656), .A3(new_n632), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n636), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n733), .A2(new_n736), .A3(new_n738), .A4(new_n680), .ZN(new_n739));
  INV_X1    g553(.A(new_n566), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n572), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n741), .A2(new_n405), .A3(new_n545), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n544), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(new_n537), .A3(new_n590), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n287), .A2(new_n623), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n745), .A2(new_n485), .A3(new_n438), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n670), .B(new_n540), .C1(new_n663), .C2(new_n746), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n744), .B(new_n747), .C1(new_n684), .C2(new_n683), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n715), .B1(new_n739), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT112), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n715), .B1(new_n748), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n736), .A2(new_n738), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n733), .A2(new_n680), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n685), .A2(KEYINPUT112), .A3(new_n747), .A4(new_n744), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n753), .A2(new_n754), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(KEYINPUT111), .B(new_n715), .C1(new_n739), .C2(new_n748), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n751), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(KEYINPUT54), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n739), .A2(new_n748), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT53), .B1(new_n719), .B2(KEYINPUT52), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n749), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n760), .B1(KEYINPUT54), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n688), .A2(new_n443), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n326), .A3(new_n652), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n620), .A2(new_n531), .A3(new_n655), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT114), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT50), .ZN(new_n772));
  INV_X1    g586(.A(new_n670), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n630), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n326), .A3(new_n444), .A4(new_n618), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n775), .A2(new_n438), .A3(new_n659), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n774), .A2(new_n766), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(new_n658), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n772), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n640), .A2(new_n534), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT113), .Z(new_n782));
  AOI211_X1 g596(.A(new_n773), .B(new_n767), .C1(new_n709), .C2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(KEYINPUT115), .B(new_n765), .C1(new_n780), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n709), .A2(new_n781), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT117), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n767), .A2(new_n773), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n709), .A2(new_n788), .A3(new_n781), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n772), .A2(new_n779), .A3(KEYINPUT116), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT116), .B1(new_n772), .B2(new_n779), .ZN(new_n792));
  OAI211_X1 g606(.A(KEYINPUT51), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n777), .A2(new_n675), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n794), .A2(KEYINPUT48), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(KEYINPUT48), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n775), .A2(new_n740), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n795), .A2(new_n441), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n765), .B1(new_n780), .B2(new_n783), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n764), .A2(new_n784), .A3(new_n793), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n767), .A2(new_n717), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n802), .A2(new_n803), .B1(G952), .B2(G953), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT49), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n640), .A2(new_n805), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n639), .A2(KEYINPUT49), .A3(new_n628), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n806), .A2(new_n687), .A3(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n326), .A2(new_n643), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n618), .A2(new_n808), .A3(new_n620), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n804), .A2(new_n810), .ZN(G75));
  NOR2_X1   g625(.A1(new_n254), .A2(G952), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n759), .A2(G210), .A3(G902), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n391), .A2(new_n394), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n392), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT55), .Z(new_n819));
  AOI21_X1  g633(.A(KEYINPUT118), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n821));
  INV_X1    g635(.A(new_n819), .ZN(new_n822));
  AOI211_X1 g636(.A(new_n821), .B(new_n822), .C1(new_n814), .C2(new_n815), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n813), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n759), .A2(G902), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n759), .A2(KEYINPUT119), .A3(G902), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT120), .B1(new_n829), .B2(new_n402), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n759), .A2(KEYINPUT119), .A3(G902), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT119), .B1(new_n759), .B2(G902), .ZN(new_n832));
  OAI211_X1 g646(.A(KEYINPUT120), .B(new_n402), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n819), .A2(KEYINPUT56), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n824), .B1(new_n835), .B2(new_n836), .ZN(G51));
  XNOR2_X1  g651(.A(new_n521), .B(KEYINPUT121), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n759), .B(KEYINPUT54), .Z(new_n839));
  XNOR2_X1  g653(.A(new_n528), .B(KEYINPUT57), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n829), .A2(G469), .A3(new_n695), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n812), .B1(new_n841), .B2(new_n842), .ZN(G54));
  NAND3_X1  g657(.A1(new_n829), .A2(KEYINPUT58), .A3(G475), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n425), .A2(new_n430), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n829), .A2(KEYINPUT58), .A3(G475), .A4(new_n845), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n847), .A2(new_n813), .A3(new_n848), .ZN(G60));
  INV_X1    g663(.A(new_n563), .ZN(new_n850));
  XNOR2_X1  g664(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n483), .A2(new_n283), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n851), .B(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n850), .B1(new_n764), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n813), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n839), .A2(new_n850), .A3(new_n853), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(G63));
  NAND2_X1  g671(.A1(G217), .A2(G902), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT60), .Z(new_n859));
  XOR2_X1   g673(.A(new_n583), .B(KEYINPUT123), .Z(new_n860));
  NAND3_X1  g674(.A1(new_n759), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n813), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT61), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n320), .B1(new_n759), .B2(new_n859), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n864), .B(new_n866), .Z(G66));
  AOI21_X1  g681(.A(new_n254), .B1(new_n446), .B2(new_n336), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n738), .A2(new_n744), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n869), .B2(new_n254), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT125), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n817), .B1(G898), .B2(new_n254), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n871), .B(new_n872), .ZN(G69));
  NAND2_X1  g687(.A1(new_n621), .A2(new_n721), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT62), .Z(new_n875));
  NOR2_X1   g689(.A1(new_n773), .A2(new_n609), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n489), .A3(new_n329), .A4(new_n741), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n705), .A3(new_n712), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n232), .B1(new_n249), .B2(KEYINPUT30), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT126), .Z(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(new_n417), .Z(new_n881));
  NAND3_X1  g695(.A1(new_n878), .A2(new_n254), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n594), .B1(new_n881), .B2(new_n509), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n694), .A2(new_n704), .B1(new_n646), .B2(new_n675), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n680), .B(new_n685), .C1(new_n884), .C2(new_n701), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n712), .A2(new_n721), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n254), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(G227), .B2(new_n254), .ZN(new_n889));
  OAI221_X1 g703(.A(new_n882), .B1(new_n254), .B2(new_n883), .C1(new_n889), .C2(new_n881), .ZN(G72));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n891));
  NAND2_X1  g705(.A1(G472), .A2(G902), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT63), .Z(new_n893));
  OAI211_X1 g707(.A(new_n891), .B(new_n893), .C1(new_n887), .C2(new_n869), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n885), .A2(new_n869), .A3(new_n886), .ZN(new_n895));
  INV_X1    g709(.A(new_n893), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT127), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n894), .A2(new_n611), .A3(new_n897), .A4(new_n264), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n611), .B2(new_n264), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n763), .B(new_n899), .C1(new_n611), .C2(new_n264), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n893), .B1(new_n878), .B2(new_n869), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n612), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n813), .A2(new_n898), .A3(new_n900), .A4(new_n902), .ZN(G57));
endmodule


