

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U557 ( .A(n820), .B(KEYINPUT102), .ZN(n822) );
  OR2_X1 U558 ( .A1(n608), .A2(n607), .ZN(n610) );
  INV_X1 U559 ( .A(KEYINPUT17), .ZN(n546) );
  NAND2_X1 U560 ( .A1(n524), .A2(n525), .ZN(n523) );
  INV_X1 U561 ( .A(KEYINPUT33), .ZN(n524) );
  XOR2_X1 U562 ( .A(n773), .B(n772), .Z(n525) );
  XNOR2_X1 U563 ( .A(n548), .B(n547), .ZN(n559) );
  XNOR2_X1 U564 ( .A(n546), .B(KEYINPUT66), .ZN(n548) );
  AND2_X1 U565 ( .A1(n766), .A2(n986), .ZN(n767) );
  INV_X1 U566 ( .A(KEYINPUT64), .ZN(n772) );
  AND2_X1 U567 ( .A1(n979), .A2(n527), .ZN(n775) );
  NAND2_X1 U568 ( .A1(n665), .A2(G54), .ZN(n601) );
  XNOR2_X1 U569 ( .A(n561), .B(n560), .ZN(n562) );
  INV_X1 U570 ( .A(KEYINPUT67), .ZN(n560) );
  NOR2_X1 U571 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U572 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U573 ( .A1(n832), .A2(n825), .ZN(n526) );
  NAND2_X1 U574 ( .A1(n698), .A2(G40), .ZN(n700) );
  NOR2_X2 U575 ( .A1(n702), .A2(n982), .ZN(n711) );
  OR2_X1 U576 ( .A1(n746), .A2(n774), .ZN(n527) );
  NOR2_X1 U577 ( .A1(n746), .A2(n770), .ZN(n528) );
  XOR2_X1 U578 ( .A(n783), .B(KEYINPUT94), .Z(n529) );
  NOR2_X1 U579 ( .A1(n734), .A2(n963), .ZN(n701) );
  INV_X1 U580 ( .A(KEYINPUT29), .ZN(n727) );
  BUF_X1 U581 ( .A(n734), .Z(n747) );
  INV_X1 U582 ( .A(KEYINPUT101), .ZN(n768) );
  INV_X1 U583 ( .A(KEYINPUT88), .ZN(n699) );
  INV_X1 U584 ( .A(KEYINPUT75), .ZN(n600) );
  AND2_X1 U585 ( .A1(n784), .A2(n529), .ZN(n785) );
  XNOR2_X1 U586 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X1 U587 ( .A1(G164), .A2(G1384), .ZN(n788) );
  INV_X1 U588 ( .A(G2105), .ZN(n553) );
  INV_X1 U589 ( .A(KEYINPUT15), .ZN(n609) );
  XOR2_X2 U590 ( .A(G543), .B(KEYINPUT0), .Z(n647) );
  INV_X1 U591 ( .A(G651), .ZN(n537) );
  NOR2_X2 U592 ( .A1(n647), .A2(n537), .ZN(n662) );
  NAND2_X1 U593 ( .A1(G76), .A2(n662), .ZN(n534) );
  XOR2_X1 U594 ( .A(KEYINPUT77), .B(KEYINPUT4), .Z(n532) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n530) );
  XOR2_X2 U596 ( .A(KEYINPUT65), .B(n530), .Z(n661) );
  NAND2_X1 U597 ( .A1(G89), .A2(n661), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(KEYINPUT5), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT78), .B(n536), .ZN(n543) );
  NOR2_X4 U602 ( .A1(G651), .A2(n647), .ZN(n665) );
  NAND2_X1 U603 ( .A1(G51), .A2(n665), .ZN(n540) );
  NOR2_X1 U604 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X2 U605 ( .A(KEYINPUT1), .B(n538), .Z(n666) );
  NAND2_X1 U606 ( .A1(G63), .A2(n666), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n541), .Z(n542) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n545) );
  XOR2_X1 U610 ( .A(KEYINPUT79), .B(KEYINPUT7), .Z(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G168) );
  INV_X1 U612 ( .A(G2104), .ZN(n552) );
  NOR2_X4 U613 ( .A1(G2105), .A2(n552), .ZN(n891) );
  NAND2_X1 U614 ( .A1(n891), .A2(G102), .ZN(n551) );
  NOR2_X1 U615 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  INV_X1 U616 ( .A(n559), .ZN(n549) );
  INV_X2 U617 ( .A(n549), .ZN(n892) );
  NAND2_X1 U618 ( .A1(G138), .A2(n892), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n557) );
  NOR2_X2 U620 ( .A1(n552), .A2(n553), .ZN(n895) );
  NAND2_X1 U621 ( .A1(G114), .A2(n895), .ZN(n555) );
  NOR2_X2 U622 ( .A1(G2104), .A2(n553), .ZN(n896) );
  NAND2_X1 U623 ( .A1(G126), .A2(n896), .ZN(n554) );
  NAND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(G164) );
  NAND2_X1 U626 ( .A1(G101), .A2(n891), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT23), .B(n558), .Z(n563) );
  NAND2_X1 U628 ( .A1(n559), .A2(G137), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G113), .A2(n895), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G125), .A2(n896), .ZN(n564) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X2 U633 ( .A1(n567), .A2(n566), .ZN(n698) );
  BUF_X1 U634 ( .A(n698), .Z(G160) );
  NAND2_X1 U635 ( .A1(n666), .A2(G64), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT69), .B(n569), .Z(n571) );
  NAND2_X1 U637 ( .A1(n665), .A2(G52), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(KEYINPUT70), .B(n572), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G90), .A2(n661), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G77), .A2(n662), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n575), .Z(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(G171) );
  AND2_X1 U645 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U646 ( .A1(G123), .A2(n896), .ZN(n578) );
  XNOR2_X1 U647 ( .A(n578), .B(KEYINPUT18), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n891), .A2(G99), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G135), .A2(n892), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n895), .A2(G111), .ZN(n581) );
  XOR2_X1 U652 ( .A(KEYINPUT80), .B(n581), .Z(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n1023) );
  XNOR2_X1 U655 ( .A(G2096), .B(n1023), .ZN(n586) );
  OR2_X1 U656 ( .A1(G2100), .A2(n586), .ZN(G156) );
  INV_X1 U657 ( .A(G57), .ZN(G237) );
  INV_X1 U658 ( .A(G132), .ZN(G219) );
  INV_X1 U659 ( .A(G82), .ZN(G220) );
  XOR2_X1 U660 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n588) );
  NAND2_X1 U661 ( .A1(G7), .A2(G661), .ZN(n587) );
  XOR2_X1 U662 ( .A(n588), .B(n587), .Z(n932) );
  NAND2_X1 U663 ( .A1(n932), .A2(G567), .ZN(n589) );
  XOR2_X1 U664 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  NAND2_X1 U665 ( .A1(n661), .A2(G81), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U667 ( .A1(G68), .A2(n662), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n593), .B(KEYINPUT13), .ZN(n599) );
  NAND2_X1 U670 ( .A1(G43), .A2(n665), .ZN(n594) );
  XOR2_X1 U671 ( .A(KEYINPUT74), .B(n594), .Z(n597) );
  NAND2_X1 U672 ( .A1(n666), .A2(G56), .ZN(n595) );
  XOR2_X1 U673 ( .A(KEYINPUT14), .B(n595), .Z(n596) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n982) );
  INV_X1 U675 ( .A(G860), .ZN(n623) );
  OR2_X1 U676 ( .A1(n982), .A2(n623), .ZN(G153) );
  INV_X1 U677 ( .A(G171), .ZN(G301) );
  NAND2_X1 U678 ( .A1(G868), .A2(G301), .ZN(n612) );
  NAND2_X1 U679 ( .A1(n662), .A2(G79), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U681 ( .A(KEYINPUT76), .B(n604), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G92), .A2(n661), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G66), .A2(n666), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X2 U685 ( .A(n610), .B(n609), .ZN(n712) );
  INV_X1 U686 ( .A(G868), .ZN(n671) );
  NAND2_X1 U687 ( .A1(n712), .A2(n671), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(G284) );
  NAND2_X1 U689 ( .A1(n665), .A2(G53), .ZN(n613) );
  XOR2_X1 U690 ( .A(KEYINPUT71), .B(n613), .Z(n615) );
  NAND2_X1 U691 ( .A1(n666), .A2(G65), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U693 ( .A(KEYINPUT72), .B(n616), .Z(n620) );
  NAND2_X1 U694 ( .A1(G91), .A2(n661), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G78), .A2(n662), .ZN(n617) );
  AND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(G299) );
  NOR2_X1 U698 ( .A1(G286), .A2(n671), .ZN(n622) );
  NOR2_X1 U699 ( .A1(G868), .A2(G299), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n622), .A2(n621), .ZN(G297) );
  NAND2_X1 U701 ( .A1(n623), .A2(G559), .ZN(n624) );
  INV_X1 U702 ( .A(n712), .ZN(n998) );
  NAND2_X1 U703 ( .A1(n624), .A2(n998), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n625), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U705 ( .A1(G868), .A2(n982), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G868), .A2(n998), .ZN(n626) );
  NOR2_X1 U707 ( .A1(G559), .A2(n626), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(G282) );
  NAND2_X1 U709 ( .A1(n998), .A2(G559), .ZN(n679) );
  XNOR2_X1 U710 ( .A(n982), .B(n679), .ZN(n629) );
  NOR2_X1 U711 ( .A1(n629), .A2(G860), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G55), .A2(n665), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G67), .A2(n666), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G93), .A2(n661), .ZN(n633) );
  NAND2_X1 U716 ( .A1(G80), .A2(n662), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n674) );
  XNOR2_X1 U719 ( .A(n636), .B(n674), .ZN(G145) );
  NAND2_X1 U720 ( .A1(G85), .A2(n661), .ZN(n638) );
  NAND2_X1 U721 ( .A1(G72), .A2(n662), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U723 ( .A1(G47), .A2(n665), .ZN(n639) );
  XOR2_X1 U724 ( .A(KEYINPUT68), .B(n639), .Z(n640) );
  NOR2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U726 ( .A1(n666), .A2(G60), .ZN(n642) );
  NAND2_X1 U727 ( .A1(n643), .A2(n642), .ZN(G290) );
  NAND2_X1 U728 ( .A1(G49), .A2(n665), .ZN(n645) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U731 ( .A1(n666), .A2(n646), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n647), .A2(G87), .ZN(n648) );
  NAND2_X1 U733 ( .A1(n649), .A2(n648), .ZN(G288) );
  NAND2_X1 U734 ( .A1(G48), .A2(n665), .ZN(n650) );
  XOR2_X1 U735 ( .A(KEYINPUT83), .B(n650), .Z(n659) );
  NAND2_X1 U736 ( .A1(G73), .A2(n662), .ZN(n651) );
  XNOR2_X1 U737 ( .A(n651), .B(KEYINPUT2), .ZN(n652) );
  XNOR2_X1 U738 ( .A(n652), .B(KEYINPUT82), .ZN(n654) );
  NAND2_X1 U739 ( .A1(G86), .A2(n661), .ZN(n653) );
  NAND2_X1 U740 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U741 ( .A1(G61), .A2(n666), .ZN(n655) );
  XNOR2_X1 U742 ( .A(KEYINPUT81), .B(n655), .ZN(n656) );
  NOR2_X1 U743 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U744 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U745 ( .A(n660), .B(KEYINPUT84), .ZN(G305) );
  NAND2_X1 U746 ( .A1(G88), .A2(n661), .ZN(n664) );
  NAND2_X1 U747 ( .A1(G75), .A2(n662), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n664), .A2(n663), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G50), .A2(n665), .ZN(n668) );
  NAND2_X1 U750 ( .A1(G62), .A2(n666), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U752 ( .A1(n670), .A2(n669), .ZN(G166) );
  INV_X1 U753 ( .A(G166), .ZN(G303) );
  NAND2_X1 U754 ( .A1(n671), .A2(n674), .ZN(n682) );
  XNOR2_X1 U755 ( .A(KEYINPUT19), .B(G290), .ZN(n672) );
  XNOR2_X1 U756 ( .A(n672), .B(G288), .ZN(n673) );
  XOR2_X1 U757 ( .A(n674), .B(n673), .Z(n676) );
  XOR2_X1 U758 ( .A(G305), .B(G303), .Z(n675) );
  XNOR2_X1 U759 ( .A(n676), .B(n675), .ZN(n677) );
  INV_X1 U760 ( .A(G299), .ZN(n723) );
  XOR2_X1 U761 ( .A(n677), .B(n723), .Z(n678) );
  XNOR2_X1 U762 ( .A(n678), .B(n982), .ZN(n908) );
  XOR2_X1 U763 ( .A(n908), .B(n679), .Z(n680) );
  NAND2_X1 U764 ( .A1(G868), .A2(n680), .ZN(n681) );
  NAND2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U766 ( .A(n683), .B(KEYINPUT85), .ZN(G295) );
  NAND2_X1 U767 ( .A1(G2078), .A2(G2084), .ZN(n684) );
  XOR2_X1 U768 ( .A(KEYINPUT20), .B(n684), .Z(n685) );
  NAND2_X1 U769 ( .A1(G2090), .A2(n685), .ZN(n686) );
  XNOR2_X1 U770 ( .A(KEYINPUT21), .B(n686), .ZN(n687) );
  NAND2_X1 U771 ( .A1(n687), .A2(G2072), .ZN(n688) );
  XNOR2_X1 U772 ( .A(KEYINPUT86), .B(n688), .ZN(G158) );
  XNOR2_X1 U773 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U774 ( .A1(G220), .A2(G219), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT22), .B(n689), .Z(n690) );
  NOR2_X1 U776 ( .A1(G218), .A2(n690), .ZN(n691) );
  NAND2_X1 U777 ( .A1(G96), .A2(n691), .ZN(n929) );
  NAND2_X1 U778 ( .A1(G2106), .A2(n929), .ZN(n695) );
  NAND2_X1 U779 ( .A1(G69), .A2(G120), .ZN(n692) );
  NOR2_X1 U780 ( .A1(G237), .A2(n692), .ZN(n693) );
  NAND2_X1 U781 ( .A1(G108), .A2(n693), .ZN(n930) );
  NAND2_X1 U782 ( .A1(G567), .A2(n930), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n862) );
  NAND2_X1 U784 ( .A1(G661), .A2(G483), .ZN(n696) );
  NOR2_X1 U785 ( .A1(n862), .A2(n696), .ZN(n697) );
  XOR2_X1 U786 ( .A(KEYINPUT87), .B(n697), .Z(n843) );
  NAND2_X1 U787 ( .A1(n843), .A2(G36), .ZN(G176) );
  XNOR2_X2 U788 ( .A(n700), .B(n699), .ZN(n787) );
  NAND2_X2 U789 ( .A1(n787), .A2(n788), .ZN(n734) );
  XOR2_X1 U790 ( .A(G1996), .B(KEYINPUT96), .Z(n963) );
  XNOR2_X1 U791 ( .A(n701), .B(KEYINPUT26), .ZN(n702) );
  INV_X1 U792 ( .A(n712), .ZN(n703) );
  NAND2_X1 U793 ( .A1(G1341), .A2(n747), .ZN(n710) );
  AND2_X1 U794 ( .A1(n703), .A2(n710), .ZN(n704) );
  AND2_X2 U795 ( .A1(n711), .A2(n704), .ZN(n705) );
  XNOR2_X1 U796 ( .A(n705), .B(KEYINPUT97), .ZN(n709) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n747), .ZN(n707) );
  INV_X1 U798 ( .A(n734), .ZN(n716) );
  NOR2_X1 U799 ( .A1(n716), .A2(G1348), .ZN(n706) );
  NOR2_X1 U800 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n721) );
  NAND2_X1 U805 ( .A1(n716), .A2(G2072), .ZN(n717) );
  XNOR2_X1 U806 ( .A(n717), .B(KEYINPUT27), .ZN(n719) );
  INV_X1 U807 ( .A(G1956), .ZN(n993) );
  NOR2_X1 U808 ( .A1(n993), .A2(n716), .ZN(n718) );
  NOR2_X1 U809 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n726) );
  NOR2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U813 ( .A(n724), .B(KEYINPUT28), .Z(n725) );
  NAND2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U815 ( .A(n728), .B(n727), .ZN(n733) );
  XOR2_X1 U816 ( .A(G2078), .B(KEYINPUT25), .Z(n964) );
  NOR2_X1 U817 ( .A1(n964), .A2(n747), .ZN(n729) );
  XNOR2_X1 U818 ( .A(n729), .B(KEYINPUT95), .ZN(n731) );
  OR2_X1 U819 ( .A1(G1961), .A2(n716), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n739) );
  NAND2_X1 U821 ( .A1(n739), .A2(G171), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n744) );
  NAND2_X1 U823 ( .A1(G8), .A2(n734), .ZN(n746) );
  NOR2_X1 U824 ( .A1(G1966), .A2(n746), .ZN(n760) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n734), .ZN(n756) );
  INV_X1 U826 ( .A(n756), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n735), .A2(G8), .ZN(n736) );
  OR2_X1 U828 ( .A1(n760), .A2(n736), .ZN(n737) );
  XNOR2_X1 U829 ( .A(KEYINPUT30), .B(n737), .ZN(n738) );
  NOR2_X1 U830 ( .A1(G168), .A2(n738), .ZN(n741) );
  NOR2_X1 U831 ( .A1(G171), .A2(n739), .ZN(n740) );
  NOR2_X1 U832 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U833 ( .A(KEYINPUT31), .B(n742), .Z(n743) );
  NAND2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n757) );
  NAND2_X1 U835 ( .A1(n757), .A2(G286), .ZN(n745) );
  XNOR2_X1 U836 ( .A(n745), .B(KEYINPUT98), .ZN(n752) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n746), .ZN(n749) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U839 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U840 ( .A1(n750), .A2(G303), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U842 ( .A1(n753), .A2(G8), .ZN(n755) );
  XOR2_X1 U843 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n754) );
  XNOR2_X1 U844 ( .A(n755), .B(n754), .ZN(n764) );
  NAND2_X1 U845 ( .A1(G8), .A2(n756), .ZN(n762) );
  BUF_X1 U846 ( .A(n757), .Z(n758) );
  INV_X1 U847 ( .A(n758), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n764), .A2(n763), .ZN(n776) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n765) );
  XOR2_X1 U852 ( .A(n765), .B(KEYINPUT100), .Z(n766) );
  NOR2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n985) );
  NAND2_X1 U854 ( .A1(n776), .A2(n767), .ZN(n769) );
  XNOR2_X1 U855 ( .A(n769), .B(n768), .ZN(n771) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U857 ( .A(n987), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n528), .ZN(n773) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n979) );
  NAND2_X1 U860 ( .A1(n985), .A2(KEYINPUT33), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n523), .A2(n775), .ZN(n786) );
  BUF_X1 U862 ( .A(n776), .Z(n779) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n777) );
  NAND2_X1 U864 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U866 ( .A1(n746), .A2(n780), .ZN(n784) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XOR2_X1 U868 ( .A(n781), .B(KEYINPUT24), .Z(n782) );
  NOR2_X1 U869 ( .A1(n746), .A2(n782), .ZN(n783) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n819) );
  INV_X1 U871 ( .A(n787), .ZN(n789) );
  NOR2_X1 U872 ( .A1(n789), .A2(n788), .ZN(n835) );
  XNOR2_X1 U873 ( .A(KEYINPUT37), .B(G2067), .ZN(n823) );
  XNOR2_X1 U874 ( .A(KEYINPUT91), .B(KEYINPUT36), .ZN(n801) );
  NAND2_X1 U875 ( .A1(n891), .A2(G104), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G140), .A2(n892), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n792), .B(KEYINPUT34), .ZN(n793) );
  XNOR2_X1 U879 ( .A(n793), .B(KEYINPUT89), .ZN(n799) );
  XNOR2_X1 U880 ( .A(KEYINPUT90), .B(KEYINPUT35), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G116), .A2(n895), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G128), .A2(n896), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U884 ( .A(n797), .B(n796), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U886 ( .A(n801), .B(n800), .ZN(n903) );
  NOR2_X1 U887 ( .A1(n823), .A2(n903), .ZN(n1026) );
  NAND2_X1 U888 ( .A1(n835), .A2(n1026), .ZN(n832) );
  NAND2_X1 U889 ( .A1(n895), .A2(G107), .ZN(n803) );
  NAND2_X1 U890 ( .A1(G131), .A2(n892), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U892 ( .A1(n891), .A2(G95), .ZN(n804) );
  XOR2_X1 U893 ( .A(KEYINPUT92), .B(n804), .Z(n805) );
  NOR2_X1 U894 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U895 ( .A1(n896), .A2(G119), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n881) );
  NAND2_X1 U897 ( .A1(n881), .A2(G1991), .ZN(n818) );
  NAND2_X1 U898 ( .A1(G105), .A2(n891), .ZN(n809) );
  XOR2_X1 U899 ( .A(KEYINPUT38), .B(n809), .Z(n814) );
  NAND2_X1 U900 ( .A1(G117), .A2(n895), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G129), .A2(n896), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U903 ( .A(KEYINPUT93), .B(n812), .Z(n813) );
  NOR2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n816) );
  NAND2_X1 U905 ( .A1(G141), .A2(n892), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n879) );
  NAND2_X1 U907 ( .A1(n879), .A2(G1996), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n1008) );
  NAND2_X1 U909 ( .A1(n1008), .A2(n835), .ZN(n825) );
  AND2_X2 U910 ( .A1(n819), .A2(n526), .ZN(n820) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U912 ( .A1(n990), .A2(n835), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n838) );
  NAND2_X1 U914 ( .A1(n823), .A2(n903), .ZN(n1009) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n879), .ZN(n824) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n824), .Z(n1017) );
  INV_X1 U917 ( .A(n825), .ZN(n828) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n881), .ZN(n1022) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n826) );
  NOR2_X1 U920 ( .A1(n1022), .A2(n826), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n1017), .A2(n829), .ZN(n830) );
  XNOR2_X1 U923 ( .A(KEYINPUT104), .B(n830), .ZN(n831) );
  XNOR2_X1 U924 ( .A(n831), .B(KEYINPUT39), .ZN(n833) );
  NAND2_X1 U925 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n1009), .A2(n834), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U928 ( .A1(n838), .A2(n837), .ZN(n840) );
  XOR2_X1 U929 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n839) );
  XNOR2_X1 U930 ( .A(n840), .B(n839), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n932), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U933 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U935 ( .A1(n843), .A2(n842), .ZN(G188) );
  XOR2_X1 U936 ( .A(G2100), .B(G2096), .Z(n845) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n844) );
  XNOR2_X1 U938 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n847) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U941 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U942 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n850) );
  XNOR2_X1 U944 ( .A(n851), .B(n850), .ZN(G227) );
  XNOR2_X1 U945 ( .A(G1971), .B(n993), .ZN(n853) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1961), .ZN(n852) );
  XNOR2_X1 U947 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U948 ( .A(G1966), .B(G1976), .Z(n855) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U950 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U951 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U952 ( .A(KEYINPUT109), .B(G2474), .ZN(n858) );
  XNOR2_X1 U953 ( .A(n859), .B(n858), .ZN(n861) );
  XOR2_X1 U954 ( .A(G1981), .B(KEYINPUT41), .Z(n860) );
  XNOR2_X1 U955 ( .A(n861), .B(n860), .ZN(G229) );
  XOR2_X1 U956 ( .A(KEYINPUT108), .B(n862), .Z(G319) );
  NAND2_X1 U957 ( .A1(G124), .A2(n896), .ZN(n863) );
  XNOR2_X1 U958 ( .A(n863), .B(KEYINPUT44), .ZN(n864) );
  XNOR2_X1 U959 ( .A(n864), .B(KEYINPUT110), .ZN(n866) );
  NAND2_X1 U960 ( .A1(G112), .A2(n895), .ZN(n865) );
  NAND2_X1 U961 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U962 ( .A1(n891), .A2(G100), .ZN(n868) );
  NAND2_X1 U963 ( .A1(G136), .A2(n892), .ZN(n867) );
  NAND2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U965 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U966 ( .A(KEYINPUT111), .B(n871), .Z(G162) );
  NAND2_X1 U967 ( .A1(G118), .A2(n895), .ZN(n873) );
  NAND2_X1 U968 ( .A1(G130), .A2(n896), .ZN(n872) );
  NAND2_X1 U969 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U970 ( .A1(n891), .A2(G106), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G142), .A2(n892), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U973 ( .A(n876), .B(KEYINPUT45), .Z(n877) );
  NOR2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n880) );
  XNOR2_X1 U975 ( .A(n880), .B(n879), .ZN(n890) );
  XNOR2_X1 U976 ( .A(G162), .B(n881), .ZN(n882) );
  XNOR2_X1 U977 ( .A(n882), .B(n1023), .ZN(n886) );
  XOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n884) );
  XNOR2_X1 U979 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U980 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U981 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U982 ( .A(G160), .B(G164), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n905) );
  NAND2_X1 U985 ( .A1(n891), .A2(G103), .ZN(n894) );
  NAND2_X1 U986 ( .A1(G139), .A2(n892), .ZN(n893) );
  NAND2_X1 U987 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U988 ( .A1(G115), .A2(n895), .ZN(n898) );
  NAND2_X1 U989 ( .A1(G127), .A2(n896), .ZN(n897) );
  NAND2_X1 U990 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U991 ( .A(KEYINPUT112), .B(n899), .Z(n900) );
  XNOR2_X1 U992 ( .A(KEYINPUT47), .B(n900), .ZN(n901) );
  NOR2_X1 U993 ( .A1(n902), .A2(n901), .ZN(n1011) );
  XNOR2_X1 U994 ( .A(n903), .B(n1011), .ZN(n904) );
  XNOR2_X1 U995 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U996 ( .A1(G37), .A2(n906), .ZN(G395) );
  XOR2_X1 U997 ( .A(G301), .B(G286), .Z(n907) );
  XNOR2_X1 U998 ( .A(n907), .B(KEYINPUT115), .ZN(n910) );
  XNOR2_X1 U999 ( .A(n998), .B(n908), .ZN(n909) );
  XNOR2_X1 U1000 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n911), .ZN(G397) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n912) );
  XNOR2_X1 U1004 ( .A(n913), .B(n912), .ZN(n926) );
  XNOR2_X1 U1005 ( .A(G2454), .B(G2446), .ZN(n922) );
  XNOR2_X1 U1006 ( .A(G2430), .B(G2443), .ZN(n920) );
  XOR2_X1 U1007 ( .A(G2435), .B(KEYINPUT106), .Z(n915) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2438), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n915), .B(n914), .ZN(n916) );
  XOR2_X1 U1010 ( .A(n916), .B(G2427), .Z(n918) );
  XNOR2_X1 U1011 ( .A(G1341), .B(G1348), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(n918), .B(n917), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(n922), .B(n921), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(n923), .A2(G14), .ZN(n924) );
  XOR2_X1 U1016 ( .A(KEYINPUT107), .B(n924), .Z(n931) );
  NAND2_X1 U1017 ( .A1(n931), .A2(G319), .ZN(n925) );
  NOR2_X1 U1018 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(G225) );
  XNOR2_X1 U1021 ( .A(KEYINPUT117), .B(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(G120), .ZN(G236) );
  INV_X1 U1024 ( .A(G96), .ZN(G221) );
  INV_X1 U1025 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(G325) );
  INV_X1 U1027 ( .A(G325), .ZN(G261) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  INV_X1 U1029 ( .A(n931), .ZN(G401) );
  INV_X1 U1030 ( .A(n932), .ZN(G223) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G21), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(G1961), .B(G5), .ZN(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n946) );
  XOR2_X1 U1034 ( .A(G1981), .B(G6), .Z(n939) );
  XOR2_X1 U1035 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n936) );
  XNOR2_X1 U1036 ( .A(KEYINPUT59), .B(G4), .ZN(n935) );
  XNOR2_X1 U1037 ( .A(n936), .B(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(G1348), .B(n937), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n943) );
  XOR2_X1 U1040 ( .A(G1341), .B(G19), .Z(n941) );
  XOR2_X1 U1041 ( .A(G1956), .B(G20), .Z(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(n944), .B(KEYINPUT60), .ZN(n945) );
  NAND2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G1986), .B(G24), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(G22), .B(G1971), .ZN(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1049 ( .A(G1976), .B(KEYINPUT127), .ZN(n949) );
  XNOR2_X1 U1050 ( .A(n949), .B(G23), .ZN(n950) );
  NAND2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1052 ( .A(KEYINPUT58), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1054 ( .A(KEYINPUT61), .B(n955), .Z(n956) );
  NOR2_X1 U1055 ( .A1(G16), .A2(n956), .ZN(n1039) );
  XOR2_X1 U1056 ( .A(G29), .B(KEYINPUT122), .Z(n977) );
  XOR2_X1 U1057 ( .A(G2090), .B(G35), .Z(n959) );
  XOR2_X1 U1058 ( .A(G34), .B(KEYINPUT54), .Z(n957) );
  XNOR2_X1 U1059 ( .A(n957), .B(G2084), .ZN(n958) );
  NAND2_X1 U1060 ( .A1(n959), .A2(n958), .ZN(n974) );
  XOR2_X1 U1061 ( .A(G1991), .B(G25), .Z(n960) );
  NAND2_X1 U1062 ( .A1(n960), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1063 ( .A(G2067), .B(G26), .ZN(n962) );
  XNOR2_X1 U1064 ( .A(G33), .B(G2072), .ZN(n961) );
  NOR2_X1 U1065 ( .A1(n962), .A2(n961), .ZN(n968) );
  XOR2_X1 U1066 ( .A(n963), .B(G32), .Z(n966) );
  XNOR2_X1 U1067 ( .A(G27), .B(n964), .ZN(n965) );
  NOR2_X1 U1068 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1071 ( .A(KEYINPUT121), .B(n971), .Z(n972) );
  XNOR2_X1 U1072 ( .A(n972), .B(KEYINPUT53), .ZN(n973) );
  NOR2_X1 U1073 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1074 ( .A(n975), .B(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1075 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1076 ( .A1(G11), .A2(n978), .ZN(n1007) );
  XNOR2_X1 U1077 ( .A(KEYINPUT56), .B(G16), .ZN(n1004) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n980) );
  NAND2_X1 U1079 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1080 ( .A(n981), .B(KEYINPUT57), .ZN(n1002) );
  XOR2_X1 U1081 ( .A(G171), .B(G1961), .Z(n984) );
  XNOR2_X1 U1082 ( .A(n982), .B(G1341), .ZN(n983) );
  NOR2_X1 U1083 ( .A1(n984), .A2(n983), .ZN(n997) );
  XOR2_X1 U1084 ( .A(G303), .B(G1971), .Z(n992) );
  INV_X1 U1085 ( .A(n985), .ZN(n986) );
  NAND2_X1 U1086 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1087 ( .A(KEYINPUT123), .B(n988), .Z(n989) );
  NOR2_X1 U1088 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1089 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1090 ( .A(n993), .B(G299), .Z(n994) );
  NOR2_X1 U1091 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1092 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1093 ( .A(G1348), .B(n998), .Z(n999) );
  NOR2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1097 ( .A(KEYINPUT124), .B(n1005), .Z(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1037) );
  INV_X1 U1099 ( .A(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1031) );
  XOR2_X1 U1101 ( .A(n1011), .B(KEYINPUT119), .Z(n1012) );
  XOR2_X1 U1102 ( .A(G2072), .B(n1012), .Z(n1014) );
  XOR2_X1 U1103 ( .A(G164), .B(G2078), .Z(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1105 ( .A(KEYINPUT50), .B(n1015), .Z(n1020) );
  XOR2_X1 U1106 ( .A(G2090), .B(G162), .Z(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(KEYINPUT51), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1029) );
  XOR2_X1 U1110 ( .A(G160), .B(G2084), .Z(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1114 ( .A(n1027), .B(KEYINPUT118), .ZN(n1028) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1117 ( .A(KEYINPUT52), .B(n1032), .Z(n1033) );
  NOR2_X1 U1118 ( .A1(KEYINPUT55), .A2(n1033), .ZN(n1034) );
  XOR2_X1 U1119 ( .A(KEYINPUT120), .B(n1034), .Z(n1035) );
  NAND2_X1 U1120 ( .A1(G29), .A2(n1035), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1122 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1040), .Z(G150) );
  INV_X1 U1124 ( .A(G150), .ZN(G311) );
endmodule

