//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  OR3_X1    g0023(.A1(new_n209), .A2(KEYINPUT64), .A3(G13), .ZN(new_n224));
  OAI21_X1  g0024(.A(KEYINPUT64), .B1(new_n209), .B2(G13), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n207), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n223), .B(new_n228), .C1(new_n230), .C2(new_n233), .ZN(G361));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XOR2_X1   g0045(.A(G58), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XOR2_X1   g0048(.A(G107), .B(G116), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT73), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT10), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n252), .A2(KEYINPUT10), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  AND2_X1   g0055(.A1(new_n255), .A2(new_n229), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT8), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n207), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT68), .ZN(new_n263));
  XNOR2_X1  g0063(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n256), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n255), .A2(new_n229), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT69), .B1(new_n207), .B2(G1), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT69), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(new_n206), .A3(G20), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n202), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT70), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(new_n277), .B2(new_n276), .ZN(new_n279));
  AOI211_X1 g0079(.A(new_n268), .B(new_n279), .C1(new_n202), .C2(new_n270), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT9), .ZN(new_n281));
  INV_X1    g0081(.A(G41), .ZN(new_n282));
  INV_X1    g0082(.A(G45), .ZN(new_n283));
  AOI21_X1  g0083(.A(G1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n284), .A2(new_n286), .A3(G274), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G222), .A2(G1698), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G223), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT3), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n286), .B1(new_n301), .B2(new_n217), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n291), .B1(new_n296), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G190), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n304), .B1(new_n305), .B2(new_n303), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n253), .B(new_n254), .C1(new_n281), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n280), .B(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n306), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n309), .A2(new_n252), .A3(KEYINPUT10), .A4(new_n310), .ZN(new_n311));
  AND2_X1   g0111(.A1(KEYINPUT71), .A2(G179), .ZN(new_n312));
  NOR2_X1   g0112(.A1(KEYINPUT71), .A2(G179), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n303), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G169), .B2(new_n303), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n280), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n307), .A2(new_n311), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n260), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n266), .B1(G20), .B2(G77), .ZN(new_n321));
  XOR2_X1   g0121(.A(KEYINPUT15), .B(G87), .Z(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n262), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n271), .B1(new_n217), .B2(new_n270), .ZN(new_n325));
  AOI211_X1 g0125(.A(new_n271), .B(new_n270), .C1(new_n275), .C2(new_n273), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G77), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n292), .A2(G232), .A3(new_n294), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n219), .B2(new_n292), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n301), .A2(new_n212), .A3(new_n294), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n287), .ZN(new_n334));
  INV_X1    g0134(.A(new_n289), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n334), .B1(G244), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n328), .B1(new_n338), .B2(G169), .ZN(new_n339));
  INV_X1    g0139(.A(new_n314), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n327), .B(new_n325), .C1(new_n338), .C2(new_n305), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT72), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n344), .A2(new_n345), .B1(new_n348), .B2(new_n337), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n319), .B(new_n343), .C1(new_n347), .C2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n292), .B2(G20), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n301), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n211), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n258), .A2(new_n211), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n356), .B2(new_n201), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n266), .A2(G159), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n351), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT78), .ZN(new_n361));
  INV_X1    g0161(.A(new_n359), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT77), .B1(new_n299), .B2(G33), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n297), .A3(KEYINPUT3), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n365), .A3(new_n300), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(new_n352), .A3(new_n207), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G68), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n352), .B1(new_n366), .B2(new_n207), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT16), .B(new_n362), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n371), .B(new_n351), .C1(new_n355), .C2(new_n359), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n361), .A2(new_n271), .A3(new_n370), .A4(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(new_n261), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n269), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n326), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n334), .B1(G232), .B2(new_n335), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n290), .A2(G1698), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(G223), .B2(G1698), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n366), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n382), .B(KEYINPUT79), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n329), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n340), .ZN(new_n386));
  INV_X1    g0186(.A(G169), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n385), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n377), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT18), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT18), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n377), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n305), .B1(new_n378), .B2(new_n384), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(G190), .B2(new_n385), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n373), .A2(new_n394), .A3(new_n376), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n373), .A2(new_n394), .A3(KEYINPUT17), .A4(new_n376), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n390), .A2(new_n392), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n264), .A2(G77), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n266), .A2(G50), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n207), .B2(G68), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n271), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT11), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n270), .A2(new_n211), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT12), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n326), .A2(G68), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n290), .A2(new_n294), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n294), .A2(G232), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n292), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(G33), .A2(G97), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n329), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT13), .ZN(new_n417));
  INV_X1    g0217(.A(G274), .ZN(new_n418));
  INV_X1    g0218(.A(new_n229), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n419), .B2(new_n285), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n335), .A2(G238), .B1(new_n420), .B2(new_n284), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n416), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n286), .B1(new_n413), .B2(new_n414), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n287), .B1(new_n289), .B2(new_n212), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT13), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n416), .A2(new_n421), .A3(KEYINPUT74), .A4(new_n417), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(G169), .A4(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT75), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n422), .A2(new_n425), .A3(G179), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n427), .A2(G169), .A3(new_n429), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n410), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n427), .A2(G200), .A3(new_n429), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n422), .A2(G190), .A3(new_n425), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n410), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n350), .A2(new_n399), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(G238), .A2(G1698), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n218), .B2(G1698), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(new_n363), .A3(new_n300), .A4(new_n365), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G116), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n286), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n283), .A2(G1), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n420), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n214), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n286), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT84), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n218), .A2(G1698), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(G238), .B2(G1698), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n450), .B1(new_n366), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n329), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n453), .A2(new_n455), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT84), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n457), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G200), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n322), .A2(new_n269), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n207), .B1(new_n414), .B2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT85), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(G97), .A2(G107), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n213), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT85), .B(new_n207), .C1(new_n414), .C2(new_n468), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G97), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n468), .B1(new_n262), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n363), .A2(new_n365), .A3(new_n207), .A4(new_n300), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n475), .B(new_n477), .C1(new_n211), .C2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n256), .B1(new_n479), .B2(KEYINPUT86), .ZN(new_n480));
  AND3_X1   g0280(.A1(new_n363), .A2(new_n365), .A3(new_n300), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n207), .A3(G68), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT86), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n475), .A4(new_n477), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n467), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n206), .A2(G33), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n269), .A2(new_n486), .A3(new_n229), .A4(new_n255), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G87), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n457), .A2(new_n464), .A3(G190), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n466), .A2(new_n485), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n465), .A2(new_n387), .ZN(new_n492));
  INV_X1    g0292(.A(new_n475), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n477), .B1(new_n478), .B2(new_n211), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT86), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n271), .A3(new_n484), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n488), .A2(new_n322), .ZN(new_n497));
  INV_X1    g0297(.A(new_n467), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n457), .A2(new_n464), .A3(new_n314), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n492), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n491), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G20), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n271), .B(new_n504), .C1(KEYINPUT87), .C2(KEYINPUT20), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n207), .B1(new_n476), .B2(G33), .ZN(new_n506));
  INV_X1    g0306(.A(G283), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT80), .B1(new_n297), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT80), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n509), .A2(G33), .A3(G283), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT87), .B(KEYINPUT20), .C1(new_n505), .C2(new_n511), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n207), .A2(G116), .B1(KEYINPUT87), .B2(KEYINPUT20), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n256), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(KEYINPUT87), .A2(KEYINPUT20), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n508), .A2(new_n510), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n514), .B(new_n515), .C1(new_n517), .C2(new_n506), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n269), .A2(new_n503), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n488), .B2(new_n503), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n512), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n220), .A2(G1698), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(G257), .B2(G1698), .ZN(new_n523));
  INV_X1    g0323(.A(G303), .ZN(new_n524));
  OAI22_X1  g0324(.A1(new_n366), .A2(new_n523), .B1(new_n524), .B2(new_n292), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n329), .ZN(new_n526));
  AND2_X1   g0326(.A1(KEYINPUT5), .A2(G41), .ZN(new_n527));
  NOR2_X1   g0327(.A1(KEYINPUT5), .A2(G41), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n452), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n286), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G270), .ZN(new_n532));
  OR2_X1    g0332(.A1(new_n527), .A2(new_n528), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n533), .A2(new_n420), .A3(new_n452), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n526), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n521), .B1(new_n535), .B2(G200), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n348), .B2(new_n535), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n526), .A2(new_n532), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(G179), .A3(new_n521), .A4(new_n534), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n521), .A3(G169), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(KEYINPUT21), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n537), .B(new_n539), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n540), .B(KEYINPUT21), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT88), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n539), .A4(new_n537), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n502), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n298), .A2(new_n300), .A3(G250), .A4(G1698), .ZN(new_n549));
  AND2_X1   g0349(.A1(KEYINPUT4), .A2(G244), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n298), .A2(new_n300), .A3(new_n550), .A4(new_n294), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n516), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n218), .A2(G1698), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n363), .A2(new_n365), .A3(new_n300), .A4(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n286), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n529), .A2(G257), .A3(new_n286), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT81), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT81), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n529), .A2(new_n560), .A3(G257), .A4(new_n286), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n534), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G190), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n476), .A2(new_n219), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(new_n472), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n219), .A2(KEYINPUT6), .A3(G97), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(G20), .B1(G77), .B2(new_n266), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n353), .A2(new_n354), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G107), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n256), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n270), .A2(new_n476), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n487), .B2(new_n476), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(G200), .B1(new_n557), .B2(new_n562), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n564), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT82), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n387), .B1(new_n557), .B2(new_n562), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n554), .A2(new_n555), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n549), .A2(new_n516), .A3(new_n551), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n329), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n561), .A2(new_n534), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n584), .A2(new_n314), .A3(new_n559), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT83), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n563), .A2(KEYINPUT83), .A3(new_n314), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n576), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n579), .B1(new_n590), .B2(new_n578), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n580), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT89), .ZN(new_n594));
  NAND2_X1  g0394(.A1(KEYINPUT22), .A2(G87), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n478), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n213), .A2(G20), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT22), .B1(new_n292), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n594), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT22), .ZN(new_n600));
  INV_X1    g0400(.A(new_n597), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n301), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(KEYINPUT89), .C1(new_n478), .C2(new_n595), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n219), .A2(KEYINPUT23), .A3(G20), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT23), .B1(new_n219), .B2(G20), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n605), .A2(new_n606), .B1(G20), .B2(new_n450), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n593), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  AOI211_X1 g0409(.A(KEYINPUT24), .B(new_n607), .C1(new_n599), .C2(new_n603), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n271), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT25), .B1(new_n270), .B2(new_n219), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n270), .A2(KEYINPUT25), .A3(new_n219), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(G107), .B2(new_n488), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT90), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n214), .A2(new_n294), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n619), .B1(G257), .B2(new_n294), .ZN(new_n620));
  INV_X1    g0420(.A(G294), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n366), .A2(new_n620), .B1(new_n297), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n329), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n531), .A2(G264), .ZN(new_n624));
  AND4_X1   g0424(.A1(G179), .A2(new_n623), .A3(new_n534), .A4(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n623), .B(new_n534), .C1(new_n220), .C2(new_n530), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n387), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n611), .A2(KEYINPUT90), .A3(new_n615), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n618), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n627), .A2(new_n348), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(G200), .B2(new_n627), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n633), .A2(new_n611), .A3(new_n615), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n548), .A2(new_n592), .A3(new_n631), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n446), .A2(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n580), .A2(new_n591), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n629), .B2(new_n616), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n461), .A2(new_n462), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n387), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n499), .A2(new_n500), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(G200), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n485), .A2(new_n489), .A3(new_n490), .A4(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n634), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n637), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n644), .A2(new_n642), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n588), .A2(new_n589), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n576), .B1(new_n648), .B2(KEYINPUT91), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT91), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n588), .A2(new_n651), .A3(new_n589), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n647), .A2(new_n649), .A3(new_n650), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n590), .A2(new_n491), .A3(new_n501), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(new_n642), .A3(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n646), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n445), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n317), .ZN(new_n659));
  INV_X1    g0459(.A(new_n392), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n391), .B1(new_n377), .B2(new_n388), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n437), .B(new_n435), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n410), .A2(new_n665), .B1(new_n443), .B2(new_n342), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n397), .A2(new_n398), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n662), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n307), .A2(new_n311), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n659), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n658), .A2(new_n671), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n544), .A2(new_n547), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(G343), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n521), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n638), .A2(new_n521), .A3(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n631), .A2(new_n634), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n618), .A2(new_n630), .A3(new_n679), .ZN(new_n688));
  INV_X1    g0488(.A(new_n679), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n687), .A2(new_n688), .B1(new_n631), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n631), .A2(new_n634), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n679), .B1(new_n545), .B2(new_n539), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n616), .A2(new_n629), .A3(new_n689), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0499(.A(new_n226), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  NOR4_X1   g0501(.A1(new_n701), .A2(new_n206), .A3(G116), .A4(new_n473), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n233), .B2(new_n701), .ZN(new_n703));
  XOR2_X1   g0503(.A(new_n703), .B(KEYINPUT28), .Z(new_n704));
  NOR2_X1   g0504(.A1(new_n628), .A2(new_n563), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n640), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n461), .A2(new_n462), .A3(KEYINPUT93), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n707), .A2(new_n314), .A3(new_n535), .A4(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(KEYINPUT94), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(KEYINPUT94), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n705), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n625), .A2(new_n563), .A3(new_n538), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n465), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT95), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n714), .A2(new_n713), .A3(new_n465), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n719), .B(new_n713), .C1(new_n714), .C2(new_n465), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n712), .A2(new_n716), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n679), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n712), .A2(new_n718), .A3(new_n715), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n724), .B(new_n726), .C1(new_n635), .C2(new_n679), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n648), .A2(KEYINPUT91), .ZN(new_n730));
  INV_X1    g0530(.A(new_n576), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n652), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n644), .A2(new_n642), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT26), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n642), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT97), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n734), .A2(new_n735), .A3(KEYINPUT97), .A4(new_n642), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n637), .A2(new_n645), .ZN(new_n740));
  INV_X1    g0540(.A(new_n631), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(new_n638), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n743), .A2(KEYINPUT98), .A3(new_n689), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT98), .B1(new_n743), .B2(new_n689), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT29), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n657), .A2(new_n689), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n729), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n704), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(G13), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n206), .B1(new_n753), .B2(G45), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n701), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT101), .Z(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n387), .A2(KEYINPUT102), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n207), .B1(KEYINPUT102), .B2(new_n387), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n229), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n247), .A2(G45), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT100), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n700), .A2(new_n481), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n768), .B(new_n769), .C1(G45), .C2(new_n232), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n700), .A2(new_n301), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n771), .A2(G355), .B1(new_n503), .B2(new_n700), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n766), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n207), .A2(new_n305), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n340), .A2(G190), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT104), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n775), .A2(KEYINPUT104), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(new_n348), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n340), .A2(new_n305), .A3(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n207), .A2(G190), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n340), .A2(new_n305), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G58), .A2(new_n783), .B1(new_n786), .B2(G77), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n780), .A2(G50), .B1(KEYINPUT103), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G179), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n781), .A2(new_n789), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G179), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G190), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n292), .B1(new_n790), .B2(new_n213), .C1(new_n794), .C2(new_n476), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n784), .A2(new_n789), .A3(G200), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n219), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n340), .A2(new_n348), .A3(new_n774), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n795), .B(new_n800), .C1(G68), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n784), .A2(new_n791), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G159), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT105), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n787), .A2(KEYINPUT103), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n788), .A2(new_n803), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n799), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n811), .A2(G283), .B1(new_n786), .B2(G311), .ZN(new_n812));
  INV_X1    g0612(.A(G329), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n301), .B1(new_n804), .B2(new_n813), .C1(new_n790), .C2(new_n524), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G294), .B2(new_n793), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT107), .B(G326), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n812), .B(new_n815), .C1(new_n779), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  XOR2_X1   g0618(.A(KEYINPUT33), .B(G317), .Z(new_n819));
  OAI22_X1  g0619(.A1(new_n818), .A2(new_n782), .B1(new_n801), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT108), .Z(new_n821));
  OAI21_X1  g0621(.A(new_n810), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n757), .B(new_n773), .C1(new_n764), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n760), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n823), .B1(new_n683), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n683), .A2(G330), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n757), .B1(new_n684), .B2(new_n685), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n342), .A2(new_n689), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n328), .A2(new_n679), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n349), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n346), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n830), .B1(new_n834), .B2(new_n342), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n747), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n830), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n831), .B1(new_n347), .B2(new_n349), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(new_n838), .B2(new_n343), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n689), .B(new_n839), .C1(new_n646), .C2(new_n656), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n729), .A2(new_n836), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT109), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n836), .A2(new_n840), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n756), .B1(new_n843), .B2(new_n728), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n759), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n846), .A2(new_n764), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n757), .B1(new_n217), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n811), .A2(G87), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G116), .A2(new_n786), .B1(new_n802), .B2(G283), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n849), .B(new_n850), .C1(new_n621), .C2(new_n782), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n779), .A2(new_n524), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n794), .A2(new_n476), .ZN(new_n853));
  INV_X1    g0653(.A(G311), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n301), .B1(new_n804), .B2(new_n854), .C1(new_n790), .C2(new_n219), .ZN(new_n855));
  NOR4_X1   g0655(.A1(new_n851), .A2(new_n852), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G150), .A2(new_n802), .B1(new_n786), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G143), .ZN(new_n858));
  INV_X1    g0658(.A(G137), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n857), .B1(new_n858), .B2(new_n782), .C1(new_n779), .C2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT34), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n794), .A2(new_n258), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n481), .B1(new_n863), .B2(new_n804), .C1(new_n202), .C2(new_n790), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n862), .B(new_n864), .C1(new_n811), .C2(G68), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n856), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n764), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n848), .B1(new_n866), .B2(new_n867), .C1(new_n839), .C2(new_n759), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n845), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G384));
  NOR2_X1   g0670(.A1(new_n753), .A2(new_n206), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n746), .A2(new_n445), .A3(new_n749), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n671), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n389), .A2(KEYINPUT112), .ZN(new_n874));
  XOR2_X1   g0674(.A(KEYINPUT113), .B(KEYINPUT37), .Z(new_n875));
  AND2_X1   g0675(.A1(new_n395), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n677), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n377), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT112), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n377), .A2(new_n388), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n874), .A2(new_n876), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n362), .B1(new_n368), .B2(new_n369), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n882), .A2(new_n351), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n370), .A2(new_n271), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n376), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n388), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n877), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(new_n395), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT37), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n881), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n887), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n399), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n439), .A2(new_n679), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n890), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n399), .A2(new_n377), .A3(new_n877), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n389), .A2(new_n878), .A3(new_n395), .ZN(new_n901));
  INV_X1    g0701(.A(new_n875), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n881), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT38), .B1(new_n900), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n899), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n897), .B(new_n898), .C1(new_n906), .C2(KEYINPUT39), .ZN(new_n907));
  INV_X1    g0707(.A(new_n662), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n677), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n895), .A2(new_n896), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n410), .A2(new_n679), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n439), .A2(new_n443), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n410), .B(new_n679), .C1(new_n665), .C2(new_n442), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n840), .A2(KEYINPUT111), .A3(new_n830), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT111), .B1(new_n840), .B2(new_n830), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n911), .B(new_n915), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n910), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n873), .B(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n881), .A2(new_n903), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n878), .B1(new_n662), .B2(new_n667), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n894), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n896), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT31), .B1(new_n721), .B2(new_n679), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n693), .A2(new_n592), .A3(new_n548), .A4(new_n689), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n835), .B1(new_n913), .B2(new_n914), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n924), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n915), .A2(new_n839), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n928), .B2(new_n927), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT40), .B1(new_n895), .B2(new_n896), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n931), .A2(KEYINPUT40), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n929), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n935), .B1(new_n446), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n548), .A2(new_n592), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n938), .A2(new_n687), .A3(new_n679), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n724), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n930), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT40), .B1(new_n942), .B2(new_n906), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n933), .A2(new_n934), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(new_n445), .A3(new_n929), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n937), .A2(new_n946), .A3(G330), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n871), .B1(new_n920), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n920), .B2(new_n947), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n569), .A2(KEYINPUT35), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n950), .A2(G116), .A3(new_n230), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT36), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n232), .A2(new_n217), .A3(new_n356), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n211), .A2(G50), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT110), .Z(new_n956));
  OAI211_X1 g0756(.A(G1), .B(new_n752), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n949), .A2(new_n953), .A3(new_n957), .ZN(G367));
  NOR3_X1   g0758(.A1(new_n238), .A2(new_n700), .A3(new_n481), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n765), .B1(new_n226), .B2(new_n323), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n756), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n790), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(G116), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT46), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n219), .B2(new_n794), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G283), .A2(new_n786), .B1(new_n783), .B2(G303), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n476), .B2(new_n799), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n481), .B1(G317), .B2(new_n805), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n621), .B2(new_n801), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n965), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n780), .A2(G311), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n780), .A2(G143), .ZN(new_n972));
  INV_X1    g0772(.A(G150), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n799), .A2(new_n217), .B1(new_n973), .B2(new_n782), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n794), .A2(new_n211), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n292), .B1(new_n804), .B2(new_n859), .C1(new_n790), .C2(new_n258), .ZN(new_n976));
  INV_X1    g0776(.A(G159), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n202), .A2(new_n785), .B1(new_n801), .B2(new_n977), .ZN(new_n978));
  NOR4_X1   g0778(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n970), .A2(new_n971), .B1(new_n972), .B2(new_n979), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT47), .Z(new_n981));
  AOI21_X1  g0781(.A(new_n961), .B1(new_n981), .B2(new_n764), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n485), .A2(new_n489), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n679), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n647), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n642), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n982), .B1(new_n824), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT114), .B(KEYINPUT43), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(KEYINPUT43), .B2(new_n986), .ZN(new_n990));
  INV_X1    g0790(.A(new_n590), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n592), .B1(new_n576), .B2(new_n689), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n649), .A2(new_n652), .A3(new_n679), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n991), .B1(new_n995), .B2(new_n631), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n693), .A3(new_n694), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n996), .A2(new_n689), .B1(KEYINPUT42), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(KEYINPUT115), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n997), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n998), .A2(KEYINPUT115), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n990), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1002), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1004), .A2(new_n1000), .A3(new_n999), .A4(new_n989), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n691), .A2(new_n995), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1006), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n995), .A2(new_n697), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT44), .Z(new_n1011));
  NOR2_X1   g0811(.A1(new_n995), .A2(new_n697), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n692), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n691), .A3(new_n1013), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n695), .B1(new_n690), .B2(new_n694), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n686), .B(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n750), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n750), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n701), .B(KEYINPUT41), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n755), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n987), .B1(new_n1009), .B2(new_n1023), .ZN(G387));
  OR2_X1    g0824(.A1(new_n690), .A2(new_n824), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n769), .B1(new_n242), .B2(new_n283), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n473), .A2(G116), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n771), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OR3_X1    g0829(.A1(new_n260), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(KEYINPUT50), .B1(new_n260), .B2(G50), .ZN(new_n1031));
  AOI21_X1  g0831(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1030), .A2(new_n1027), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1029), .A2(new_n1033), .B1(new_n219), .B2(new_n700), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n756), .B1(new_n1034), .B2(new_n766), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n780), .A2(G159), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n962), .A2(G77), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n973), .B2(new_n804), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n794), .A2(new_n323), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1038), .A2(new_n1039), .A3(new_n366), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n811), .A2(G97), .B1(G50), .B2(new_n783), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G68), .A2(new_n786), .B1(new_n802), .B2(new_n261), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1036), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G311), .A2(new_n802), .B1(new_n783), .B2(G317), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n524), .B2(new_n785), .C1(new_n779), .C2(new_n818), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n794), .A2(new_n507), .B1(new_n790), .B2(new_n621), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1050));
  NAND3_X1  g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n366), .B1(new_n816), .B2(new_n804), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n811), .B2(G116), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1050), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1043), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1035), .B1(new_n1056), .B2(new_n764), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1019), .A2(new_n755), .B1(new_n1025), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1020), .A2(new_n701), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n750), .A2(new_n1019), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(G393));
  AND2_X1   g0861(.A1(new_n769), .A2(new_n250), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n765), .B1(new_n476), .B2(new_n226), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n756), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n780), .A2(G317), .B1(G311), .B2(new_n783), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT117), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n301), .B1(new_n804), .B2(new_n818), .C1(new_n790), .C2(new_n507), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n800), .B1(G303), .B2(new_n802), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n621), .B2(new_n785), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1068), .B(new_n1070), .C1(G116), .C2(new_n793), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n779), .A2(new_n973), .B1(new_n977), .B2(new_n782), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT51), .Z(new_n1075));
  OAI221_X1 g0875(.A(new_n849), .B1(new_n202), .B2(new_n801), .C1(new_n260), .C2(new_n785), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n794), .A2(new_n217), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n481), .B1(new_n858), .B2(new_n804), .C1(new_n211), .C2(new_n790), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1072), .A2(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1064), .B1(new_n1080), .B2(new_n764), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n994), .B2(new_n824), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n701), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1082), .B1(new_n754), .B2(new_n1017), .C1(new_n1083), .C2(new_n1084), .ZN(G390));
  AOI21_X1  g0885(.A(new_n685), .B1(new_n927), .B2(new_n928), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n445), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n872), .A2(new_n671), .A3(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n727), .A2(G330), .A3(new_n839), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n915), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1086), .A2(new_n930), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n917), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n840), .A2(KEYINPUT111), .A3(new_n830), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n743), .A2(new_n689), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT98), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n743), .A2(KEYINPUT98), .A3(new_n689), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n830), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n834), .A2(new_n342), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n915), .B1(new_n1086), .B2(new_n839), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1095), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1088), .A2(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT39), .B1(new_n923), .B2(new_n896), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n898), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1100), .A2(new_n1102), .A3(new_n915), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n906), .A2(new_n898), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1114), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1104), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1108), .B(new_n1119), .C1(new_n1117), .C2(new_n1092), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n872), .A2(new_n671), .A3(new_n1087), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1095), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1117), .A2(new_n1092), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1104), .B(new_n1114), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1120), .A2(new_n1128), .A3(new_n701), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n757), .B1(new_n374), .B2(new_n847), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT118), .Z(new_n1131));
  NOR2_X1   g0931(.A1(new_n1111), .A2(new_n759), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1133));
  OR3_X1    g0933(.A1(new_n790), .A2(new_n1133), .A3(new_n973), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n790), .B2(new_n973), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n301), .B1(new_n805), .B2(G125), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n793), .A2(G159), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .A4(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT54), .B(G143), .Z(new_n1139));
  AOI22_X1  g0939(.A1(G132), .A2(new_n783), .B1(new_n786), .B2(new_n1139), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n202), .B2(new_n799), .C1(new_n859), .C2(new_n801), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1138), .B(new_n1141), .C1(G128), .C2(new_n780), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n292), .B1(new_n962), .B2(G87), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1143), .A2(KEYINPUT120), .B1(new_n783), .B2(G116), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(KEYINPUT120), .B2(new_n1143), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G97), .A2(new_n786), .B1(new_n802), .B2(G107), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1077), .B1(G294), .B2(new_n805), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n211), .C2(new_n799), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n1145), .B(new_n1148), .C1(G283), .C2(new_n780), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1131), .B(new_n1132), .C1(new_n764), .C2(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n1152), .B2(new_n755), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1129), .A2(new_n1153), .ZN(G378));
  AOI21_X1  g0954(.A(new_n1088), .B1(new_n1152), .B2(new_n1108), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n280), .A2(new_n677), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n318), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n307), .A2(new_n311), .A3(new_n317), .A4(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1160), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n945), .B2(G330), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n685), .B(new_n1163), .C1(new_n943), .C2(new_n944), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n919), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1163), .B1(new_n935), .B2(new_n685), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n918), .A2(new_n909), .A3(new_n907), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n945), .A2(G330), .A3(new_n1164), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1167), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT57), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n701), .B1(new_n1155), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT57), .B1(new_n1175), .B2(new_n1172), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1163), .A2(new_n846), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n780), .A2(G116), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1037), .B1(new_n507), .B2(new_n804), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n366), .A2(new_n282), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1180), .A2(new_n975), .A3(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n811), .A2(G58), .B1(G97), .B2(new_n802), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G107), .A2(new_n783), .B1(new_n786), .B2(new_n322), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT58), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G50), .B1(new_n297), .B2(new_n282), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1185), .A2(new_n1186), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G128), .A2(new_n783), .B1(new_n802), .B2(G132), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n962), .A2(new_n1139), .B1(new_n793), .B2(G150), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1191), .C1(new_n859), .C2(new_n785), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G125), .B2(new_n780), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT59), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1189), .B1(new_n977), .B2(new_n799), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1193), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1196), .A2(KEYINPUT59), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1188), .B1(new_n1186), .B2(new_n1185), .C1(new_n1195), .C2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n764), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n847), .A2(new_n202), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1178), .A2(new_n756), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n1172), .B2(new_n755), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1177), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1088), .A2(new_n1107), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1125), .A2(new_n1022), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1090), .A2(new_n846), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n846), .A2(G68), .A3(new_n764), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n780), .A2(G294), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n301), .B1(new_n804), .B2(new_n524), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n1212), .B(new_n1039), .C1(G97), .C2(new_n962), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n811), .A2(G77), .B1(G283), .B2(new_n783), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G107), .A2(new_n786), .B1(new_n802), .B2(G116), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n779), .A2(new_n863), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT122), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n790), .A2(new_n977), .B1(new_n804), .B2(new_n1219), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n366), .B(new_n1220), .C1(G50), .C2(new_n793), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n811), .A2(G58), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G137), .A2(new_n783), .B1(new_n802), .B2(new_n1139), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n786), .A2(G150), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1221), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1216), .B1(new_n1218), .B2(new_n1225), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n757), .B(new_n1210), .C1(new_n1226), .C2(new_n764), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1209), .A2(new_n1227), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n754), .B(KEYINPUT121), .Z(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1107), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1208), .A2(new_n1231), .ZN(G381));
  NOR2_X1   g1032(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1082), .B1(new_n1017), .B2(new_n754), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n869), .ZN(new_n1236));
  OR2_X1    g1036(.A1(G393), .A2(G396), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1236), .A2(G387), .A3(G381), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G378), .A2(KEYINPUT123), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT123), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1129), .A2(new_n1240), .A3(new_n1153), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(new_n1205), .A3(new_n1243), .ZN(G407));
  NAND2_X1  g1044(.A1(new_n678), .A2(G213), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT124), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1205), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G407), .A2(new_n1247), .A3(G213), .ZN(G409));
  INV_X1    g1048(.A(KEYINPUT127), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G390), .B(new_n987), .C1(new_n1023), .C2(new_n1009), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(G387), .A2(new_n1235), .ZN(new_n1251));
  XOR2_X1   g1051(.A(G393), .B(G396), .Z(new_n1252));
  AND3_X1   g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1249), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1252), .ZN(new_n1256));
  AND2_X1   g1056(.A1(G387), .A2(new_n1235), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(G387), .A2(new_n1235), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(KEYINPUT127), .A3(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1255), .A2(new_n1261), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1263));
  OAI211_X1 g1063(.A(new_n1022), .B(new_n1172), .C1(new_n1263), .C2(new_n1088), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1229), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1169), .B1(new_n1170), .B2(new_n1168), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1265), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT125), .B1(new_n1268), .B2(new_n1201), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1229), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT125), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1270), .A2(new_n1271), .A3(new_n1202), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1269), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1264), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1239), .A2(new_n1274), .A3(new_n1241), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G378), .B(new_n1203), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1088), .A2(new_n1107), .A3(KEYINPUT60), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1279), .A2(new_n701), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1107), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1207), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1283), .B2(new_n1231), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n869), .B(new_n1230), .C1(new_n1280), .C2(new_n1282), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1278), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1279), .A2(new_n701), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1207), .B2(new_n1281), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n869), .B1(new_n1288), .B2(new_n1230), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1283), .A2(G384), .A3(new_n1231), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(KEYINPUT126), .A3(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1286), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1277), .A2(new_n1245), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1246), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1294), .B1(new_n1286), .B2(new_n1291), .ZN(new_n1296));
  AOI22_X1  g1096(.A1(new_n1293), .A2(new_n1294), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n678), .A2(G213), .A3(G2897), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1284), .A2(new_n1285), .A3(new_n1278), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT126), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(G2897), .A3(new_n1246), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1298), .B1(new_n1305), .B2(new_n1295), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1262), .B1(new_n1297), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1259), .A2(new_n1298), .A3(new_n1260), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1292), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1308), .B1(new_n1295), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1293), .A2(new_n1310), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1277), .A2(new_n1245), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n1302), .A3(new_n1304), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1307), .A2(new_n1316), .ZN(G405));
  OAI211_X1 g1117(.A(new_n1303), .B(new_n1276), .C1(new_n1205), .C2(new_n1242), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1276), .B1(new_n1205), .B2(new_n1242), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1318), .B1(new_n1320), .B2(new_n1309), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(new_n1262), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1255), .A2(new_n1261), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1323), .B(new_n1318), .C1(new_n1309), .C2(new_n1320), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(G402));
endmodule


