

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U555 ( .A1(KEYINPUT33), .A2(n701), .ZN(n702) );
  OR2_X1 U556 ( .A1(n752), .A2(n751), .ZN(n773) );
  BUF_X1 U557 ( .A(n727), .Z(n728) );
  INV_X1 U558 ( .A(G2105), .ZN(n528) );
  BUF_X2 U559 ( .A(n637), .Z(n678) );
  NOR2_X1 U560 ( .A1(n653), .A2(n652), .ZN(n656) );
  INV_X1 U561 ( .A(KEYINPUT28), .ZN(n657) );
  NOR2_X2 U562 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  XNOR2_X1 U563 ( .A(KEYINPUT66), .B(G543), .ZN(n535) );
  XNOR2_X1 U564 ( .A(n550), .B(n549), .ZN(n552) );
  INV_X1 U565 ( .A(KEYINPUT23), .ZN(n549) );
  NAND2_X1 U566 ( .A1(G160), .A2(G40), .ZN(n523) );
  INV_X1 U567 ( .A(KEYINPUT26), .ZN(n638) );
  INV_X1 U568 ( .A(KEYINPUT30), .ZN(n667) );
  XNOR2_X1 U569 ( .A(n667), .B(KEYINPUT101), .ZN(n668) );
  XNOR2_X1 U570 ( .A(n669), .B(n668), .ZN(n670) );
  INV_X1 U571 ( .A(KEYINPUT0), .ZN(n534) );
  XNOR2_X1 U572 ( .A(n535), .B(n534), .ZN(n584) );
  BUF_X1 U573 ( .A(n608), .Z(G164) );
  XOR2_X2 U574 ( .A(KEYINPUT17), .B(n524), .Z(n905) );
  NAND2_X1 U575 ( .A1(n905), .A2(G138), .ZN(n527) );
  NOR2_X1 U576 ( .A1(G2104), .A2(n528), .ZN(n727) );
  NAND2_X1 U577 ( .A1(G126), .A2(n727), .ZN(n525) );
  XOR2_X1 U578 ( .A(KEYINPUT91), .B(n525), .Z(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n532) );
  AND2_X4 U580 ( .A1(n528), .A2(G2104), .ZN(n906) );
  NAND2_X1 U581 ( .A1(G102), .A2(n906), .ZN(n530) );
  AND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n909) );
  NAND2_X1 U583 ( .A1(G114), .A2(n909), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n608) );
  NOR2_X1 U586 ( .A1(G651), .A2(G543), .ZN(n817) );
  NAND2_X1 U587 ( .A1(n817), .A2(G89), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n533), .B(KEYINPUT4), .ZN(n537) );
  INV_X1 U589 ( .A(G651), .ZN(n539) );
  NOR2_X1 U590 ( .A1(n539), .A2(n584), .ZN(n615) );
  BUF_X1 U591 ( .A(n615), .Z(n818) );
  NAND2_X1 U592 ( .A1(G76), .A2(n818), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U594 ( .A(n538), .B(KEYINPUT5), .ZN(n547) );
  NOR2_X1 U595 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U596 ( .A(KEYINPUT1), .B(n540), .Z(n813) );
  NAND2_X1 U597 ( .A1(G63), .A2(n813), .ZN(n544) );
  NOR2_X1 U598 ( .A1(G651), .A2(n584), .ZN(n541) );
  XNOR2_X1 U599 ( .A(n541), .B(KEYINPUT64), .ZN(n613) );
  INV_X1 U600 ( .A(n613), .ZN(n542) );
  INV_X1 U601 ( .A(n542), .ZN(n814) );
  NAND2_X1 U602 ( .A1(G51), .A2(n814), .ZN(n543) );
  NAND2_X1 U603 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U608 ( .A(KEYINPUT65), .ZN(n554) );
  NAND2_X1 U609 ( .A1(n906), .A2(G101), .ZN(n550) );
  NAND2_X1 U610 ( .A1(n727), .A2(G125), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n554), .B(n553), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G137), .A2(n905), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G113), .A2(n909), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X2 U616 ( .A1(n558), .A2(n557), .ZN(G160) );
  NAND2_X1 U617 ( .A1(G90), .A2(n817), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G77), .A2(n818), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT9), .ZN(n566) );
  NAND2_X1 U621 ( .A1(G64), .A2(n813), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G52), .A2(n814), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U624 ( .A(KEYINPUT68), .B(n564), .Z(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(n567), .B(KEYINPUT69), .ZN(G171) );
  NAND2_X1 U627 ( .A1(G65), .A2(n813), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G53), .A2(n814), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT70), .B(n570), .Z(n574) );
  NAND2_X1 U631 ( .A1(G91), .A2(n817), .ZN(n572) );
  NAND2_X1 U632 ( .A1(G78), .A2(n818), .ZN(n571) );
  AND2_X1 U633 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(G299) );
  NAND2_X1 U635 ( .A1(n814), .A2(G50), .ZN(n575) );
  XNOR2_X1 U636 ( .A(n575), .B(KEYINPUT84), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G88), .A2(n817), .ZN(n577) );
  NAND2_X1 U638 ( .A1(G75), .A2(n818), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G62), .A2(n813), .ZN(n578) );
  XNOR2_X1 U641 ( .A(KEYINPUT83), .B(n578), .ZN(n579) );
  NOR2_X1 U642 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U644 ( .A(KEYINPUT85), .B(n583), .Z(G303) );
  INV_X1 U645 ( .A(G303), .ZN(G166) );
  NAND2_X1 U646 ( .A1(G87), .A2(n584), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G651), .A2(G74), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G49), .A2(n814), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U650 ( .A1(n813), .A2(n587), .ZN(n588) );
  NAND2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U652 ( .A(KEYINPUT81), .B(n590), .Z(G288) );
  NAND2_X1 U653 ( .A1(G86), .A2(n817), .ZN(n592) );
  NAND2_X1 U654 ( .A1(G61), .A2(n813), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT82), .B(n593), .ZN(n596) );
  NAND2_X1 U657 ( .A1(n818), .A2(G73), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT2), .B(n594), .Z(n595) );
  NOR2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U660 ( .A1(G48), .A2(n814), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(G305) );
  NAND2_X1 U662 ( .A1(G85), .A2(n817), .ZN(n600) );
  NAND2_X1 U663 ( .A1(G72), .A2(n818), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U665 ( .A(KEYINPUT67), .B(n601), .ZN(n605) );
  NAND2_X1 U666 ( .A1(n814), .A2(G47), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G60), .A2(n813), .ZN(n602) );
  AND2_X1 U668 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U669 ( .A1(n605), .A2(n604), .ZN(G290) );
  INV_X1 U670 ( .A(G40), .ZN(n606) );
  OR2_X1 U671 ( .A1(n606), .A2(G1384), .ZN(n607) );
  NOR2_X1 U672 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U673 ( .A1(G160), .A2(n609), .ZN(n637) );
  XOR2_X1 U674 ( .A(n637), .B(KEYINPUT100), .Z(n651) );
  XNOR2_X1 U675 ( .A(G2078), .B(KEYINPUT25), .ZN(n937) );
  NAND2_X1 U676 ( .A1(n651), .A2(n937), .ZN(n612) );
  INV_X1 U677 ( .A(G1961), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n610), .A2(n678), .ZN(n611) );
  NAND2_X1 U679 ( .A1(n612), .A2(n611), .ZN(n671) );
  NAND2_X1 U680 ( .A1(n671), .A2(G171), .ZN(n664) );
  NAND2_X1 U681 ( .A1(n613), .A2(G54), .ZN(n614) );
  XNOR2_X1 U682 ( .A(n614), .B(KEYINPUT76), .ZN(n618) );
  NAND2_X1 U683 ( .A1(n615), .A2(G79), .ZN(n616) );
  XOR2_X1 U684 ( .A(KEYINPUT75), .B(n616), .Z(n617) );
  NAND2_X1 U685 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U686 ( .A(n619), .B(KEYINPUT77), .ZN(n624) );
  AND2_X1 U687 ( .A1(G66), .A2(n813), .ZN(n622) );
  NAND2_X1 U688 ( .A1(n817), .A2(G92), .ZN(n620) );
  XOR2_X1 U689 ( .A(KEYINPUT74), .B(n620), .Z(n621) );
  NOR2_X1 U690 ( .A1(n622), .A2(n621), .ZN(n623) );
  AND2_X1 U691 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X2 U692 ( .A(KEYINPUT15), .B(n625), .Z(n1008) );
  NAND2_X1 U693 ( .A1(n813), .A2(G56), .ZN(n626) );
  XNOR2_X1 U694 ( .A(n626), .B(KEYINPUT14), .ZN(n633) );
  XNOR2_X1 U695 ( .A(KEYINPUT13), .B(KEYINPUT72), .ZN(n631) );
  NAND2_X1 U696 ( .A1(n817), .A2(G81), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n627), .B(KEYINPUT12), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G68), .A2(n818), .ZN(n628) );
  NAND2_X1 U699 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(n632) );
  NAND2_X1 U701 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(KEYINPUT73), .ZN(n636) );
  NAND2_X1 U703 ( .A1(G43), .A2(n814), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n1010) );
  INV_X1 U705 ( .A(G1996), .ZN(n934) );
  NOR2_X1 U706 ( .A1(n678), .A2(n934), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n641) );
  NAND2_X1 U708 ( .A1(n678), .A2(G1341), .ZN(n640) );
  NAND2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U710 ( .A1(n1010), .A2(n642), .ZN(n647) );
  NAND2_X1 U711 ( .A1(n1008), .A2(n647), .ZN(n646) );
  NAND2_X1 U712 ( .A1(G2067), .A2(n651), .ZN(n644) );
  NAND2_X1 U713 ( .A1(G1348), .A2(n678), .ZN(n643) );
  NAND2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U715 ( .A1(n646), .A2(n645), .ZN(n649) );
  OR2_X1 U716 ( .A1(n1008), .A2(n647), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n655) );
  INV_X1 U718 ( .A(G299), .ZN(n1023) );
  NAND2_X1 U719 ( .A1(G2072), .A2(n651), .ZN(n650) );
  XNOR2_X1 U720 ( .A(n650), .B(KEYINPUT27), .ZN(n653) );
  INV_X1 U721 ( .A(G1956), .ZN(n984) );
  NOR2_X1 U722 ( .A1(n651), .A2(n984), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n1023), .A2(n656), .ZN(n654) );
  NAND2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n660) );
  NOR2_X1 U725 ( .A1(n1023), .A2(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U727 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U728 ( .A(KEYINPUT29), .B(n661), .ZN(n662) );
  INV_X1 U729 ( .A(n662), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n676) );
  NAND2_X1 U731 ( .A1(n678), .A2(G8), .ZN(n722) );
  NOR2_X1 U732 ( .A1(G1966), .A2(n722), .ZN(n691) );
  NOR2_X1 U733 ( .A1(G2084), .A2(n678), .ZN(n665) );
  XOR2_X1 U734 ( .A(KEYINPUT99), .B(n665), .Z(n688) );
  NOR2_X1 U735 ( .A1(n691), .A2(n688), .ZN(n666) );
  NAND2_X1 U736 ( .A1(G8), .A2(n666), .ZN(n669) );
  NOR2_X1 U737 ( .A1(G168), .A2(n670), .ZN(n673) );
  NOR2_X1 U738 ( .A1(G171), .A2(n671), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U740 ( .A(KEYINPUT31), .B(n674), .Z(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n689) );
  NAND2_X1 U742 ( .A1(G286), .A2(n689), .ZN(n677) );
  XNOR2_X1 U743 ( .A(n677), .B(KEYINPUT102), .ZN(n685) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n722), .ZN(n680) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n678), .ZN(n679) );
  NOR2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(KEYINPUT103), .ZN(n682) );
  NOR2_X1 U748 ( .A1(G166), .A2(n682), .ZN(n683) );
  XOR2_X1 U749 ( .A(KEYINPUT104), .B(n683), .Z(n684) );
  NAND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n686), .A2(G8), .ZN(n687) );
  XNOR2_X1 U752 ( .A(n687), .B(KEYINPUT32), .ZN(n710) );
  NAND2_X1 U753 ( .A1(G8), .A2(n688), .ZN(n693) );
  INV_X1 U754 ( .A(n689), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n711) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n1021) );
  AND2_X1 U758 ( .A1(n711), .A2(n1021), .ZN(n694) );
  NAND2_X1 U759 ( .A1(n710), .A2(n694), .ZN(n700) );
  INV_X1 U760 ( .A(n1021), .ZN(n698) );
  NOR2_X1 U761 ( .A1(G1976), .A2(G288), .ZN(n1020) );
  NOR2_X1 U762 ( .A1(G1971), .A2(G303), .ZN(n695) );
  XOR2_X1 U763 ( .A(n695), .B(KEYINPUT105), .Z(n696) );
  NOR2_X1 U764 ( .A1(n1020), .A2(n696), .ZN(n697) );
  OR2_X1 U765 ( .A1(n698), .A2(n697), .ZN(n699) );
  AND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  INV_X1 U767 ( .A(n722), .ZN(n703) );
  NAND2_X1 U768 ( .A1(n702), .A2(n703), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n1020), .A2(n703), .ZN(n704) );
  NAND2_X1 U770 ( .A1(n704), .A2(KEYINPUT33), .ZN(n705) );
  NAND2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n707), .B(KEYINPUT106), .ZN(n709) );
  XNOR2_X1 U773 ( .A(G1981), .B(KEYINPUT107), .ZN(n708) );
  XNOR2_X1 U774 ( .A(n708), .B(G305), .ZN(n1013) );
  NAND2_X1 U775 ( .A1(n709), .A2(n1013), .ZN(n717) );
  NAND2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U777 ( .A1(G2090), .A2(G303), .ZN(n712) );
  NAND2_X1 U778 ( .A1(G8), .A2(n712), .ZN(n713) );
  NAND2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n722), .A2(n715), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U782 ( .A(n718), .B(KEYINPUT108), .ZN(n752) );
  NOR2_X1 U783 ( .A1(G1981), .A2(G305), .ZN(n719) );
  XOR2_X1 U784 ( .A(n719), .B(KEYINPUT24), .Z(n720) );
  XNOR2_X1 U785 ( .A(KEYINPUT98), .B(n720), .ZN(n721) );
  NOR2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n750) );
  NAND2_X1 U787 ( .A1(G105), .A2(n906), .ZN(n723) );
  XNOR2_X1 U788 ( .A(n723), .B(KEYINPUT96), .ZN(n724) );
  XNOR2_X1 U789 ( .A(n724), .B(KEYINPUT38), .ZN(n726) );
  NAND2_X1 U790 ( .A1(G117), .A2(n909), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n732) );
  NAND2_X1 U792 ( .A1(G129), .A2(n728), .ZN(n730) );
  NAND2_X1 U793 ( .A1(G141), .A2(n905), .ZN(n729) );
  NAND2_X1 U794 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U795 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U796 ( .A(KEYINPUT97), .B(n733), .Z(n901) );
  AND2_X1 U797 ( .A1(n934), .A2(n901), .ZN(n734) );
  XOR2_X1 U798 ( .A(KEYINPUT109), .B(n734), .Z(n961) );
  NOR2_X1 U799 ( .A1(G164), .A2(G1384), .ZN(n735) );
  NOR2_X1 U800 ( .A1(n523), .A2(n735), .ZN(n736) );
  XNOR2_X1 U801 ( .A(n736), .B(KEYINPUT92), .ZN(n775) );
  INV_X1 U802 ( .A(n775), .ZN(n764) );
  NAND2_X1 U803 ( .A1(G131), .A2(n905), .ZN(n738) );
  NAND2_X1 U804 ( .A1(G95), .A2(n906), .ZN(n737) );
  NAND2_X1 U805 ( .A1(n738), .A2(n737), .ZN(n742) );
  NAND2_X1 U806 ( .A1(G119), .A2(n728), .ZN(n740) );
  NAND2_X1 U807 ( .A1(G107), .A2(n909), .ZN(n739) );
  NAND2_X1 U808 ( .A1(n740), .A2(n739), .ZN(n741) );
  OR2_X1 U809 ( .A1(n742), .A2(n741), .ZN(n896) );
  AND2_X1 U810 ( .A1(n896), .A2(G1991), .ZN(n744) );
  NOR2_X1 U811 ( .A1(n934), .A2(n901), .ZN(n743) );
  NOR2_X1 U812 ( .A1(n744), .A2(n743), .ZN(n971) );
  NOR2_X1 U813 ( .A1(n764), .A2(n971), .ZN(n766) );
  NOR2_X1 U814 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n896), .ZN(n969) );
  NOR2_X1 U816 ( .A1(n745), .A2(n969), .ZN(n746) );
  NOR2_X1 U817 ( .A1(n766), .A2(n746), .ZN(n747) );
  NOR2_X1 U818 ( .A1(n961), .A2(n747), .ZN(n748) );
  XNOR2_X1 U819 ( .A(n748), .B(KEYINPUT39), .ZN(n749) );
  AND2_X1 U820 ( .A1(n749), .A2(n775), .ZN(n769) );
  OR2_X1 U821 ( .A1(n750), .A2(n769), .ZN(n751) );
  XOR2_X1 U822 ( .A(G2067), .B(KEYINPUT37), .Z(n774) );
  NAND2_X1 U823 ( .A1(n728), .A2(G128), .ZN(n753) );
  XNOR2_X1 U824 ( .A(n753), .B(KEYINPUT94), .ZN(n755) );
  NAND2_X1 U825 ( .A1(G116), .A2(n909), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U827 ( .A(n756), .B(KEYINPUT35), .ZN(n761) );
  NAND2_X1 U828 ( .A1(G140), .A2(n905), .ZN(n758) );
  NAND2_X1 U829 ( .A1(G104), .A2(n906), .ZN(n757) );
  NAND2_X1 U830 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U831 ( .A(KEYINPUT34), .B(n759), .Z(n760) );
  NAND2_X1 U832 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U833 ( .A(n762), .B(KEYINPUT36), .ZN(n918) );
  NAND2_X1 U834 ( .A1(n774), .A2(n918), .ZN(n965) );
  NOR2_X1 U835 ( .A1(n764), .A2(n965), .ZN(n763) );
  XNOR2_X1 U836 ( .A(n763), .B(KEYINPUT95), .ZN(n771) );
  XOR2_X1 U837 ( .A(G1986), .B(G290), .Z(n1028) );
  NOR2_X1 U838 ( .A1(n764), .A2(n1028), .ZN(n765) );
  XOR2_X1 U839 ( .A(KEYINPUT93), .B(n765), .Z(n767) );
  NOR2_X1 U840 ( .A1(n767), .A2(n766), .ZN(n768) );
  OR2_X1 U841 ( .A1(n769), .A2(n768), .ZN(n770) );
  AND2_X1 U842 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U843 ( .A1(n773), .A2(n772), .ZN(n777) );
  NOR2_X1 U844 ( .A1(n774), .A2(n918), .ZN(n963) );
  NAND2_X1 U845 ( .A1(n775), .A2(n963), .ZN(n776) );
  NAND2_X1 U846 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U847 ( .A(n778), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U848 ( .A(G2443), .B(G2446), .Z(n780) );
  XNOR2_X1 U849 ( .A(G2427), .B(G2451), .ZN(n779) );
  XNOR2_X1 U850 ( .A(n780), .B(n779), .ZN(n786) );
  XOR2_X1 U851 ( .A(G2430), .B(G2454), .Z(n782) );
  XNOR2_X1 U852 ( .A(G1341), .B(G1348), .ZN(n781) );
  XNOR2_X1 U853 ( .A(n782), .B(n781), .ZN(n784) );
  XOR2_X1 U854 ( .A(G2435), .B(G2438), .Z(n783) );
  XNOR2_X1 U855 ( .A(n784), .B(n783), .ZN(n785) );
  XOR2_X1 U856 ( .A(n786), .B(n785), .Z(n787) );
  AND2_X1 U857 ( .A1(G14), .A2(n787), .ZN(G401) );
  AND2_X1 U858 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U859 ( .A(G82), .ZN(G220) );
  INV_X1 U860 ( .A(G57), .ZN(G237) );
  NAND2_X1 U861 ( .A1(G7), .A2(G661), .ZN(n788) );
  XNOR2_X1 U862 ( .A(n788), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U863 ( .A(G223), .ZN(n853) );
  NAND2_X1 U864 ( .A1(n853), .A2(G567), .ZN(n789) );
  XOR2_X1 U865 ( .A(KEYINPUT11), .B(n789), .Z(G234) );
  INV_X1 U866 ( .A(G860), .ZN(n795) );
  OR2_X1 U867 ( .A1(n1010), .A2(n795), .ZN(G153) );
  INV_X1 U868 ( .A(G171), .ZN(G301) );
  INV_X1 U869 ( .A(n1008), .ZN(n798) );
  INV_X1 U870 ( .A(G868), .ZN(n833) );
  NAND2_X1 U871 ( .A1(n798), .A2(n833), .ZN(n790) );
  XNOR2_X1 U872 ( .A(n790), .B(KEYINPUT78), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G868), .A2(G301), .ZN(n791) );
  NAND2_X1 U874 ( .A1(n792), .A2(n791), .ZN(G284) );
  NOR2_X1 U875 ( .A1(G286), .A2(n833), .ZN(n794) );
  NOR2_X1 U876 ( .A1(G868), .A2(G299), .ZN(n793) );
  NOR2_X1 U877 ( .A1(n794), .A2(n793), .ZN(G297) );
  NAND2_X1 U878 ( .A1(n795), .A2(G559), .ZN(n796) );
  NAND2_X1 U879 ( .A1(n796), .A2(n1008), .ZN(n797) );
  XNOR2_X1 U880 ( .A(n797), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U881 ( .A1(n798), .A2(n833), .ZN(n799) );
  XNOR2_X1 U882 ( .A(n799), .B(KEYINPUT79), .ZN(n800) );
  NOR2_X1 U883 ( .A1(G559), .A2(n800), .ZN(n802) );
  NOR2_X1 U884 ( .A1(G868), .A2(n1010), .ZN(n801) );
  NOR2_X1 U885 ( .A1(n802), .A2(n801), .ZN(G282) );
  NAND2_X1 U886 ( .A1(G135), .A2(n905), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G111), .A2(n909), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U889 ( .A1(n728), .A2(G123), .ZN(n805) );
  XOR2_X1 U890 ( .A(KEYINPUT18), .B(n805), .Z(n806) );
  NOR2_X1 U891 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U892 ( .A1(n906), .A2(G99), .ZN(n808) );
  NAND2_X1 U893 ( .A1(n809), .A2(n808), .ZN(n966) );
  XNOR2_X1 U894 ( .A(G2096), .B(n966), .ZN(n810) );
  NOR2_X1 U895 ( .A1(G2100), .A2(n810), .ZN(n811) );
  XOR2_X1 U896 ( .A(KEYINPUT80), .B(n811), .Z(G156) );
  NAND2_X1 U897 ( .A1(n1008), .A2(G559), .ZN(n830) );
  XNOR2_X1 U898 ( .A(n1010), .B(n830), .ZN(n812) );
  NOR2_X1 U899 ( .A1(n812), .A2(G860), .ZN(n823) );
  NAND2_X1 U900 ( .A1(G67), .A2(n813), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G55), .A2(n814), .ZN(n815) );
  NAND2_X1 U902 ( .A1(n816), .A2(n815), .ZN(n822) );
  NAND2_X1 U903 ( .A1(G93), .A2(n817), .ZN(n820) );
  NAND2_X1 U904 ( .A1(G80), .A2(n818), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U906 ( .A1(n822), .A2(n821), .ZN(n832) );
  XNOR2_X1 U907 ( .A(n823), .B(n832), .ZN(G145) );
  XOR2_X1 U908 ( .A(KEYINPUT19), .B(n832), .Z(n824) );
  XNOR2_X1 U909 ( .A(G288), .B(n824), .ZN(n825) );
  XNOR2_X1 U910 ( .A(G166), .B(n825), .ZN(n828) );
  XNOR2_X1 U911 ( .A(n1023), .B(G290), .ZN(n826) );
  XNOR2_X1 U912 ( .A(n826), .B(G305), .ZN(n827) );
  XNOR2_X1 U913 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U914 ( .A(n829), .B(n1010), .ZN(n922) );
  XNOR2_X1 U915 ( .A(n830), .B(n922), .ZN(n831) );
  NAND2_X1 U916 ( .A1(n831), .A2(G868), .ZN(n835) );
  NAND2_X1 U917 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U918 ( .A1(n835), .A2(n834), .ZN(n836) );
  XOR2_X1 U919 ( .A(KEYINPUT86), .B(n836), .Z(G295) );
  NAND2_X1 U920 ( .A1(G2078), .A2(G2084), .ZN(n837) );
  XOR2_X1 U921 ( .A(KEYINPUT20), .B(n837), .Z(n838) );
  NAND2_X1 U922 ( .A1(G2090), .A2(n838), .ZN(n840) );
  XOR2_X1 U923 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n839) );
  XNOR2_X1 U924 ( .A(n840), .B(n839), .ZN(n841) );
  NAND2_X1 U925 ( .A1(G2072), .A2(n841), .ZN(G158) );
  XNOR2_X1 U926 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U927 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  NAND2_X1 U928 ( .A1(G120), .A2(G69), .ZN(n842) );
  NOR2_X1 U929 ( .A1(G237), .A2(n842), .ZN(n843) );
  XNOR2_X1 U930 ( .A(KEYINPUT90), .B(n843), .ZN(n844) );
  NAND2_X1 U931 ( .A1(n844), .A2(G108), .ZN(n858) );
  NAND2_X1 U932 ( .A1(n858), .A2(G567), .ZN(n851) );
  NOR2_X1 U933 ( .A1(G220), .A2(G219), .ZN(n845) );
  XOR2_X1 U934 ( .A(KEYINPUT88), .B(n845), .Z(n846) );
  XNOR2_X1 U935 ( .A(n846), .B(KEYINPUT22), .ZN(n847) );
  NOR2_X1 U936 ( .A1(G218), .A2(n847), .ZN(n848) );
  XOR2_X1 U937 ( .A(KEYINPUT89), .B(n848), .Z(n849) );
  NAND2_X1 U938 ( .A1(G96), .A2(n849), .ZN(n859) );
  NAND2_X1 U939 ( .A1(n859), .A2(G2106), .ZN(n850) );
  NAND2_X1 U940 ( .A1(n851), .A2(n850), .ZN(n860) );
  NAND2_X1 U941 ( .A1(G483), .A2(G661), .ZN(n852) );
  NOR2_X1 U942 ( .A1(n860), .A2(n852), .ZN(n855) );
  NAND2_X1 U943 ( .A1(n855), .A2(G36), .ZN(G176) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n853), .ZN(G217) );
  AND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n854) );
  NAND2_X1 U946 ( .A1(G661), .A2(n854), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G1), .A2(G3), .ZN(n856) );
  NAND2_X1 U948 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U949 ( .A(n857), .B(KEYINPUT110), .ZN(G188) );
  INV_X1 U951 ( .A(G120), .ZN(G236) );
  INV_X1 U952 ( .A(G108), .ZN(G238) );
  INV_X1 U953 ( .A(G96), .ZN(G221) );
  INV_X1 U954 ( .A(G69), .ZN(G235) );
  NOR2_X1 U955 ( .A1(n859), .A2(n858), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  INV_X1 U957 ( .A(n860), .ZN(G319) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2678), .Z(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2090), .Z(n864) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n863) );
  XNOR2_X1 U963 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U964 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U965 ( .A(G2096), .B(G2100), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n870) );
  XOR2_X1 U967 ( .A(G2078), .B(G2084), .Z(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(G227) );
  XOR2_X1 U969 ( .A(G1971), .B(G1956), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1986), .B(G1976), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n873), .B(G2474), .Z(n875) );
  XNOR2_X1 U973 ( .A(G1981), .B(G1966), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U975 ( .A(KEYINPUT41), .B(G1961), .Z(n877) );
  XNOR2_X1 U976 ( .A(G1996), .B(G1991), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U978 ( .A(n879), .B(n878), .ZN(G229) );
  NAND2_X1 U979 ( .A1(n728), .A2(G124), .ZN(n880) );
  XNOR2_X1 U980 ( .A(n880), .B(KEYINPUT44), .ZN(n882) );
  NAND2_X1 U981 ( .A1(G112), .A2(n909), .ZN(n881) );
  NAND2_X1 U982 ( .A1(n882), .A2(n881), .ZN(n886) );
  NAND2_X1 U983 ( .A1(G136), .A2(n905), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G100), .A2(n906), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U986 ( .A1(n886), .A2(n885), .ZN(G162) );
  NAND2_X1 U987 ( .A1(G130), .A2(n728), .ZN(n888) );
  NAND2_X1 U988 ( .A1(G118), .A2(n909), .ZN(n887) );
  NAND2_X1 U989 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U990 ( .A(KEYINPUT113), .B(n889), .Z(n894) );
  NAND2_X1 U991 ( .A1(G142), .A2(n905), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G106), .A2(n906), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(n892), .B(KEYINPUT45), .Z(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n895), .B(n966), .ZN(n900) );
  XOR2_X1 U997 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n898) );
  XOR2_X1 U998 ( .A(n896), .B(KEYINPUT114), .Z(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n903) );
  XNOR2_X1 U1001 ( .A(G164), .B(n901), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1003 ( .A(n904), .B(G162), .Z(n916) );
  NAND2_X1 U1004 ( .A1(G139), .A2(n905), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n906), .ZN(n907) );
  NAND2_X1 U1006 ( .A1(n908), .A2(n907), .ZN(n914) );
  NAND2_X1 U1007 ( .A1(G127), .A2(n728), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(G115), .A2(n909), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1010 ( .A(KEYINPUT47), .B(n912), .Z(n913) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n955) );
  XNOR2_X1 U1012 ( .A(G160), .B(n955), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1014 ( .A(n918), .B(n917), .Z(n919) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n919), .ZN(n920) );
  XOR2_X1 U1016 ( .A(KEYINPUT115), .B(n920), .Z(G395) );
  XNOR2_X1 U1017 ( .A(G171), .B(n1008), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(n921), .B(G286), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n924), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(KEYINPUT116), .B(n925), .ZN(G397) );
  NOR2_X1 U1022 ( .A1(G227), .A2(G229), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(KEYINPUT49), .B(n926), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G401), .A2(n927), .ZN(n928) );
  AND2_X1 U1025 ( .A1(G319), .A2(n928), .ZN(n930) );
  NOR2_X1 U1026 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1028 ( .A(G225), .ZN(G308) );
  INV_X1 U1029 ( .A(G29), .ZN(n952) );
  XOR2_X1 U1030 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n979) );
  XOR2_X1 U1031 ( .A(G2084), .B(G34), .Z(n931) );
  XNOR2_X1 U1032 ( .A(KEYINPUT54), .B(n931), .ZN(n948) );
  XNOR2_X1 U1033 ( .A(G2090), .B(G35), .ZN(n946) );
  XOR2_X1 U1034 ( .A(G2067), .B(G26), .Z(n932) );
  NAND2_X1 U1035 ( .A1(n932), .A2(G28), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(KEYINPUT119), .B(G2072), .ZN(n933) );
  XNOR2_X1 U1037 ( .A(n933), .B(G33), .ZN(n941) );
  XOR2_X1 U1038 ( .A(G1991), .B(G25), .Z(n936) );
  XNOR2_X1 U1039 ( .A(n934), .B(G32), .ZN(n935) );
  NAND2_X1 U1040 ( .A1(n936), .A2(n935), .ZN(n939) );
  XOR2_X1 U1041 ( .A(G27), .B(n937), .Z(n938) );
  NOR2_X1 U1042 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(n944), .ZN(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(n949), .B(KEYINPUT120), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(n979), .B(n950), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n953), .A2(G11), .ZN(n954) );
  XNOR2_X1 U1052 ( .A(n954), .B(KEYINPUT121), .ZN(n983) );
  XNOR2_X1 U1053 ( .A(G2072), .B(n955), .ZN(n958) );
  XOR2_X1 U1054 ( .A(G164), .B(G2078), .Z(n956) );
  XNOR2_X1 U1055 ( .A(KEYINPUT117), .B(n956), .ZN(n957) );
  NAND2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(n959), .B(KEYINPUT50), .ZN(n977) );
  XOR2_X1 U1058 ( .A(G2090), .B(G162), .Z(n960) );
  NOR2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1060 ( .A(KEYINPUT51), .B(n962), .Z(n975) );
  INV_X1 U1061 ( .A(n963), .ZN(n964) );
  NAND2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(G160), .B(G2084), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT52), .B(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(n981), .A2(G29), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n1039) );
  XNOR2_X1 U1074 ( .A(G20), .B(n984), .ZN(n988) );
  XNOR2_X1 U1075 ( .A(G1981), .B(G6), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(G1341), .B(G19), .ZN(n985) );
  NOR2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1079 ( .A(KEYINPUT59), .B(G1348), .Z(n989) );
  XNOR2_X1 U1080 ( .A(G4), .B(n989), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n992), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT60), .ZN(n997) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G21), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(G1961), .B(G5), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n1005) );
  XNOR2_X1 U1088 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(G1976), .B(G23), .Z(n1001) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1094 ( .A(n1003), .B(n1002), .Z(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(KEYINPUT61), .B(n1006), .Z(n1007) );
  NOR2_X1 U1097 ( .A1(G16), .A2(n1007), .ZN(n1036) );
  XOR2_X1 U1098 ( .A(G16), .B(KEYINPUT56), .Z(n1033) );
  XNOR2_X1 U1099 ( .A(G1348), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(n1009), .B(KEYINPUT122), .ZN(n1019) );
  XOR2_X1 U1101 ( .A(n1010), .B(G1341), .Z(n1012) );
  XNOR2_X1 U1102 ( .A(G166), .B(G1971), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G1966), .B(G168), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1106 ( .A(KEYINPUT57), .B(n1015), .Z(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1031) );
  INV_X1 U1109 ( .A(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1023), .B(G1956), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(G171), .B(G1961), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1116 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1117 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1118 ( .A(KEYINPUT123), .B(n1034), .Z(n1035) );
  NOR2_X1 U1119 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1120 ( .A(n1037), .B(KEYINPUT126), .Z(n1038) );
  NOR2_X1 U1121 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1040), .Z(n1041) );
  XNOR2_X1 U1123 ( .A(KEYINPUT127), .B(n1041), .ZN(G311) );
  INV_X1 U1124 ( .A(G311), .ZN(G150) );
endmodule

