

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  XNOR2_X1 U325 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U326 ( .A(n376), .B(n375), .ZN(n378) );
  INV_X1 U327 ( .A(G190GAT), .ZN(n464) );
  XOR2_X1 U328 ( .A(n460), .B(n441), .Z(n524) );
  XNOR2_X1 U329 ( .A(n464), .B(KEYINPUT58), .ZN(n465) );
  XNOR2_X1 U330 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT7), .B(KEYINPUT67), .Z(n294) );
  XNOR2_X1 U332 ( .A(G43GAT), .B(G29GAT), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U334 ( .A(KEYINPUT8), .B(n295), .Z(n412) );
  XOR2_X1 U335 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n297) );
  XNOR2_X1 U336 ( .A(KEYINPUT10), .B(KEYINPUT74), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n299) );
  INV_X1 U338 ( .A(KEYINPUT73), .ZN(n298) );
  XNOR2_X1 U339 ( .A(n299), .B(n298), .ZN(n301) );
  XOR2_X1 U340 ( .A(G50GAT), .B(G162GAT), .Z(n321) );
  XNOR2_X1 U341 ( .A(G134GAT), .B(n321), .ZN(n300) );
  XNOR2_X1 U342 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U343 ( .A(n412), .B(n302), .ZN(n313) );
  XOR2_X1 U344 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n304) );
  NAND2_X1 U345 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U347 ( .A(n305), .B(KEYINPUT77), .Z(n311) );
  XNOR2_X1 U348 ( .A(G92GAT), .B(G85GAT), .ZN(n307) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G106GAT), .ZN(n306) );
  XNOR2_X1 U350 ( .A(n307), .B(n306), .ZN(n361) );
  INV_X1 U351 ( .A(n361), .ZN(n359) );
  XOR2_X1 U352 ( .A(KEYINPUT76), .B(G218GAT), .Z(n309) );
  XNOR2_X1 U353 ( .A(G36GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n430) );
  XNOR2_X1 U355 ( .A(n359), .B(n430), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U357 ( .A(n313), .B(n312), .Z(n562) );
  XOR2_X1 U358 ( .A(n562), .B(KEYINPUT78), .Z(n549) );
  XOR2_X1 U359 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n315) );
  XNOR2_X1 U360 ( .A(KEYINPUT92), .B(KEYINPUT90), .ZN(n314) );
  XNOR2_X1 U361 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U362 ( .A(n316), .B(G106GAT), .Z(n318) );
  XOR2_X1 U363 ( .A(G148GAT), .B(G78GAT), .Z(n360) );
  XNOR2_X1 U364 ( .A(n360), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n320) );
  XNOR2_X1 U366 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n319), .B(KEYINPUT3), .ZN(n333) );
  XOR2_X1 U368 ( .A(n320), .B(n333), .Z(n323) );
  XOR2_X1 U369 ( .A(G141GAT), .B(G22GAT), .Z(n401) );
  XNOR2_X1 U370 ( .A(n401), .B(n321), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U372 ( .A(KEYINPUT22), .B(KEYINPUT93), .Z(n325) );
  NAND2_X1 U373 ( .A1(G228GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U375 ( .A(n327), .B(n326), .Z(n332) );
  XOR2_X1 U376 ( .A(KEYINPUT91), .B(G211GAT), .Z(n329) );
  XNOR2_X1 U377 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U379 ( .A(G197GAT), .B(n330), .Z(n438) );
  XNOR2_X1 U380 ( .A(n438), .B(KEYINPUT23), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n478) );
  XOR2_X1 U382 ( .A(G85GAT), .B(n333), .Z(n335) );
  XNOR2_X1 U383 ( .A(G29GAT), .B(G162GAT), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U385 ( .A(G141GAT), .B(n336), .ZN(n357) );
  XOR2_X1 U386 ( .A(KEYINPUT98), .B(KEYINPUT96), .Z(n338) );
  XNOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT97), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U389 ( .A(G148GAT), .B(G120GAT), .Z(n340) );
  XNOR2_X1 U390 ( .A(G1GAT), .B(G127GAT), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n355) );
  XOR2_X1 U393 ( .A(KEYINPUT5), .B(KEYINPUT99), .Z(n344) );
  XNOR2_X1 U394 ( .A(KEYINPUT94), .B(KEYINPUT4), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U396 ( .A(KEYINPUT95), .B(n345), .Z(n347) );
  NAND2_X1 U397 ( .A1(G225GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U399 ( .A(n348), .B(KEYINPUT6), .Z(n353) );
  XOR2_X1 U400 ( .A(KEYINPUT82), .B(G134GAT), .Z(n350) );
  XNOR2_X1 U401 ( .A(KEYINPUT83), .B(KEYINPUT0), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U403 ( .A(G113GAT), .B(n351), .ZN(n461) );
  XOR2_X1 U404 ( .A(n461), .B(KEYINPUT1), .Z(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U407 ( .A(n357), .B(n356), .Z(n477) );
  INV_X1 U408 ( .A(n477), .ZN(n534) );
  XNOR2_X1 U409 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n425) );
  INV_X1 U410 ( .A(n360), .ZN(n358) );
  NAND2_X1 U411 ( .A1(n359), .A2(n358), .ZN(n363) );
  NAND2_X1 U412 ( .A1(n361), .A2(n360), .ZN(n362) );
  NAND2_X1 U413 ( .A1(n363), .A2(n362), .ZN(n365) );
  NAND2_X1 U414 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U416 ( .A(G176GAT), .B(G64GAT), .Z(n432) );
  NAND2_X1 U417 ( .A1(n366), .A2(n432), .ZN(n370) );
  INV_X1 U418 ( .A(n366), .ZN(n368) );
  INV_X1 U419 ( .A(n432), .ZN(n367) );
  NAND2_X1 U420 ( .A1(n368), .A2(n367), .ZN(n369) );
  NAND2_X1 U421 ( .A1(n370), .A2(n369), .ZN(n376) );
  XOR2_X1 U422 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n372) );
  XNOR2_X1 U423 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n374) );
  XOR2_X1 U425 ( .A(G204GAT), .B(KEYINPUT32), .Z(n373) );
  XOR2_X1 U426 ( .A(G120GAT), .B(G71GAT), .Z(n453) );
  XOR2_X1 U427 ( .A(G57GAT), .B(KEYINPUT13), .Z(n384) );
  XOR2_X1 U428 ( .A(n453), .B(n384), .Z(n377) );
  XNOR2_X1 U429 ( .A(n378), .B(n377), .ZN(n583) );
  XNOR2_X1 U430 ( .A(KEYINPUT36), .B(n549), .ZN(n592) );
  XOR2_X1 U431 ( .A(G64GAT), .B(G71GAT), .Z(n380) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(G183GAT), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n396) );
  XOR2_X1 U434 ( .A(G15GAT), .B(G127GAT), .Z(n452) );
  XOR2_X1 U435 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n382) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n452), .B(n383), .ZN(n394) );
  XOR2_X1 U439 ( .A(n384), .B(G78GAT), .Z(n386) );
  XOR2_X1 U440 ( .A(G1GAT), .B(KEYINPUT68), .Z(n398) );
  XNOR2_X1 U441 ( .A(n398), .B(G155GAT), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U443 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n388) );
  XNOR2_X1 U444 ( .A(KEYINPUT80), .B(KEYINPUT12), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U446 ( .A(n390), .B(n389), .Z(n392) );
  XNOR2_X1 U447 ( .A(G22GAT), .B(G211GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U449 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U450 ( .A(n396), .B(n395), .Z(n587) );
  INV_X1 U451 ( .A(n587), .ZN(n574) );
  NOR2_X1 U452 ( .A1(n592), .A2(n574), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n397), .B(KEYINPUT45), .ZN(n413) );
  XOR2_X1 U454 ( .A(G169GAT), .B(G8GAT), .Z(n431) );
  XOR2_X1 U455 ( .A(n398), .B(n431), .Z(n400) );
  NAND2_X1 U456 ( .A1(G229GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U458 ( .A(n402), .B(n401), .Z(n410) );
  XOR2_X1 U459 ( .A(G15GAT), .B(G197GAT), .Z(n404) );
  XNOR2_X1 U460 ( .A(G50GAT), .B(G36GAT), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n406) );
  XNOR2_X1 U463 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U467 ( .A(n412), .B(n411), .Z(n509) );
  INV_X1 U468 ( .A(n509), .ZN(n578) );
  NAND2_X1 U469 ( .A1(n413), .A2(n578), .ZN(n414) );
  NOR2_X1 U470 ( .A1(n583), .A2(n414), .ZN(n415) );
  XOR2_X1 U471 ( .A(KEYINPUT114), .B(n415), .Z(n423) );
  XNOR2_X1 U472 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n583), .B(n416), .ZN(n570) );
  NOR2_X1 U474 ( .A1(n570), .A2(n578), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n417), .B(KEYINPUT46), .ZN(n418) );
  NOR2_X1 U476 ( .A1(n418), .A2(n587), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n419), .B(KEYINPUT113), .ZN(n420) );
  NOR2_X1 U478 ( .A1(n420), .A2(n562), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n421), .B(KEYINPUT47), .ZN(n422) );
  NAND2_X1 U480 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n536) );
  INV_X1 U482 ( .A(n536), .ZN(n442) );
  XNOR2_X1 U483 ( .A(KEYINPUT87), .B(KEYINPUT17), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n426), .B(G183GAT), .ZN(n427) );
  XOR2_X1 U485 ( .A(n427), .B(KEYINPUT86), .Z(n429) );
  XNOR2_X1 U486 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n460) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U490 ( .A(KEYINPUT79), .B(KEYINPUT100), .Z(n435) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U493 ( .A(n437), .B(n436), .Z(n440) );
  XNOR2_X1 U494 ( .A(n438), .B(G92GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  NAND2_X1 U496 ( .A1(n442), .A2(n524), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n443), .B(KEYINPUT54), .ZN(n444) );
  NOR2_X1 U498 ( .A1(n534), .A2(n444), .ZN(n577) );
  NAND2_X1 U499 ( .A1(n478), .A2(n577), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n445), .B(KEYINPUT55), .ZN(n463) );
  XOR2_X1 U501 ( .A(KEYINPUT20), .B(G190GAT), .Z(n447) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(G99GAT), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT84), .Z(n449) );
  XNOR2_X1 U505 ( .A(KEYINPUT85), .B(KEYINPUT88), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U507 ( .A(n451), .B(n450), .Z(n458) );
  XOR2_X1 U508 ( .A(n453), .B(n452), .Z(n455) );
  NAND2_X1 U509 ( .A1(G227GAT), .A2(G233GAT), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U511 ( .A(G169GAT), .B(n456), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U514 ( .A(n462), .B(n461), .ZN(n537) );
  NAND2_X1 U515 ( .A1(n463), .A2(n537), .ZN(n573) );
  NOR2_X1 U516 ( .A1(n549), .A2(n573), .ZN(n466) );
  XNOR2_X1 U517 ( .A(G1GAT), .B(KEYINPUT103), .ZN(n467) );
  XNOR2_X1 U518 ( .A(n467), .B(KEYINPUT102), .ZN(n468) );
  XOR2_X1 U519 ( .A(KEYINPUT34), .B(n468), .Z(n487) );
  NOR2_X1 U520 ( .A1(n578), .A2(n583), .ZN(n469) );
  XNOR2_X1 U521 ( .A(n469), .B(KEYINPUT71), .ZN(n498) );
  XNOR2_X1 U522 ( .A(KEYINPUT27), .B(KEYINPUT101), .ZN(n470) );
  XOR2_X1 U523 ( .A(n470), .B(n524), .Z(n533) );
  NOR2_X1 U524 ( .A1(n537), .A2(n478), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n471), .B(KEYINPUT26), .ZN(n576) );
  NAND2_X1 U526 ( .A1(n533), .A2(n576), .ZN(n475) );
  NAND2_X1 U527 ( .A1(n524), .A2(n537), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n478), .A2(n472), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n473), .Z(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U531 ( .A1(n477), .A2(n476), .ZN(n483) );
  XOR2_X1 U532 ( .A(n478), .B(KEYINPUT65), .Z(n479) );
  XOR2_X1 U533 ( .A(KEYINPUT28), .B(n479), .Z(n529) );
  INV_X1 U534 ( .A(n529), .ZN(n539) );
  NAND2_X1 U535 ( .A1(n539), .A2(n533), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n537), .A2(n480), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n534), .A2(n481), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n483), .A2(n482), .ZN(n495) );
  NAND2_X1 U539 ( .A1(n587), .A2(n549), .ZN(n484) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n484), .Z(n485) );
  NAND2_X1 U541 ( .A1(n495), .A2(n485), .ZN(n511) );
  NOR2_X1 U542 ( .A1(n498), .A2(n511), .ZN(n492) );
  NAND2_X1 U543 ( .A1(n492), .A2(n534), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n492), .A2(n524), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U548 ( .A1(n492), .A2(n537), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n491), .ZN(G1326GAT) );
  XOR2_X1 U551 ( .A(G22GAT), .B(KEYINPUT105), .Z(n494) );
  NAND2_X1 U552 ( .A1(n492), .A2(n529), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  NAND2_X1 U554 ( .A1(n495), .A2(n574), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n592), .A2(n496), .ZN(n497) );
  XNOR2_X1 U556 ( .A(KEYINPUT37), .B(n497), .ZN(n520) );
  NOR2_X1 U557 ( .A1(n520), .A2(n498), .ZN(n500) );
  XNOR2_X1 U558 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(n507) );
  NAND2_X1 U560 ( .A1(n507), .A2(n534), .ZN(n503) );
  XNOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n501), .B(KEYINPUT107), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n507), .A2(n524), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n537), .A2(n507), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U569 ( .A1(n529), .A2(n507), .ZN(n508) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(n508), .ZN(G1331GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n513) );
  NOR2_X1 U572 ( .A1(n509), .A2(n570), .ZN(n510) );
  XOR2_X1 U573 ( .A(KEYINPUT108), .B(n510), .Z(n521) );
  NOR2_X1 U574 ( .A1(n521), .A2(n511), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n517), .A2(n534), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NAND2_X1 U578 ( .A1(n517), .A2(n524), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U580 ( .A1(n537), .A2(n517), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U583 ( .A1(n517), .A2(n529), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n530) );
  NAND2_X1 U586 ( .A1(n530), .A2(n534), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  XOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT111), .Z(n526) );
  NAND2_X1 U590 ( .A1(n530), .A2(n524), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1337GAT) );
  NAND2_X1 U592 ( .A1(n537), .A2(n530), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT112), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  NAND2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n553) );
  NAND2_X1 U600 ( .A1(n553), .A2(n537), .ZN(n538) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(n538), .Z(n540) );
  NAND2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n548) );
  NOR2_X1 U603 ( .A1(n578), .A2(n548), .ZN(n541) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n541), .Z(G1340GAT) );
  NOR2_X1 U605 ( .A1(n548), .A2(n570), .ZN(n545) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n543) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT118), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U610 ( .A1(n574), .A2(n548), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n551) );
  XNOR2_X1 U614 ( .A(KEYINPUT51), .B(KEYINPUT119), .ZN(n550) );
  XNOR2_X1 U615 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n576), .ZN(n563) );
  NOR2_X1 U618 ( .A1(n578), .A2(n563), .ZN(n554) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  NOR2_X1 U620 ( .A1(n570), .A2(n563), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT52), .B(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U626 ( .A1(n574), .A2(n563), .ZN(n560) );
  XOR2_X1 U627 ( .A(KEYINPUT122), .B(n560), .Z(n561) );
  XNOR2_X1 U628 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  INV_X1 U629 ( .A(n562), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(G162GAT), .B(n565), .Z(G1347GAT) );
  NOR2_X1 U632 ( .A1(n578), .A2(n573), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT56), .Z(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n572) );
  NOR2_X1 U638 ( .A1(n570), .A2(n573), .ZN(n571) );
  XOR2_X1 U639 ( .A(n572), .B(n571), .Z(G1349GAT) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(G183GAT), .B(n575), .Z(G1350GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n591) );
  NOR2_X1 U643 ( .A1(n591), .A2(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U649 ( .A(n591), .ZN(n588) );
  NAND2_X1 U650 ( .A1(n588), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U653 ( .A(G211GAT), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1354GAT) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

