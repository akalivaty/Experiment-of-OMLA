//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G50), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G116), .ZN(new_n212));
  INV_X1    g0012(.A(G270), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n209), .B1(new_n210), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n208), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(G50), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT65), .Z(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n206), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g0033(.A1(new_n223), .A2(new_n224), .A3(new_n228), .A4(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  INV_X1    g0045(.A(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT68), .B(G50), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(G223), .A3(G1698), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n256), .B(new_n257), .C1(new_n216), .C2(new_n254), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  OAI211_X1 g0062(.A(G1), .B(G13), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G274), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OR2_X1    g0065(.A1(KEYINPUT69), .A2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(KEYINPUT69), .A2(G45), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  AND3_X1   g0068(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n205), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT70), .B1(new_n268), .B2(new_n205), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G226), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n260), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT71), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n260), .A2(new_n271), .A3(KEYINPUT71), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G190), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(G200), .A3(new_n279), .ZN(new_n282));
  INV_X1    g0082(.A(G13), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n283), .A2(new_n206), .A3(G1), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n210), .ZN(new_n285));
  OAI21_X1  g0085(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G150), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n206), .A2(G33), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n286), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n231), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n284), .A2(new_n293), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT72), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n205), .A2(G20), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT72), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n284), .B2(new_n293), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n285), .B(new_n294), .C1(new_n300), .C2(new_n210), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT9), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n281), .A2(new_n282), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n281), .A2(new_n305), .A3(new_n282), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n278), .A2(new_n308), .A3(new_n279), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n301), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(G179), .B1(new_n278), .B2(new_n279), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n309), .A2(KEYINPUT73), .A3(new_n301), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n312), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n307), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G68), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n246), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(G20), .B1(new_n320), .B2(new_n201), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n287), .A2(G159), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT82), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n261), .B2(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT82), .A3(G33), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n206), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G68), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n330), .B2(new_n206), .ZN(new_n334));
  OAI211_X1 g0134(.A(KEYINPUT16), .B(new_n324), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n331), .B1(new_n254), .B2(G20), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n328), .A2(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n327), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n319), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n336), .B1(new_n341), .B2(new_n323), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n335), .A2(new_n293), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n290), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n300), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n284), .B2(new_n344), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n273), .A2(new_n237), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT70), .ZN(new_n348));
  AND2_X1   g0148(.A1(KEYINPUT69), .A2(G45), .ZN(new_n349));
  NOR2_X1   g0149(.A1(KEYINPUT69), .A2(G45), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n349), .A2(new_n350), .A3(G41), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n351), .B2(G1), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n205), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n347), .B1(new_n354), .B2(new_n265), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G87), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n211), .A2(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G223), .B2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n357), .B1(new_n330), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT83), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT83), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n362), .B(new_n357), .C1(new_n330), .C2(new_n359), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n363), .A3(new_n259), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n355), .A2(new_n356), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(G200), .B1(new_n355), .B2(new_n364), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n343), .B(new_n346), .C1(new_n365), .C2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT17), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n343), .A2(new_n346), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n361), .A2(new_n259), .A3(new_n363), .ZN(new_n372));
  INV_X1    g0172(.A(new_n347), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n271), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n371), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n355), .A2(new_n364), .A3(new_n356), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT17), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n369), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(G169), .B1(new_n372), .B2(new_n374), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n355), .A2(new_n364), .A3(G179), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT18), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n343), .A2(new_n346), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n293), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n344), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n391), .A2(new_n289), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n389), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n295), .A2(G77), .A3(new_n297), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT75), .B1(new_n284), .B2(new_n216), .ZN(new_n395));
  AND3_X1   g0195(.A1(new_n284), .A2(KEYINPUT75), .A3(new_n216), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n254), .A2(G238), .A3(G1698), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n400), .C1(new_n218), .C2(new_n254), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(new_n259), .B1(G244), .B2(new_n274), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n271), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n398), .B1(new_n403), .B2(new_n308), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G179), .B2(new_n403), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(G200), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n406), .B(new_n398), .C1(new_n356), .C2(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  OR3_X1    g0208(.A1(new_n318), .A2(new_n388), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n274), .A2(G238), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n271), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n211), .A2(new_n255), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n237), .A2(G1698), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n327), .A2(new_n412), .A3(new_n338), .A4(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G97), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT76), .B1(new_n416), .B2(new_n259), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  AOI211_X1 g0218(.A(new_n418), .B(new_n263), .C1(new_n414), .C2(new_n415), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT13), .B1(new_n411), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n415), .ZN(new_n422));
  NOR2_X1   g0222(.A1(G226), .A2(G1698), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n237), .B2(G1698), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n422), .B1(new_n424), .B2(new_n254), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n418), .B1(new_n425), .B2(new_n263), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n416), .A2(KEYINPUT76), .A3(new_n259), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n271), .A4(new_n410), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n421), .A2(G179), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n421), .A2(KEYINPUT77), .A3(new_n430), .ZN(new_n433));
  INV_X1    g0233(.A(new_n411), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT77), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n429), .A4(new_n428), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(G169), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT14), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n433), .A2(KEYINPUT14), .A3(G169), .A4(new_n436), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n295), .A2(G68), .A3(new_n297), .ZN(new_n442));
  INV_X1    g0242(.A(new_n284), .ZN(new_n443));
  NOR3_X1   g0243(.A1(new_n443), .A2(KEYINPUT12), .A3(G68), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT12), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n284), .B2(new_n319), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n289), .A2(new_n216), .B1(new_n206), .B2(G68), .ZN(new_n450));
  INV_X1    g0250(.A(new_n287), .ZN(new_n451));
  OAI22_X1  g0251(.A1(new_n450), .A2(KEYINPUT78), .B1(new_n210), .B2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n450), .A2(KEYINPUT78), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n293), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT11), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(KEYINPUT11), .B(new_n293), .C1(new_n452), .C2(new_n453), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n442), .B(KEYINPUT79), .C1(new_n444), .C2(new_n446), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n449), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n441), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n430), .A2(G190), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n462), .B2(new_n421), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n433), .A2(G200), .A3(new_n436), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT80), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT80), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT81), .B1(new_n461), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT80), .ZN(new_n469));
  INV_X1    g0269(.A(new_n464), .ZN(new_n470));
  INV_X1    g0270(.A(new_n421), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n430), .A2(G190), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n469), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT80), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n477), .C1(new_n460), .C2(new_n441), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n409), .B1(new_n468), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n255), .A2(G244), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n330), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n263), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g0287(.A(KEYINPUT5), .B(G41), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n488), .A2(new_n263), .A3(G274), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n263), .ZN(new_n493));
  INV_X1    g0293(.A(G257), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n308), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n486), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n259), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(KEYINPUT84), .ZN(new_n499));
  INV_X1    g0299(.A(G179), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT84), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n501), .B(new_n491), .C1(new_n493), .C2(new_n494), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  INV_X1    g0304(.A(G97), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n504), .A2(new_n505), .A3(G107), .ZN(new_n506));
  XNOR2_X1  g0306(.A(G97), .B(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n508), .A2(new_n206), .B1(new_n216), .B2(new_n451), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n218), .B1(new_n337), .B2(new_n340), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n293), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n284), .A2(new_n505), .ZN(new_n512));
  AOI211_X1 g0312(.A(new_n293), .B(new_n284), .C1(new_n205), .C2(G33), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G97), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n496), .A2(new_n503), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT85), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT85), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n496), .A2(new_n503), .A3(new_n515), .A4(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n487), .A2(new_n495), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  INV_X1    g0323(.A(new_n515), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n521), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n517), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT86), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n517), .A2(new_n525), .A3(KEYINPUT86), .A4(new_n519), .ZN(new_n529));
  XNOR2_X1  g0329(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n261), .A2(new_n212), .A3(G20), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT23), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n206), .B2(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n218), .A2(KEYINPUT23), .A3(G20), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n206), .A2(G87), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n537), .B1(new_n339), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n326), .A2(new_n329), .A3(new_n206), .A4(new_n327), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n541), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n531), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .A3(new_n206), .A4(G87), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(new_n530), .A3(new_n539), .A4(new_n536), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n389), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n295), .B1(G1), .B2(new_n261), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT25), .B1(new_n284), .B2(new_n218), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n218), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n549), .A2(new_n218), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n493), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n494), .A2(G1698), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(G250), .B2(G1698), .ZN(new_n556));
  INV_X1    g0356(.A(G294), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n330), .A2(new_n556), .B1(new_n261), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n554), .A2(G264), .B1(new_n558), .B2(new_n259), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n491), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(G190), .ZN(new_n561));
  AOI21_X1  g0361(.A(G200), .B1(new_n559), .B2(new_n491), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n553), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n308), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n559), .A2(new_n500), .A3(new_n491), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n548), .C2(new_n552), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT19), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n542), .A2(new_n505), .A3(new_n218), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n415), .A2(new_n206), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n289), .A2(KEYINPUT19), .A3(new_n505), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(new_n541), .B2(new_n319), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n293), .B1(new_n284), .B2(new_n391), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n391), .B2(new_n549), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n217), .A2(G1698), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G238), .B2(G1698), .ZN(new_n577));
  OAI22_X1  g0377(.A1(new_n330), .A2(new_n577), .B1(new_n261), .B2(new_n212), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n259), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n265), .A2(new_n490), .ZN(new_n580));
  INV_X1    g0380(.A(G250), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n490), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n263), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n308), .ZN(new_n585));
  INV_X1    g0385(.A(new_n490), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n583), .B1(new_n264), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n259), .B2(new_n578), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n500), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n575), .A2(new_n585), .A3(new_n589), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n584), .A2(KEYINPUT87), .A3(new_n356), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT87), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n588), .B2(G190), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n513), .A2(G87), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n574), .B(new_n595), .C1(new_n588), .C2(new_n371), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n590), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n443), .A2(G116), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n600), .B1(new_n549), .B2(new_n212), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n292), .A2(new_n231), .B1(G20), .B2(new_n212), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n481), .B(new_n206), .C1(G33), .C2(new_n505), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(KEYINPUT20), .B(new_n602), .C1(new_n605), .C2(new_n606), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n601), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n219), .A2(G1698), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(G257), .B2(G1698), .ZN(new_n613));
  INV_X1    g0413(.A(G303), .ZN(new_n614));
  OAI22_X1  g0414(.A1(new_n330), .A2(new_n613), .B1(new_n614), .B2(new_n254), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n259), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n491), .B1(new_n493), .B2(new_n213), .ZN(new_n618));
  OAI21_X1  g0418(.A(G169), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n598), .B1(new_n611), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n599), .B1(new_n513), .B2(G116), .ZN(new_n621));
  INV_X1    g0421(.A(new_n610), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n603), .B(new_n604), .ZN(new_n623));
  AOI21_X1  g0423(.A(KEYINPUT20), .B1(new_n623), .B2(new_n602), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n621), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n616), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n625), .A2(KEYINPUT21), .A3(G169), .A4(new_n627), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n617), .A2(new_n618), .A3(new_n500), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(G190), .A3(new_n616), .ZN(new_n631));
  OAI21_X1  g0431(.A(G200), .B1(new_n617), .B2(new_n618), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n611), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n620), .A2(new_n628), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n567), .A2(new_n597), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n479), .A2(new_n528), .A3(new_n529), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT90), .Z(G372));
  AOI21_X1  g0437(.A(new_n597), .B1(new_n517), .B2(new_n519), .ZN(new_n638));
  XOR2_X1   g0438(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n597), .ZN(new_n641));
  INV_X1    g0441(.A(new_n516), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n638), .A2(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n591), .A2(new_n593), .ZN(new_n646));
  INV_X1    g0446(.A(new_n596), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n566), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n620), .A2(new_n628), .A3(new_n630), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n563), .B(new_n648), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n590), .B1(new_n651), .B2(new_n526), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n479), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n317), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n470), .A2(new_n473), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(new_n405), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n379), .B1(new_n461), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT92), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n385), .B2(new_n386), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n355), .A2(G179), .A3(new_n364), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n308), .B1(new_n355), .B2(new_n364), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(KEYINPUT18), .B1(new_n662), .B2(new_n370), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(KEYINPUT92), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n657), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n654), .B1(new_n667), .B2(new_n307), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n653), .A2(new_n668), .ZN(G369));
  NAND3_X1  g0469(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n611), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT93), .B1(new_n650), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n634), .B2(new_n677), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n650), .A2(KEYINPUT93), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G330), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n567), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n553), .B2(new_n676), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n566), .B2(new_n676), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n650), .A2(new_n676), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n688), .A2(new_n684), .B1(new_n649), .B2(new_n676), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n225), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n569), .A2(G116), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G1), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n229), .B2(new_n693), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT28), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n676), .B1(new_n645), .B2(new_n652), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT95), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT29), .ZN(new_n701));
  OAI211_X1 g0501(.A(KEYINPUT95), .B(new_n676), .C1(new_n645), .C2(new_n652), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n638), .A2(new_n640), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n643), .A2(new_n644), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI211_X1 g0506(.A(KEYINPUT29), .B(new_n676), .C1(new_n706), .C2(new_n652), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n635), .A2(new_n528), .A3(new_n529), .A4(new_n676), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n588), .A2(new_n559), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n520), .A3(KEYINPUT30), .A4(new_n629), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  INV_X1    g0511(.A(new_n495), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n498), .A2(new_n588), .A3(new_n559), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n626), .A2(G179), .A3(new_n616), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n711), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n588), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n522), .A2(new_n716), .A3(new_n627), .A4(new_n560), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n710), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(KEYINPUT31), .B1(new_n718), .B2(new_n675), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n718), .A2(new_n675), .ZN(new_n720));
  XOR2_X1   g0520(.A(KEYINPUT94), .B(KEYINPUT31), .Z(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n708), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n703), .A2(new_n707), .B1(G330), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n697), .B1(new_n725), .B2(G1), .ZN(G364));
  INV_X1    g0526(.A(new_n681), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n283), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n205), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n692), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n728), .A2(new_n683), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n727), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n691), .A2(new_n339), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT96), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(G355), .ZN(new_n742));
  AND2_X1   g0542(.A1(G355), .A2(new_n741), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n743), .B1(G116), .B2(new_n225), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n249), .A2(new_n489), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n691), .A2(new_n545), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n266), .A2(new_n267), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(new_n230), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n744), .B1(new_n745), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n231), .B1(G20), .B2(new_n308), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n736), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n732), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n206), .A2(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(new_n356), .A3(new_n371), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n254), .B1(new_n758), .B2(G329), .ZN(new_n759));
  INV_X1    g0559(.A(G283), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n206), .A2(new_n371), .A3(G179), .A4(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(G20), .A2(G179), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n356), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G326), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n766), .A2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(KEYINPUT33), .B(G317), .Z(new_n771));
  OAI21_X1  g0571(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n356), .A2(G179), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n206), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n756), .A2(G190), .A3(G200), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n774), .A2(new_n557), .B1(new_n775), .B2(new_n614), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n763), .A2(new_n772), .A3(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n779));
  AOI21_X1  g0579(.A(G200), .B1(new_n764), .B2(KEYINPUT97), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(new_n356), .A3(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G322), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n779), .A2(G190), .A3(new_n780), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n783), .A2(KEYINPUT98), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(KEYINPUT98), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n777), .B1(new_n778), .B2(new_n781), .C1(new_n782), .C2(new_n787), .ZN(new_n788));
  OR2_X1    g0588(.A1(new_n788), .A2(KEYINPUT99), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n758), .A2(KEYINPUT32), .A3(G159), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT32), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n791), .B1(new_n757), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n770), .A2(new_n319), .B1(new_n505), .B2(new_n774), .ZN(new_n795));
  INV_X1    g0595(.A(new_n767), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n796), .A2(new_n210), .B1(new_n775), .B2(new_n542), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n254), .B1(new_n762), .B2(new_n218), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n794), .A2(new_n795), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n799), .B1(new_n246), .B2(new_n787), .C1(new_n216), .C2(new_n781), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n788), .A2(KEYINPUT99), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n789), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n755), .B1(new_n802), .B2(new_n752), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n733), .B1(new_n739), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  INV_X1    g0605(.A(new_n732), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n407), .B1(new_n398), .B2(new_n676), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n405), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n405), .A2(new_n675), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n700), .A2(new_n702), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n810), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n676), .B(new_n812), .C1(new_n645), .C2(new_n652), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n724), .A2(G330), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n806), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n816), .A2(KEYINPUT101), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(KEYINPUT101), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n752), .A2(new_n734), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n806), .B1(new_n216), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n752), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n545), .B1(new_n822), .B2(new_n757), .ZN(new_n823));
  INV_X1    g0623(.A(new_n774), .ZN(new_n824));
  AOI22_X1  g0624(.A1(new_n824), .A2(G58), .B1(G68), .B2(new_n761), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n210), .B2(new_n775), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G137), .A2(new_n767), .B1(new_n769), .B2(G150), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n792), .B2(new_n781), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G143), .B2(new_n786), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n823), .B(new_n826), .C1(new_n829), .C2(KEYINPUT34), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n831));
  INV_X1    g0631(.A(new_n781), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(G116), .B1(new_n769), .B2(G283), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT100), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n339), .B1(new_n757), .B2(new_n778), .C1(new_n774), .C2(new_n505), .ZN(new_n836));
  INV_X1    g0636(.A(new_n775), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G107), .B1(new_n761), .B2(G87), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n614), .B2(new_n796), .ZN(new_n839));
  NOR3_X1   g0639(.A1(new_n835), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n786), .A2(G294), .B1(new_n833), .B2(new_n834), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n830), .A2(new_n831), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n820), .B1(new_n821), .B2(new_n842), .C1(new_n812), .C2(new_n735), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n818), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT102), .Z(G384));
  INV_X1    g0645(.A(new_n508), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT35), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n847), .A2(G116), .A3(new_n232), .A4(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT36), .Z(new_n850));
  OR3_X1    g0650(.A1(new_n229), .A2(new_n216), .A3(new_n320), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n210), .A2(G68), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n205), .B(G13), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n813), .A2(new_n809), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n439), .A2(new_n440), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n431), .C1(new_n465), .C2(new_n466), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n459), .A2(new_n675), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n858), .B1(new_n470), .B2(new_n473), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n460), .B2(new_n441), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n855), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n673), .B1(new_n343), .B2(new_n346), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n370), .B2(new_n377), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n382), .A2(new_n384), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n384), .B1(new_n376), .B2(new_n375), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n324), .B1(new_n333), .B2(new_n334), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n336), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n293), .A3(new_n335), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n346), .A2(new_n876), .B1(new_n380), .B2(new_n381), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n872), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n335), .A2(new_n293), .ZN(new_n879));
  INV_X1    g0679(.A(new_n334), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(G68), .A3(new_n332), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT16), .B1(new_n881), .B2(new_n324), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n346), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n382), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(KEYINPUT103), .A3(new_n367), .ZN(new_n885));
  INV_X1    g0685(.A(new_n673), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n878), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n871), .B1(new_n888), .B2(KEYINPUT37), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n887), .B1(new_n379), .B2(new_n387), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n866), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n887), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n388), .A2(new_n892), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n370), .A2(new_n377), .B1(new_n382), .B2(new_n883), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n892), .B1(new_n894), .B2(KEYINPUT103), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n869), .B1(new_n895), .B2(new_n878), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n893), .B(KEYINPUT38), .C1(new_n896), .C2(new_n871), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n865), .A2(new_n898), .B1(new_n666), .B2(new_n886), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n889), .A2(new_n890), .A3(new_n866), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n659), .A2(new_n379), .A3(new_n665), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n867), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n868), .A2(new_n658), .A3(KEYINPUT37), .A4(new_n870), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n384), .A2(new_n886), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n367), .A2(KEYINPUT92), .A3(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(KEYINPUT37), .A2(new_n906), .B1(new_n868), .B2(new_n870), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n902), .B2(new_n908), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n900), .A2(new_n909), .A3(KEYINPUT39), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n891), .B2(new_n897), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT104), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT104), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n907), .B(new_n904), .C1(new_n901), .C2(new_n867), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n897), .B(new_n911), .C1(new_n915), .C2(KEYINPUT38), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n914), .B(new_n916), .C1(new_n898), .C2(new_n911), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n461), .A2(new_n676), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n899), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n703), .A2(new_n479), .A3(new_n707), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n668), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n921), .B(new_n923), .Z(new_n924));
  AOI21_X1  g0724(.A(new_n722), .B1(new_n718), .B2(new_n675), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(KEYINPUT31), .B2(new_n720), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n708), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n858), .B1(new_n476), .B2(new_n441), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n856), .A2(new_n431), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n861), .B1(new_n929), .B2(new_n459), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n927), .B(new_n812), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n897), .B1(new_n915), .B2(KEYINPUT38), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n864), .A2(new_n935), .A3(new_n812), .A4(new_n927), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n891), .A2(new_n897), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n934), .A2(KEYINPUT40), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n479), .A2(new_n927), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n682), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n924), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n205), .B2(new_n729), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n924), .A2(new_n943), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n854), .B1(new_n945), .B2(new_n946), .ZN(G367));
  OAI221_X1 g0747(.A(new_n753), .B1(new_n225), .B2(new_n391), .C1(new_n747), .C2(new_n243), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n948), .A2(new_n732), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT105), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n574), .A2(new_n595), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n675), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n950), .B1(new_n597), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n641), .A2(KEYINPUT105), .A3(new_n952), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n590), .C2(new_n952), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G143), .A2(new_n767), .B1(new_n769), .B2(G159), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n246), .B2(new_n775), .C1(new_n216), .C2(new_n762), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n774), .A2(new_n319), .ZN(new_n959));
  INV_X1    g0759(.A(G137), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n254), .B1(new_n757), .B2(new_n960), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(G150), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n962), .B1(new_n210), .B2(new_n781), .C1(new_n963), .C2(new_n787), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G294), .A2(new_n769), .B1(new_n767), .B2(G311), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n761), .A2(G97), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(new_n218), .C2(new_n774), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G283), .B2(new_n832), .ZN(new_n968));
  INV_X1    g0768(.A(G317), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n775), .A2(new_n212), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n330), .B1(new_n969), .B2(new_n757), .C1(new_n970), .C2(KEYINPUT46), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(KEYINPUT46), .B2(new_n970), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n968), .B(new_n972), .C1(new_n614), .C2(new_n787), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n964), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT110), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT47), .Z(new_n976));
  OAI221_X1 g0776(.A(new_n949), .B1(new_n737), .B2(new_n956), .C1(new_n976), .C2(new_n821), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n524), .A2(new_n676), .ZN(new_n978));
  OR2_X1    g0778(.A1(new_n526), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n642), .A2(new_n675), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n689), .ZN(new_n982));
  XNOR2_X1  g0782(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n982), .B(new_n983), .Z(new_n984));
  INV_X1    g0784(.A(KEYINPUT109), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  OR3_X1    g0786(.A1(new_n981), .A2(new_n689), .A3(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n984), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n687), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n688), .A2(new_n684), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n686), .B2(new_n688), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(new_n683), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n725), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n725), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n692), .B(KEYINPUT41), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n731), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n981), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1001), .A2(new_n994), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT42), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1001), .A2(new_n566), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n517), .A2(new_n519), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n676), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n956), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(KEYINPUT43), .B2(new_n956), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1003), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n687), .A2(new_n1001), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1012), .C1(KEYINPUT107), .C2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(KEYINPUT107), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n977), .B1(new_n1000), .B2(new_n1016), .ZN(G387));
  OR2_X1    g0817(.A1(new_n240), .A2(new_n749), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n694), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1018), .A2(new_n746), .B1(new_n1019), .B2(new_n740), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1021));
  AND3_X1   g0821(.A1(new_n344), .A2(new_n210), .A3(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n694), .B(new_n489), .C1(new_n319), .C2(new_n216), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1021), .B1(new_n344), .B2(new_n210), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n218), .B2(new_n691), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n732), .B1(new_n1027), .B2(new_n754), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n686), .A2(new_n737), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n966), .B1(new_n391), .B2(new_n774), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n545), .B1(new_n963), .B2(new_n757), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n770), .A2(new_n290), .B1(new_n775), .B2(new_n216), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n796), .A2(new_n792), .ZN(new_n1033));
  NOR4_X1   g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n210), .B2(new_n787), .C1(new_n319), .C2(new_n781), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n545), .B1(G326), .B2(new_n758), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n774), .A2(new_n760), .B1(new_n775), .B2(new_n557), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G311), .A2(new_n769), .B1(new_n767), .B2(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1038), .B1(new_n614), .B2(new_n781), .C1(new_n787), .C2(new_n969), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT49), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1036), .B1(new_n212), .B2(new_n762), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1035), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1028), .B(new_n1029), .C1(new_n752), .C2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n996), .B2(new_n731), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n997), .A2(new_n692), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n725), .A2(new_n996), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT112), .ZN(G393));
  NAND2_X1  g0852(.A1(new_n993), .A2(new_n997), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n997), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n693), .B1(new_n992), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n753), .B1(new_n505), .B2(new_n225), .C1(new_n747), .C2(new_n252), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1057), .A2(new_n732), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n786), .A2(G159), .B1(G150), .B2(new_n767), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT51), .Z(new_n1060));
  AOI22_X1  g0860(.A1(new_n832), .A2(new_n344), .B1(new_n769), .B2(G50), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1061), .A2(KEYINPUT113), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(KEYINPUT113), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n824), .A2(G77), .B1(G87), .B2(new_n761), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n330), .B1(new_n758), .B2(G143), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1064), .B(new_n1065), .C1(new_n319), .C2(new_n775), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1062), .A2(new_n1063), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n786), .A2(G311), .B1(G317), .B2(new_n767), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI221_X1 g0869(.A(new_n339), .B1(new_n782), .B2(new_n757), .C1(new_n762), .C2(new_n218), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G303), .A2(new_n769), .B1(new_n837), .B2(G283), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n212), .B2(new_n774), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G294), .C2(new_n832), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1060), .A2(new_n1067), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1058), .B1(new_n821), .B2(new_n1074), .C1(new_n981), .C2(new_n737), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n993), .B2(new_n730), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1056), .A2(new_n1076), .ZN(G390));
  NAND2_X1  g0877(.A1(new_n865), .A2(new_n919), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n913), .A2(new_n917), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n676), .B(new_n808), .C1(new_n706), .C2(new_n652), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n809), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n864), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n919), .A3(new_n933), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1079), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n810), .B1(new_n860), .B2(new_n863), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(G330), .A3(new_n927), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n815), .A2(new_n810), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1089), .A2(KEYINPUT114), .A3(new_n864), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT114), .B1(new_n1089), .B2(new_n864), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n479), .A2(G330), .A3(new_n927), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n922), .A2(new_n1095), .A3(new_n668), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n864), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n927), .A2(G330), .A3(new_n812), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1081), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1086), .B1(new_n864), .B2(new_n1089), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n855), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1096), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1094), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1088), .A2(new_n1093), .A3(new_n1103), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n692), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1088), .A2(new_n731), .A3(new_n1093), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n819), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n732), .B1(new_n344), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n254), .B1(new_n757), .B2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n824), .A2(G159), .B1(new_n769), .B2(G137), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n210), .B2(new_n762), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(G128), .C2(new_n767), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n837), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT53), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n775), .B2(new_n963), .ZN(new_n1118));
  XOR2_X1   g0918(.A(KEYINPUT54), .B(G143), .Z(new_n1119));
  AOI22_X1  g0919(.A1(new_n1116), .A2(new_n1118), .B1(new_n832), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1115), .B(new_n1120), .C1(new_n822), .C2(new_n787), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n787), .A2(new_n212), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n339), .B1(new_n775), .B2(new_n542), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n796), .A2(new_n760), .B1(new_n216), .B2(new_n774), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1123), .B(new_n1124), .C1(G107), .C2(new_n769), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n762), .A2(new_n319), .B1(new_n757), .B2(new_n557), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1126), .A2(KEYINPUT115), .B1(G97), .B2(new_n832), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(KEYINPUT115), .C2(new_n1126), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1121), .B1(new_n1122), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1110), .B1(new_n1129), .B2(new_n752), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n918), .B2(new_n735), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1107), .A2(new_n1108), .A3(new_n1131), .ZN(G378));
  INV_X1    g0932(.A(new_n1096), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1106), .A2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g0934(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n301), .A2(new_n886), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT55), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n307), .A2(new_n317), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1138), .B1(new_n307), .B2(new_n317), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1138), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n318), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n1135), .A3(new_n1139), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n939), .B2(new_n682), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT119), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1140), .A2(new_n1141), .A3(new_n1136), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1135), .B1(new_n1144), .B2(new_n1139), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1142), .A2(new_n1145), .A3(KEYINPUT119), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n935), .B1(new_n932), .B2(new_n933), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n898), .A2(new_n936), .ZN(new_n1155));
  OAI211_X1 g0955(.A(G330), .B(new_n1153), .C1(new_n1154), .C2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n919), .B1(new_n913), .B2(new_n917), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1147), .B(new_n1156), .C1(new_n1157), .C2(new_n899), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n937), .A2(new_n938), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n900), .A2(new_n909), .ZN(new_n1160));
  OAI21_X1  g0960(.A(KEYINPUT40), .B1(new_n1160), .B2(new_n931), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n682), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1146), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n921), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1158), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1134), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n693), .B1(new_n1134), .B2(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1164), .A2(new_n921), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1164), .A2(new_n921), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n731), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n758), .C2(G124), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1175), .B1(new_n792), .B2(new_n762), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n824), .A2(G150), .B1(new_n769), .B2(G132), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n767), .A2(G125), .B1(new_n837), .B2(new_n1119), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n960), .C2(new_n781), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G128), .B2(new_n786), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT116), .Z(new_n1181));
  AOI21_X1  g0981(.A(new_n1176), .B1(new_n1181), .B2(KEYINPUT59), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(KEYINPUT59), .B2(new_n1181), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n767), .A2(G116), .B1(G58), .B2(new_n761), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1184), .B1(new_n505), .B2(new_n770), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n775), .A2(new_n216), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n330), .B(new_n262), .C1(new_n757), .C2(new_n760), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1185), .A2(new_n959), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n218), .B2(new_n787), .C1(new_n391), .C2(new_n781), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT58), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n545), .A2(G33), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G50), .B1(new_n1193), .B2(new_n262), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n821), .B1(new_n1183), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT117), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n806), .B(new_n1198), .C1(new_n210), .C2(new_n819), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1153), .A2(new_n734), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT120), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT120), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1203), .A3(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT121), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1174), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n730), .B1(new_n1158), .B2(new_n1165), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT121), .B1(new_n1209), .B2(new_n1205), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1169), .A2(new_n1171), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(G375));
  NAND3_X1  g1012(.A1(new_n1100), .A2(new_n1096), .A3(new_n1102), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT122), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n999), .A3(new_n1104), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n730), .B1(new_n1102), .B2(new_n1100), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1097), .A2(new_n734), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n732), .B1(G68), .B2(new_n1109), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n796), .A2(new_n822), .B1(new_n246), .B2(new_n762), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n330), .B(new_n1219), .C1(G128), .C2(new_n758), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n774), .A2(new_n210), .B1(new_n775), .B2(new_n792), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n769), .B2(new_n1119), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n963), .C2(new_n781), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n787), .A2(new_n960), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n787), .A2(new_n760), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n339), .B1(new_n614), .B2(new_n757), .C1(new_n762), .C2(new_n216), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n770), .A2(new_n212), .B1(new_n391), .B2(new_n774), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n796), .A2(new_n557), .B1(new_n775), .B2(new_n505), .ZN(new_n1228));
  NOR3_X1   g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n218), .B2(new_n781), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1223), .A2(new_n1224), .B1(new_n1225), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1218), .B1(new_n1231), .B2(new_n752), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1216), .B1(new_n1217), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1215), .A2(new_n1233), .ZN(G381));
  OR2_X1    g1034(.A1(G393), .A2(G396), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G384), .A2(new_n1235), .A3(G387), .A4(G390), .ZN(new_n1236));
  INV_X1    g1036(.A(G378), .ZN(new_n1237));
  INV_X1    g1037(.A(G381), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1211), .A4(new_n1238), .ZN(G407));
  NAND2_X1  g1039(.A1(new_n674), .A2(G213), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1211), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(G213), .A3(new_n1242), .ZN(G409));
  NOR2_X1   g1043(.A1(new_n1056), .A2(new_n1076), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G387), .B(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(G393), .B(G396), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT126), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(G387), .B2(new_n1244), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1245), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1246), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(G387), .B(G390), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1158), .A2(new_n1165), .A3(KEYINPUT124), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1255), .A2(new_n731), .A3(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(KEYINPUT125), .A3(new_n1201), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1106), .A2(new_n1133), .B1(new_n1165), .B2(new_n1158), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n999), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT125), .B1(new_n1257), .B2(new_n1201), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1237), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT123), .B1(new_n1211), .B2(G378), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1134), .A2(new_n1170), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(new_n692), .C1(KEYINPUT57), .C2(new_n1259), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1267));
  AND4_X1   g1067(.A1(KEYINPUT123), .A2(new_n1266), .A3(G378), .A4(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1263), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1240), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1214), .B1(new_n1271), .B2(new_n1103), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n692), .C1(new_n1271), .C2(new_n1213), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1233), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n844), .B(KEYINPUT102), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G384), .A2(new_n1273), .A3(new_n1233), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1241), .A2(G2897), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1270), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1277), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G384), .B1(new_n1233), .B2(new_n1273), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1269), .A2(new_n1285), .A3(new_n1240), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1253), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1266), .A2(new_n1267), .A3(G378), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT123), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1211), .A2(KEYINPUT123), .A3(G378), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1241), .B1(new_n1295), .B2(new_n1263), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT63), .B1(new_n1296), .B2(new_n1285), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1283), .A2(new_n1284), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1269), .A2(new_n1240), .A3(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1297), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT127), .B1(new_n1303), .B2(new_n1282), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1253), .B1(new_n1296), .B2(new_n1299), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1286), .A2(new_n1298), .ZN(new_n1306));
  AND4_X1   g1106(.A1(KEYINPUT127), .A2(new_n1282), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1290), .B1(new_n1304), .B2(new_n1307), .ZN(G405));
  OAI21_X1  g1108(.A(new_n1295), .B1(G378), .B2(new_n1211), .ZN(new_n1309));
  XOR2_X1   g1109(.A(new_n1309), .B(new_n1285), .Z(new_n1310));
  XNOR2_X1  g1110(.A(new_n1310), .B(new_n1301), .ZN(G402));
endmodule


