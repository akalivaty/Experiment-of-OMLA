//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G113), .B(G122), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT87), .B(G104), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(G237), .A2(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G214), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n195), .A2(KEYINPUT83), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n194), .B(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT18), .A2(G131), .ZN(new_n198));
  XNOR2_X1  g012(.A(new_n197), .B(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n200), .B(KEYINPUT75), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n200), .A2(new_n202), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n199), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT85), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT19), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n200), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT19), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n208), .B1(new_n213), .B2(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n197), .A2(new_n215), .A3(G131), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n197), .B2(G131), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n216), .A2(new_n217), .B1(G131), .B2(new_n197), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT73), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n219), .B1(new_n211), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n200), .A2(KEYINPUT73), .A3(KEYINPUT16), .ZN(new_n222));
  INV_X1    g036(.A(G125), .ZN(new_n223));
  OR2_X1    g037(.A1(new_n223), .A2(G140), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n221), .B(new_n222), .C1(KEYINPUT16), .C2(new_n224), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n225), .A2(new_n202), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n210), .A2(KEYINPUT85), .A3(new_n202), .A4(new_n212), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n214), .A2(new_n218), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT86), .B1(new_n207), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n207), .A2(new_n228), .A3(KEYINPUT86), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n192), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n216), .A2(new_n217), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT17), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(KEYINPUT17), .B2(new_n218), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n225), .B(new_n202), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n207), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(new_n191), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n187), .B(new_n188), .C1(new_n232), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT20), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n231), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n191), .B1(new_n242), .B2(new_n229), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n191), .B2(new_n237), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n244), .A2(KEYINPUT20), .A3(new_n187), .A4(new_n188), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n191), .A2(KEYINPUT88), .ZN(new_n246));
  AOI21_X1  g060(.A(G902), .B1(new_n237), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n246), .B2(new_n237), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G475), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n241), .A2(new_n245), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G478), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(KEYINPUT15), .ZN(new_n252));
  INV_X1    g066(.A(G116), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT14), .A3(G122), .ZN(new_n254));
  XNOR2_X1  g068(.A(G116), .B(G122), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(G107), .B(new_n254), .C1(new_n256), .C2(KEYINPUT14), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n195), .A2(G128), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G143), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT65), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n261), .A2(new_n266), .ZN(new_n269));
  OAI221_X1 g083(.A(new_n257), .B1(G107), .B2(new_n256), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n258), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n272), .A2(KEYINPUT90), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(KEYINPUT90), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n260), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n258), .A2(new_n271), .ZN(new_n276));
  OAI21_X1  g090(.A(G134), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n267), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n255), .B(G107), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT89), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n270), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  XOR2_X1   g095(.A(KEYINPUT9), .B(G234), .Z(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G217), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n283), .A2(new_n284), .A3(G953), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n281), .A2(new_n286), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n188), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n252), .B1(new_n289), .B2(KEYINPUT91), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT91), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  MUX2_X1   g106(.A(new_n252), .B(new_n290), .S(new_n292), .Z(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G952), .ZN(new_n295));
  NAND2_X1  g109(.A1(G234), .A2(G237), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT93), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT21), .B(G898), .Z(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(G902), .A3(G953), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n299), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT94), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n250), .A2(new_n293), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G469), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G140), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n294), .A2(G227), .ZN(new_n311));
  XOR2_X1   g125(.A(new_n310), .B(new_n311), .Z(new_n312));
  INV_X1    g126(.A(KEYINPUT11), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n264), .A2(G134), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n315));
  OAI21_X1  g129(.A(G137), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n262), .A2(G137), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n313), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT65), .B(G134), .ZN(new_n320));
  INV_X1    g134(.A(G137), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT11), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G131), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n321), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n313), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n317), .B1(new_n266), .B2(G137), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n325), .B(new_n326), .C1(new_n313), .C2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(KEYINPUT66), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n330), .B(G131), .C1(new_n319), .C2(new_n322), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G104), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n334), .B2(G107), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n336));
  INV_X1    g150(.A(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G104), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n335), .B(new_n338), .C1(G104), .C2(new_n337), .ZN(new_n339));
  XOR2_X1   g153(.A(KEYINPUT77), .B(G101), .Z(new_n340));
  OR2_X1    g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n337), .A2(G104), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n334), .A2(G107), .ZN(new_n343));
  OAI21_X1  g157(.A(G101), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n341), .A2(KEYINPUT10), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n202), .A2(G143), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT64), .B1(new_n195), .B2(G146), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n259), .B1(new_n347), .B2(KEYINPUT1), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT67), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT67), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n195), .A2(G146), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT64), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n202), .B2(G143), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n195), .A2(KEYINPUT64), .A3(G146), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n354), .B1(new_n359), .B2(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n195), .A2(G146), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n347), .A2(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(KEYINPUT1), .A3(new_n259), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n346), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g180(.A(KEYINPUT68), .B(new_n364), .C1(new_n353), .C2(new_n360), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n345), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(KEYINPUT78), .B(new_n345), .C1(new_n366), .C2(new_n367), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n339), .A2(G101), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n341), .A2(KEYINPUT4), .A3(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n363), .A2(new_n259), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT0), .B(G128), .Z(new_n376));
  AOI22_X1  g190(.A1(KEYINPUT0), .A2(new_n375), .B1(new_n350), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(new_n373), .A2(KEYINPUT4), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n341), .A2(new_n344), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n364), .B1(new_n363), .B2(new_n352), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n379), .B1(new_n382), .B2(KEYINPUT10), .ZN(new_n383));
  OAI211_X1 g197(.A(KEYINPUT79), .B(new_n333), .C1(new_n372), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n383), .B1(new_n370), .B2(new_n371), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n332), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n332), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n312), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n364), .B1(new_n353), .B2(new_n360), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n382), .B1(new_n391), .B2(new_n380), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(new_n332), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(KEYINPUT12), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n389), .A2(new_n312), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n309), .B(new_n188), .C1(new_n390), .C2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n396), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n388), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n312), .B1(new_n394), .B2(new_n389), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(G469), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n309), .A2(new_n188), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n398), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G221), .B1(new_n283), .B2(G902), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G214), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G119), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G116), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n253), .A2(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT2), .B(G113), .Z(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n415), .A2(KEYINPUT5), .ZN(new_n418));
  OAI21_X1  g232(.A(G113), .B1(new_n412), .B2(KEYINPUT5), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OR3_X1    g234(.A1(new_n420), .A2(new_n380), .A3(KEYINPUT80), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT80), .B1(new_n420), .B2(new_n380), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n415), .A2(new_n416), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n417), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n374), .A2(new_n424), .A3(new_n378), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n421), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(G110), .B(G122), .Z(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n421), .A2(new_n429), .A3(new_n425), .A4(new_n422), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n391), .A2(new_n223), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n223), .B2(new_n377), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n294), .A2(G224), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n433), .A2(new_n435), .ZN(new_n437));
  OR2_X1    g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n426), .A2(new_n439), .A3(new_n427), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n431), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  OAI22_X1  g255(.A1(new_n436), .A2(new_n437), .B1(KEYINPUT7), .B2(new_n435), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n418), .B(KEYINPUT81), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n417), .B1(new_n443), .B2(new_n419), .ZN(new_n444));
  INV_X1    g258(.A(new_n380), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n427), .B(KEYINPUT8), .Z(new_n447));
  OAI211_X1 g261(.A(new_n446), .B(new_n447), .C1(new_n445), .C2(new_n420), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT7), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n433), .A2(new_n449), .A3(new_n434), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n442), .A2(new_n448), .A3(new_n430), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n441), .A2(new_n451), .A3(new_n188), .ZN(new_n452));
  OAI21_X1  g266(.A(G210), .B1(G237), .B2(G902), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT82), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n454), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n441), .A2(new_n451), .A3(new_n188), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n410), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n308), .A2(new_n408), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n259), .A2(G119), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT23), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n411), .A2(G128), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(G110), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n461), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT24), .B(G110), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n236), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT74), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(G110), .B2(new_n466), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n226), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n470), .B1(new_n205), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT22), .B(G137), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n475), .B(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT25), .B1(new_n480), .B2(G902), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n284), .B1(G234), .B2(new_n188), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n475), .B(new_n478), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n188), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n483), .B(new_n188), .C1(new_n284), .C2(G234), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT72), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT32), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n324), .B1(G134), .B2(new_n321), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G131), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n328), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n366), .B2(new_n367), .ZN(new_n494));
  INV_X1    g308(.A(new_n424), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n329), .A2(new_n331), .A3(new_n377), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n391), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n495), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g314(.A(KEYINPUT70), .B(KEYINPUT28), .C1(new_n497), .C2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT70), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n497), .B2(KEYINPUT28), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n496), .A2(new_n499), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n424), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n501), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n193), .A2(G210), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n511), .B(G101), .Z(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n505), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n496), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n424), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n514), .A2(KEYINPUT69), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n507), .A3(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n518), .A2(KEYINPUT31), .A3(new_n507), .A4(new_n519), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n510), .A2(new_n514), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G472), .A2(G902), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n490), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n522), .A2(new_n523), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n501), .B(new_n514), .C1(new_n503), .C2(new_n508), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT32), .A3(new_n525), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT32), .B1(new_n531), .B2(new_n525), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT71), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G472), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n518), .A2(new_n514), .A3(new_n507), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n509), .B2(new_n514), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n497), .A2(new_n542), .ZN(new_n543));
  MUX2_X1   g357(.A(new_n497), .B(new_n543), .S(KEYINPUT28), .Z(new_n544));
  NOR2_X1   g358(.A1(new_n514), .A2(new_n540), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n537), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n489), .B1(new_n536), .B2(new_n548), .ZN(new_n549));
  AOI211_X1 g363(.A(KEYINPUT72), .B(new_n547), .C1(new_n533), .C2(new_n535), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n460), .B(new_n488), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n340), .ZN(G3));
  AND2_X1   g366(.A1(new_n406), .A2(new_n407), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n554));
  AOI21_X1  g368(.A(G902), .B1(new_n529), .B2(new_n530), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n537), .ZN(new_n556));
  OAI211_X1 g370(.A(KEYINPUT95), .B(G472), .C1(new_n524), .C2(G902), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n531), .A2(new_n525), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT96), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n553), .A2(new_n560), .A3(new_n561), .A4(new_n488), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n488), .A2(new_n558), .A3(new_n556), .A4(new_n557), .ZN(new_n563));
  OAI21_X1  g377(.A(KEYINPUT96), .B1(new_n563), .B2(new_n408), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n287), .A2(new_n288), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT33), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n281), .B2(KEYINPUT97), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n567), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n251), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n289), .A2(G478), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n251), .A2(new_n188), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n250), .A2(new_n458), .A3(new_n305), .A4(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n562), .A2(new_n564), .A3(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT34), .B(G104), .Z(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(G6));
  NAND4_X1  g393(.A1(new_n293), .A2(new_n249), .A3(new_n241), .A4(new_n245), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n580), .A2(new_n459), .A3(new_n306), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n562), .A2(new_n564), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT35), .B(G107), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G9));
  NOR2_X1   g398(.A1(new_n479), .A2(KEYINPUT36), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n475), .B(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(new_n188), .C1(new_n284), .C2(G234), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT98), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n486), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n460), .A2(new_n560), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G110), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT99), .B(KEYINPUT37), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G12));
  AOI211_X1 g409(.A(new_n528), .B(KEYINPUT32), .C1(new_n531), .C2(new_n525), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n490), .B(new_n526), .C1(new_n529), .C2(new_n530), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n534), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n596), .B1(new_n598), .B2(new_n528), .ZN(new_n599));
  OAI21_X1  g413(.A(KEYINPUT72), .B1(new_n599), .B2(new_n547), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n536), .A2(new_n489), .A3(new_n548), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n408), .A2(new_n459), .ZN(new_n603));
  INV_X1    g417(.A(G900), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n299), .B1(new_n604), .B2(new_n303), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n580), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n602), .A2(new_n603), .A3(new_n591), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G128), .ZN(G30));
  XOR2_X1   g422(.A(new_n605), .B(KEYINPUT39), .Z(new_n609));
  NAND2_X1  g423(.A1(new_n553), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n610), .B(KEYINPUT40), .Z(new_n611));
  NAND2_X1  g425(.A1(new_n455), .A2(new_n457), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT38), .Z(new_n613));
  NAND2_X1  g427(.A1(new_n250), .A2(new_n293), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n518), .A2(new_n507), .ZN(new_n616));
  INV_X1    g430(.A(new_n514), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n543), .A2(new_n514), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n618), .A2(new_n188), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(G472), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n536), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n591), .A2(new_n410), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n611), .A2(new_n615), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G143), .ZN(G45));
  INV_X1    g439(.A(new_n605), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n250), .A2(new_n574), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n602), .A2(new_n603), .A3(new_n591), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT100), .B(G146), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G48));
  OR2_X1    g444(.A1(new_n390), .A2(new_n397), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n188), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(G469), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n631), .B(new_n188), .C1(KEYINPUT101), .C2(new_n309), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n407), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n602), .A2(new_n488), .A3(new_n576), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT41), .B(G113), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G15));
  NAND4_X1  g455(.A1(new_n602), .A2(new_n488), .A3(new_n581), .A4(new_n638), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G116), .ZN(G18));
  NOR3_X1   g457(.A1(new_n636), .A2(new_n459), .A3(new_n637), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n602), .A2(new_n307), .A3(new_n591), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G119), .ZN(G21));
  NAND3_X1  g460(.A1(new_n250), .A2(new_n458), .A3(new_n293), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT102), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n555), .A2(new_n537), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n544), .A2(new_n617), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n526), .B1(new_n651), .B2(new_n529), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n653), .A2(new_n488), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n649), .A2(new_n638), .A3(new_n305), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT103), .B(G122), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G24));
  AND2_X1   g471(.A1(new_n653), .A2(new_n591), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n644), .A2(new_n627), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G125), .ZN(G27));
  OR2_X1    g474(.A1(new_n408), .A2(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n408), .A2(KEYINPUT104), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n612), .A2(new_n410), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n627), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n602), .A3(new_n488), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n598), .A2(new_n548), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n488), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n667), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n666), .A2(new_n667), .B1(new_n665), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n326), .ZN(G33));
  OAI211_X1 g486(.A(new_n488), .B(new_n663), .C1(new_n549), .C2(new_n550), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n661), .A2(new_n606), .A3(new_n662), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(G134), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G36));
  INV_X1    g491(.A(new_n398), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n396), .B1(new_n387), .B2(new_n384), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n679), .B1(new_n680), .B2(new_n401), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n400), .A2(KEYINPUT45), .A3(new_n402), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(G469), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT106), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n681), .A2(new_n682), .A3(new_n685), .A4(G469), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n405), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n678), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n689), .B(new_n404), .C1(new_n684), .C2(new_n686), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n407), .A3(new_n609), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n574), .A2(new_n241), .A3(new_n249), .A4(new_n245), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT43), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT43), .B1(new_n696), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(KEYINPUT44), .A3(new_n559), .A4(new_n591), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT108), .ZN(new_n702));
  INV_X1    g516(.A(new_n663), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(new_n559), .A3(new_n591), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n695), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G137), .ZN(G39));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n693), .A2(KEYINPUT109), .A3(new_n709), .A4(new_n407), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n404), .B1(new_n684), .B2(new_n686), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n398), .B1(new_n711), .B2(KEYINPUT46), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n709), .B(new_n407), .C1(new_n712), .C2(new_n691), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n627), .A2(new_n663), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n602), .A2(new_n488), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n407), .B1(new_n712), .B2(new_n691), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(KEYINPUT110), .A3(KEYINPUT47), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT110), .B1(new_n719), .B2(KEYINPUT47), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n716), .B(new_n718), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G140), .ZN(G42));
  AND2_X1   g538(.A1(new_n636), .A2(KEYINPUT49), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n636), .A2(KEYINPUT49), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n488), .A2(new_n409), .A3(new_n407), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n622), .ZN(new_n729));
  INV_X1    g543(.A(new_n696), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n613), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n648), .A2(new_n408), .ZN(new_n732));
  INV_X1    g546(.A(new_n591), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n626), .A4(new_n622), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n607), .A2(new_n628), .A3(new_n659), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n733), .B1(new_n600), .B2(new_n601), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(new_n603), .C1(new_n606), .C2(new_n627), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(KEYINPUT52), .A3(new_n659), .A4(new_n734), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n737), .A2(KEYINPUT114), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n408), .A2(new_n703), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n250), .A2(new_n293), .A3(new_n605), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n742), .B(new_n743), .C1(new_n549), .C2(new_n550), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n661), .A2(new_n664), .A3(new_n653), .A4(new_n662), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n591), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n673), .A2(new_n674), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n733), .B1(new_n744), .B2(new_n745), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT113), .B1(new_n751), .B2(new_n675), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n671), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n639), .A2(new_n642), .A3(new_n645), .A4(new_n655), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n575), .B(KEYINPUT111), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n562), .A2(new_n755), .A3(new_n564), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n551), .A2(new_n582), .A3(new_n756), .A4(new_n592), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n582), .A2(new_n592), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(KEYINPUT112), .A3(new_n551), .A4(new_n756), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n754), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n607), .A2(new_n628), .A3(new_n659), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT52), .A4(new_n734), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n741), .A2(new_n753), .A3(new_n762), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT53), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n737), .A2(new_n740), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n753), .A2(new_n768), .A3(new_n762), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT54), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n766), .A2(new_n769), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT115), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n753), .A2(new_n768), .A3(new_n762), .A4(KEYINPUT53), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT115), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n766), .A2(new_n775), .A3(new_n769), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n771), .B1(new_n777), .B2(KEYINPUT54), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n698), .A2(new_n699), .A3(new_n298), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n644), .A2(new_n654), .A3(new_n779), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n780), .B(KEYINPUT118), .Z(new_n781));
  AND2_X1   g595(.A1(new_n250), .A2(new_n574), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n636), .A2(new_n637), .A3(new_n703), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n488), .A3(new_n299), .A4(new_n729), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n781), .B(new_n295), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n638), .A2(new_n654), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n410), .A3(new_n613), .A4(new_n779), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT50), .Z(new_n789));
  NAND3_X1  g603(.A1(new_n784), .A2(new_n658), .A3(new_n779), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n785), .A2(new_n250), .A3(new_n574), .ZN(new_n791));
  AND4_X1   g605(.A1(KEYINPUT51), .A2(new_n789), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n716), .B1(new_n721), .B2(new_n722), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n793), .B(new_n794), .C1(new_n407), .C2(new_n636), .ZN(new_n795));
  INV_X1    g609(.A(new_n722), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n796), .A2(new_n720), .B1(new_n710), .B2(new_n715), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n636), .A2(new_n407), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT117), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n779), .A2(new_n654), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n703), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n786), .B1(new_n792), .B2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n804));
  INV_X1    g618(.A(new_n801), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n798), .B1(new_n793), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n797), .A2(KEYINPUT116), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n789), .A2(new_n790), .A3(new_n791), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n784), .A2(new_n779), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n669), .ZN(new_n813));
  XOR2_X1   g627(.A(new_n813), .B(KEYINPUT48), .Z(new_n814));
  AND3_X1   g628(.A1(new_n803), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n778), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(G952), .A2(G953), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n731), .B1(new_n816), .B2(new_n817), .ZN(G75));
  NAND2_X1  g632(.A1(new_n767), .A2(new_n770), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n188), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n454), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n431), .A2(new_n440), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n438), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT55), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n821), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n825), .B1(new_n821), .B2(new_n822), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n294), .A2(G952), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT119), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(G51));
  NAND3_X1  g644(.A1(new_n767), .A2(KEYINPUT54), .A3(new_n770), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n771), .ZN(new_n833));
  XOR2_X1   g647(.A(new_n404), .B(KEYINPUT57), .Z(new_n834));
  OAI21_X1  g648(.A(new_n631), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n820), .A2(new_n686), .A3(new_n684), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n828), .B1(new_n835), .B2(new_n836), .ZN(G54));
  NAND3_X1  g651(.A1(new_n820), .A2(KEYINPUT58), .A3(G475), .ZN(new_n838));
  INV_X1    g652(.A(new_n244), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n840), .A2(new_n841), .A3(new_n828), .ZN(G60));
  NAND2_X1  g656(.A1(new_n568), .A2(new_n569), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT120), .ZN(new_n844));
  XOR2_X1   g658(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n573), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n778), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n844), .A2(new_n846), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n819), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n850), .B1(new_n852), .B2(new_n831), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n848), .B1(new_n853), .B2(new_n829), .ZN(new_n854));
  INV_X1    g668(.A(new_n829), .ZN(new_n855));
  OAI211_X1 g669(.A(KEYINPUT122), .B(new_n855), .C1(new_n833), .C2(new_n850), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n847), .A2(new_n854), .A3(new_n856), .ZN(G63));
  INV_X1    g671(.A(new_n819), .ZN(new_n858));
  NAND2_X1  g672(.A1(G217), .A2(G902), .ZN(new_n859));
  XOR2_X1   g673(.A(new_n859), .B(KEYINPUT60), .Z(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n480), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n858), .A2(new_n586), .A3(new_n860), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n855), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n862), .A2(KEYINPUT61), .A3(new_n855), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(G66));
  AOI21_X1  g682(.A(new_n294), .B1(new_n300), .B2(G224), .ZN(new_n869));
  INV_X1    g683(.A(new_n762), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n869), .B1(new_n870), .B2(new_n294), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n823), .B1(G898), .B2(new_n294), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n871), .B(new_n872), .Z(G69));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n875));
  INV_X1    g689(.A(new_n624), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n739), .A2(new_n659), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n874), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n763), .A2(new_n624), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n673), .B1(new_n783), .B2(new_n580), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n553), .A3(new_n609), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n723), .A2(new_n707), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(G953), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n516), .A2(new_n517), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(new_n213), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT124), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n890));
  INV_X1    g704(.A(new_n888), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n723), .A2(new_n707), .A3(new_n884), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n878), .B2(new_n881), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n890), .B(new_n891), .C1(new_n893), .C2(G953), .ZN(new_n894));
  NAND2_X1  g708(.A1(G900), .A2(G953), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n671), .A2(new_n877), .A3(new_n675), .ZN(new_n896));
  OR3_X1    g710(.A1(new_n694), .A2(new_n648), .A3(new_n669), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n896), .A2(new_n707), .A3(new_n723), .A4(new_n897), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n888), .B(new_n895), .C1(new_n898), .C2(G953), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n889), .A2(new_n894), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT126), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n889), .A2(new_n894), .A3(new_n902), .A4(new_n899), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n889), .A2(new_n894), .A3(KEYINPUT125), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n901), .A2(new_n905), .A3(new_n906), .A4(new_n903), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(G72));
  NAND2_X1  g724(.A1(new_n893), .A2(new_n762), .ZN(new_n911));
  NAND2_X1  g725(.A1(G472), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT63), .Z(new_n913));
  AOI21_X1  g727(.A(new_n618), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n898), .B2(new_n870), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n538), .B(KEYINPUT127), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n777), .A2(new_n538), .A3(new_n618), .A4(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(new_n828), .ZN(G57));
endmodule


