//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT65), .Z(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(G325));
  XNOR2_X1  g033(.A(G325), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g034(.A(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n467), .A2(new_n469), .A3(G137), .A4(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n466), .A2(G2105), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n475), .A2(KEYINPUT69), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n471), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n479));
  NAND2_X1  g054(.A1(G113), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n470), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n478), .A2(new_n481), .ZN(G160));
  NAND2_X1  g057(.A1(new_n467), .A2(new_n469), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n470), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n486), .A2(KEYINPUT70), .A3(G136), .ZN(new_n492));
  AND4_X1   g067(.A1(new_n485), .A2(new_n489), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(KEYINPUT71), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  NAND4_X1  g072(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n470), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .ZN(new_n501));
  NAND2_X1  g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT3), .B(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G114), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n509), .A3(G2105), .ZN(new_n510));
  OAI21_X1  g085(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n500), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  XNOR2_X1  g090(.A(KEYINPUT6), .B(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G50), .A3(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT73), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(new_n516), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G88), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT5), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G62), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n518), .A2(new_n531), .ZN(G166));
  NAND3_X1  g107(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT74), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(KEYINPUT7), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n520), .A2(G89), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n537), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n519), .A2(new_n516), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n544), .A2(new_n545), .B1(new_n534), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  INV_X1    g127(.A(G43), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n544), .A2(new_n552), .B1(new_n534), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n549), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  NAND3_X1  g138(.A1(new_n516), .A2(G53), .A3(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n519), .A2(new_n516), .A3(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n568), .B2(new_n549), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n566), .A2(new_n569), .ZN(G299));
  OR2_X1    g145(.A1(new_n547), .A2(new_n550), .ZN(G301));
  OR2_X1    g146(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n572), .A2(new_n530), .A3(new_n521), .A4(new_n573), .ZN(G303));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n549), .B1(new_n527), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(G87), .B2(new_n520), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n534), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n534), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(KEYINPUT75), .A3(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT76), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n577), .A2(new_n585), .A3(new_n582), .A4(new_n580), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G288));
  AND3_X1   g162(.A1(new_n524), .A2(new_n526), .A3(G61), .ZN(new_n588));
  INV_X1    g163(.A(G73), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT77), .B1(new_n589), .B2(new_n523), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n591), .A2(G73), .A3(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n519), .A2(new_n516), .A3(G86), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n544), .A2(new_n598), .B1(new_n534), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n549), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n600), .A2(new_n602), .ZN(G290));
  XOR2_X1   g178(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n604));
  NAND3_X1  g179(.A1(new_n520), .A2(G92), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n581), .A2(G54), .ZN(new_n606));
  INV_X1    g181(.A(new_n604), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n544), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n527), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n605), .A2(new_n606), .A3(new_n609), .A4(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n615), .B2(G171), .ZN(G284));
  OAI21_X1  g192(.A(new_n616), .B1(new_n615), .B2(G171), .ZN(G321));
  NAND2_X1  g193(.A1(G299), .A2(new_n615), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G168), .B2(new_n615), .ZN(G280));
  XOR2_X1   g195(.A(G280), .B(KEYINPUT79), .Z(G297));
  INV_X1    g196(.A(new_n614), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  INV_X1    g199(.A(new_n557), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(new_n615), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n614), .A2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n504), .A2(new_n473), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n484), .A2(G123), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n486), .A2(G135), .ZN(new_n635));
  OR2_X1    g210(.A1(G99), .A2(G2105), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n636), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(G2096), .Z(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n639), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT15), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2435), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2435), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(KEYINPUT14), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2451), .B(G2454), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n648), .A2(new_n650), .ZN(new_n655));
  OR3_X1    g230(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n652), .B2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT80), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT81), .B(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n663), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n671));
  OAI221_X1 g246(.A(new_n667), .B1(new_n661), .B2(new_n670), .C1(new_n671), .C2(new_n668), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2096), .B(G2100), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT19), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT82), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n683), .B1(new_n681), .B2(new_n679), .C1(new_n687), .C2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n690), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT83), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NAND2_X1  g272(.A1(new_n484), .A2(G129), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n473), .A2(G105), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n486), .A2(G141), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT26), .Z(new_n702));
  NAND4_X1  g277(.A1(new_n698), .A2(new_n699), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(KEYINPUT90), .A3(G29), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT27), .B(G1996), .Z(new_n706));
  OAI21_X1  g281(.A(KEYINPUT90), .B1(G29), .B2(G32), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  AND3_X1   g284(.A1(new_n705), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n706), .B1(new_n705), .B2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n708), .A2(G33), .ZN(new_n713));
  NAND2_X1  g288(.A1(G115), .A2(G2104), .ZN(new_n714));
  INV_X1    g289(.A(G127), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n483), .B2(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n716), .A2(G2105), .B1(G139), .B2(new_n486), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n473), .A2(G103), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT25), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n713), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT89), .B(G2072), .Z(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n722), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n537), .A2(G16), .A3(new_n541), .ZN(new_n726));
  OR2_X1    g301(.A1(G16), .A2(G21), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT91), .B(G1966), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G171), .A2(G16), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G5), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1961), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT30), .B(G28), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n733), .A2(new_n734), .B1(new_n708), .B2(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n712), .A2(new_n725), .A3(new_n731), .A4(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT31), .B(G11), .Z(new_n738));
  NOR2_X1   g313(.A1(new_n733), .A2(new_n734), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n708), .A2(G27), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G164), .B2(new_n708), .ZN(new_n741));
  INV_X1    g316(.A(G2078), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  NOR4_X1   g319(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n728), .A2(new_n730), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT92), .ZN(new_n747));
  OR2_X1    g322(.A1(KEYINPUT24), .A2(G34), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT24), .A2(G34), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n748), .A2(new_n708), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G160), .B2(new_n708), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n638), .A2(new_n708), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n745), .A2(new_n747), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(KEYINPUT93), .ZN(new_n757));
  INV_X1    g332(.A(new_n732), .ZN(new_n758));
  NOR2_X1   g333(.A1(G5), .A2(G16), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n734), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n735), .A2(new_n708), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n729), .B1(new_n726), .B2(new_n727), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n764), .A2(new_n743), .A3(new_n725), .A4(new_n712), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n765), .A2(new_n754), .A3(new_n738), .A4(new_n739), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n766), .A2(new_n767), .A3(new_n747), .A4(new_n753), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n708), .B1(new_n494), .B2(new_n495), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n708), .A2(G35), .ZN(new_n770));
  OAI21_X1  g345(.A(KEYINPUT29), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n769), .A2(KEYINPUT29), .A3(new_n770), .ZN(new_n773));
  OAI21_X1  g348(.A(G2090), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G16), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n775), .A2(KEYINPUT23), .A3(G20), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT23), .ZN(new_n777));
  INV_X1    g352(.A(G20), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G16), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n566), .A2(new_n569), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n776), .B(new_n779), .C1(new_n780), .C2(new_n775), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT94), .Z(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G1956), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n784));
  INV_X1    g359(.A(G26), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G29), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n785), .A2(G29), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n484), .A2(G128), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n486), .A2(G140), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n470), .A2(G116), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n787), .B1(new_n792), .B2(G29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n786), .B1(new_n793), .B2(new_n784), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n782), .A2(G1956), .B1(G2067), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n774), .A2(new_n783), .A3(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n772), .A2(G2090), .A3(new_n773), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n757), .A2(new_n768), .A3(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G24), .B(G290), .S(G16), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1986), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n484), .A2(G119), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n486), .A2(G131), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n470), .A2(G107), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n802), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G25), .B(new_n806), .S(G29), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT35), .B(G1991), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  OR2_X1    g386(.A1(G16), .A2(G23), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n583), .B2(new_n775), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT33), .B(G1976), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G22), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT84), .B1(new_n816), .B2(G16), .ZN(new_n817));
  OR3_X1    g392(.A1(new_n816), .A2(KEYINPUT84), .A3(G16), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n817), .B(new_n818), .C1(G166), .C2(new_n775), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(G1971), .ZN(new_n820));
  INV_X1    g395(.A(G305), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G16), .ZN(new_n822));
  OR2_X1    g397(.A1(G6), .A2(G16), .ZN(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT32), .B(G1981), .ZN(new_n824));
  AND3_X1   g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n824), .B1(new_n822), .B2(new_n823), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n819), .A2(G1971), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n815), .A2(new_n820), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G1971), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n819), .B(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n833), .A2(KEYINPUT85), .A3(new_n815), .A4(new_n827), .ZN(new_n834));
  AOI211_X1 g409(.A(KEYINPUT86), .B(new_n811), .C1(new_n831), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n811), .A2(KEYINPUT86), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n811), .A2(KEYINPUT86), .ZN(new_n837));
  AND4_X1   g412(.A1(new_n834), .A2(new_n831), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n810), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT87), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n841), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n839), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n775), .A2(G19), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n557), .B2(new_n775), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(G1341), .Z(new_n848));
  OAI211_X1 g423(.A(new_n842), .B(new_n810), .C1(new_n835), .C2(new_n838), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n799), .A2(new_n845), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n794), .A2(G2067), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n622), .A2(G16), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(G4), .B2(G16), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT88), .B(G1348), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n850), .A2(new_n852), .A3(new_n857), .ZN(G311));
  INV_X1    g433(.A(new_n845), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n849), .A2(new_n768), .A3(new_n757), .A4(new_n798), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n861), .A2(new_n851), .A3(new_n856), .A4(new_n848), .ZN(G150));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n527), .B2(new_n864), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT95), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G651), .ZN(new_n867));
  XNOR2_X1  g442(.A(KEYINPUT96), .B(G55), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n581), .A2(new_n869), .B1(new_n520), .B2(G93), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT98), .B(G860), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NOR2_X1   g449(.A1(new_n614), .A2(new_n623), .ZN(new_n875));
  XNOR2_X1  g450(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT39), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n875), .B(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n867), .A2(new_n625), .A3(new_n870), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n865), .B(KEYINPUT95), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(new_n549), .ZN(new_n881));
  INV_X1    g456(.A(new_n870), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n557), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n878), .B(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n874), .B1(new_n885), .B2(new_n872), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT99), .ZN(G145));
  XNOR2_X1  g462(.A(new_n792), .B(G164), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n717), .A2(KEYINPUT100), .A3(new_n720), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n486), .A2(G142), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n484), .A2(G130), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(KEYINPUT101), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(KEYINPUT101), .ZN(new_n894));
  OR2_X1    g469(.A1(G106), .A2(G2105), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n895), .B(G2104), .C1(G118), .C2(new_n470), .ZN(new_n896));
  AND4_X1   g471(.A1(new_n891), .A2(new_n893), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n890), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n890), .A2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n631), .B(KEYINPUT102), .Z(new_n901));
  XNOR2_X1  g476(.A(new_n496), .B(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n904), .A2(new_n898), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(G160), .B(new_n638), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n806), .B(new_n703), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n907), .B(new_n908), .Z(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(G37), .ZN(new_n911));
  INV_X1    g486(.A(new_n909), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n903), .A2(new_n912), .A3(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g490(.A1(new_n871), .A2(new_n615), .ZN(new_n916));
  NAND2_X1  g491(.A1(G299), .A2(new_n614), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n622), .A2(new_n780), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n921), .A3(new_n918), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n924), .A3(KEYINPUT41), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n884), .B(new_n627), .Z(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g503(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(KEYINPUT105), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n929), .B(new_n930), .C1(new_n919), .C2(new_n927), .ZN(new_n931));
  XOR2_X1   g506(.A(G290), .B(new_n583), .Z(new_n932));
  XNOR2_X1  g507(.A(G303), .B(new_n821), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n932), .B(new_n933), .Z(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  XNOR2_X1  g510(.A(new_n931), .B(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n916), .B1(new_n936), .B2(new_n615), .ZN(G295));
  OAI21_X1  g512(.A(new_n916), .B1(new_n936), .B2(new_n615), .ZN(G331));
  NAND2_X1  g513(.A1(G286), .A2(G171), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n537), .A2(new_n541), .A3(G301), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n939), .A2(new_n879), .A3(new_n883), .A4(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n940), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n884), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n944), .A2(new_n884), .A3(KEYINPUT107), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n926), .ZN(new_n951));
  INV_X1    g526(.A(new_n934), .ZN(new_n952));
  INV_X1    g527(.A(new_n945), .ZN(new_n953));
  INV_X1    g528(.A(new_n941), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n954), .A3(new_n919), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n923), .A2(new_n925), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n943), .B2(new_n949), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n934), .B1(new_n959), .B2(new_n955), .ZN(new_n960));
  INV_X1    g535(.A(G37), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n953), .A2(new_n954), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n920), .A2(new_n922), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n950), .A2(new_n919), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n934), .ZN(new_n968));
  AND4_X1   g543(.A1(KEYINPUT43), .A2(new_n968), .A3(new_n911), .A4(new_n957), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT44), .B1(new_n964), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n968), .A2(new_n963), .A3(new_n957), .A4(new_n911), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(G397));
  OR2_X1    g551(.A1(new_n806), .A2(new_n808), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n514), .A2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT108), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n478), .A2(new_n982), .A3(new_n481), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n984), .A2(G1996), .A3(new_n703), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n984), .B(KEYINPUT109), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n792), .B(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1996), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n704), .ZN(new_n990));
  AOI211_X1 g565(.A(new_n977), .B(new_n985), .C1(new_n986), .C2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n792), .A2(G2067), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT125), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT125), .ZN(new_n994));
  INV_X1    g569(.A(new_n992), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n986), .A2(new_n990), .ZN(new_n996));
  INV_X1    g571(.A(new_n985), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n994), .B(new_n995), .C1(new_n998), .C2(new_n977), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n999), .A3(new_n986), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n806), .B(new_n808), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(new_n1001), .B2(new_n986), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n984), .A2(G1986), .A3(G290), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n988), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n986), .B1(new_n703), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n981), .A2(new_n989), .A3(new_n983), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT46), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1012));
  XNOR2_X1  g587(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1000), .A2(new_n1006), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(G166), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n1021));
  NAND4_X1  g596(.A1(G303), .A2(new_n1021), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n514), .B2(new_n978), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT69), .B1(new_n475), .B2(new_n476), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n473), .A2(new_n472), .A3(G101), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n486), .A2(G137), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n481), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(G40), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1025), .B1(new_n1027), .B2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n512), .A2(new_n510), .B1(new_n503), .B2(new_n504), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n1034), .B2(new_n500), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n983), .B(KEYINPUT115), .C1(new_n1035), .C2(new_n1026), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n514), .A2(new_n1026), .A3(new_n978), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1033), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n979), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n514), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n983), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n832), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1024), .B1(new_n1045), .B2(new_n1019), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1038), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n983), .B1(new_n1027), .B2(KEYINPUT110), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(G2090), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1044), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1023), .B(G8), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G1976), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n583), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n983), .A2(new_n1035), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(G8), .ZN(new_n1058));
  AOI211_X1 g633(.A(KEYINPUT112), .B(new_n1019), .C1(new_n983), .C2(new_n1035), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n594), .B2(KEYINPUT113), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT49), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n594), .A2(new_n1064), .A3(new_n595), .A4(new_n596), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1061), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1032), .B2(new_n979), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT112), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1057), .A2(new_n1056), .A3(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1060), .A2(KEYINPUT52), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1054), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(new_n1072), .A3(new_n1055), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1046), .A2(new_n1053), .A3(new_n1073), .A4(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1032), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1077));
  AOI211_X1 g652(.A(KEYINPUT50), .B(G1384), .C1(new_n1034), .C2(new_n500), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT110), .B1(new_n1078), .B2(new_n1027), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1079), .A3(new_n752), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1043), .A2(new_n730), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1077), .A2(new_n1079), .A3(KEYINPUT116), .A4(new_n752), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G286), .A2(new_n1019), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1015), .B1(new_n1076), .B2(new_n1087), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n1053), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1087), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(KEYINPUT117), .A4(new_n1046), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(G8), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n1094), .B2(new_n1024), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1089), .A2(new_n1090), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1976), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(new_n584), .A3(new_n586), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n821), .A2(new_n1062), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1099), .A2(new_n1100), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1102), .A2(new_n1053), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n1104));
  OR3_X1    g679(.A1(new_n1101), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1097), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1033), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1109));
  INV_X1    g684(.A(G1956), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g686(.A(KEYINPUT118), .B(new_n567), .C1(new_n568), .C2(new_n549), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1117));
  OAI21_X1  g692(.A(G299), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1117), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n780), .A3(new_n1115), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1040), .B(G1384), .C1(new_n1034), .C2(new_n500), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT45), .B1(new_n514), .B2(new_n978), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1032), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1111), .A2(new_n1121), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1348), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1057), .A2(G2067), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n614), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1111), .A2(new_n1126), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1121), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1133), .A2(KEYINPUT120), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT120), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n1140));
  AOI21_X1  g715(.A(G1348), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1141), .B2(new_n1130), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1130), .B1(new_n1143), .B2(new_n1128), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n614), .B1(new_n1144), .B2(KEYINPUT60), .ZN(new_n1145));
  NOR4_X1   g720(.A1(new_n1141), .A2(new_n1140), .A3(new_n622), .A4(new_n1130), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1041), .A2(new_n989), .A3(new_n983), .A4(new_n1042), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT121), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n989), .A4(new_n983), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  NAND2_X1  g728(.A1(new_n1057), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1149), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n557), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1155), .A2(new_n1158), .A3(new_n557), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1111), .A2(new_n1121), .A3(new_n1126), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1121), .B1(new_n1111), .B2(new_n1126), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1136), .A2(KEYINPUT61), .A3(new_n1127), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1147), .A2(new_n1160), .A3(new_n1164), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1139), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT51), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1082), .A2(G168), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1169), .B2(G8), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(G8), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1168), .B1(new_n1085), .B2(G286), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1171), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1124), .A2(new_n742), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT53), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT122), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1143), .A2(new_n734), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1178), .B(new_n1179), .C1(new_n1176), .C2(new_n1175), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G301), .B(KEYINPUT54), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1179), .B(KEYINPUT123), .Z(new_n1183));
  INV_X1    g758(.A(new_n1181), .ZN(new_n1184));
  OAI21_X1  g759(.A(G40), .B1(new_n478), .B2(KEYINPUT124), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n981), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n481), .B1(new_n478), .B2(KEYINPUT124), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1122), .A2(new_n1176), .A3(G2078), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1183), .A2(new_n1178), .A3(new_n1184), .A4(new_n1189), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1167), .A2(new_n1174), .A3(new_n1182), .A4(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1173), .A2(new_n1172), .ZN(new_n1192));
  OAI21_X1  g767(.A(KEYINPUT62), .B1(new_n1192), .B2(new_n1170), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1171), .B(new_n1194), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1193), .A2(new_n1195), .A3(G171), .A4(new_n1180), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1191), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1076), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1108), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  XOR2_X1   g774(.A(G290), .B(G1986), .Z(new_n1200));
  OAI21_X1  g775(.A(new_n1002), .B1(new_n984), .B2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1014), .B1(new_n1199), .B2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g777(.A1(new_n464), .A2(G227), .ZN(new_n1204));
  AND3_X1   g778(.A1(new_n914), .A2(new_n658), .A3(new_n1204), .ZN(new_n1205));
  AND3_X1   g779(.A1(new_n696), .A2(new_n1205), .A3(new_n973), .ZN(G308));
  NAND3_X1  g780(.A1(new_n696), .A2(new_n1205), .A3(new_n973), .ZN(G225));
endmodule


