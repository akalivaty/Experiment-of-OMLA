

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753;

  XNOR2_X1 U366 ( .A(n422), .B(G119), .ZN(n468) );
  XNOR2_X2 U367 ( .A(n731), .B(n491), .ZN(n617) );
  INV_X1 U368 ( .A(G953), .ZN(n744) );
  NOR2_X1 U369 ( .A1(n720), .A2(G953), .ZN(n721) );
  OR2_X1 U370 ( .A1(n572), .A2(n573), .ZN(n352) );
  XNOR2_X1 U371 ( .A(n611), .B(KEYINPUT122), .ZN(n612) );
  XNOR2_X1 U372 ( .A(n487), .B(n414), .ZN(n737) );
  XNOR2_X1 U373 ( .A(KEYINPUT16), .B(G122), .ZN(n478) );
  AND2_X1 U374 ( .A1(n751), .A2(n559), .ZN(n356) );
  NAND2_X1 U375 ( .A1(n532), .A2(n700), .ZN(n533) );
  XNOR2_X2 U376 ( .A(n481), .B(n480), .ZN(n731) );
  BUF_X1 U377 ( .A(n605), .Z(n672) );
  XNOR2_X1 U378 ( .A(G113), .B(KEYINPUT69), .ZN(n467) );
  XNOR2_X1 U379 ( .A(n404), .B(n380), .ZN(n677) );
  XNOR2_X1 U380 ( .A(n454), .B(KEYINPUT25), .ZN(n404) );
  NOR2_X1 U381 ( .A1(n723), .A2(G902), .ZN(n380) );
  NOR2_X1 U382 ( .A1(n659), .A2(n584), .ZN(n586) );
  NAND2_X1 U383 ( .A1(n560), .A2(n561), .ZN(n573) );
  INV_X1 U384 ( .A(KEYINPUT80), .ZN(n426) );
  XNOR2_X1 U385 ( .A(n419), .B(n418), .ZN(n510) );
  INV_X1 U386 ( .A(KEYINPUT8), .ZN(n418) );
  NAND2_X1 U387 ( .A1(n744), .A2(G234), .ZN(n419) );
  XNOR2_X1 U388 ( .A(n415), .B(G125), .ZN(n487) );
  INV_X1 U389 ( .A(G146), .ZN(n415) );
  XNOR2_X1 U390 ( .A(n411), .B(n412), .ZN(n703) );
  INV_X1 U391 ( .A(KEYINPUT100), .ZN(n412) );
  NOR2_X1 U392 ( .A1(n549), .A2(n548), .ZN(n411) );
  XNOR2_X1 U393 ( .A(n421), .B(n479), .ZN(n632) );
  XNOR2_X1 U394 ( .A(n473), .B(n472), .ZN(n421) );
  XNOR2_X1 U395 ( .A(n410), .B(KEYINPUT32), .ZN(n751) );
  NOR2_X1 U396 ( .A1(n477), .A2(n476), .ZN(n546) );
  NOR2_X1 U397 ( .A1(n570), .A2(n749), .ZN(n371) );
  NOR2_X1 U398 ( .A1(n588), .A2(n384), .ZN(n383) );
  XNOR2_X1 U399 ( .A(n424), .B(n423), .ZN(n605) );
  INV_X1 U400 ( .A(KEYINPUT45), .ZN(n423) );
  XNOR2_X1 U401 ( .A(G143), .B(G128), .ZN(n486) );
  XNOR2_X1 U402 ( .A(KEYINPUT65), .B(G131), .ZN(n506) );
  XNOR2_X1 U403 ( .A(G101), .B(G107), .ZN(n437) );
  XNOR2_X1 U404 ( .A(n547), .B(n494), .ZN(n701) );
  NAND2_X1 U405 ( .A1(n492), .A2(G214), .ZN(n700) );
  XNOR2_X1 U406 ( .A(n361), .B(n360), .ZN(n359) );
  INV_X1 U407 ( .A(KEYINPUT101), .ZN(n360) );
  NOR2_X1 U408 ( .A1(n703), .A2(n531), .ZN(n361) );
  NAND2_X1 U409 ( .A1(n396), .A2(n395), .ZN(n394) );
  AND2_X1 U410 ( .A1(n399), .A2(n398), .ZN(n397) );
  NAND2_X1 U411 ( .A1(n445), .A2(G902), .ZN(n398) );
  NAND2_X1 U412 ( .A1(n433), .A2(KEYINPUT0), .ZN(n432) );
  OR2_X2 U413 ( .A1(n585), .A2(n429), .ZN(n428) );
  NAND2_X1 U414 ( .A1(n345), .A2(n430), .ZN(n429) );
  INV_X1 U415 ( .A(KEYINPUT0), .ZN(n430) );
  XOR2_X1 U416 ( .A(KEYINPUT7), .B(G122), .Z(n514) );
  XNOR2_X1 U417 ( .A(n486), .B(G134), .ZN(n515) );
  NOR2_X1 U418 ( .A1(n715), .A2(n374), .ZN(n416) );
  NAND2_X1 U419 ( .A1(n389), .A2(n388), .ZN(n593) );
  NOR2_X1 U420 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X1 U421 ( .A1(n348), .A2(n397), .ZN(n388) );
  NOR2_X1 U422 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U423 ( .A(n413), .B(n509), .ZN(n549) );
  OR2_X1 U424 ( .A1(n632), .A2(G902), .ZN(n420) );
  NOR2_X1 U425 ( .A1(n562), .A2(n368), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n452), .B(n381), .ZN(n723) );
  XNOR2_X1 U427 ( .A(n451), .B(n737), .ZN(n381) );
  AND2_X1 U428 ( .A1(n407), .A2(n674), .ZN(n722) );
  AND2_X1 U429 ( .A1(n614), .A2(G953), .ZN(n725) );
  NOR2_X1 U430 ( .A1(n753), .A2(n581), .ZN(n582) );
  INV_X1 U431 ( .A(G237), .ZN(n474) );
  XNOR2_X1 U432 ( .A(n406), .B(n405), .ZN(n455) );
  XNOR2_X1 U433 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n405) );
  NAND2_X1 U434 ( .A1(n602), .A2(G234), .ZN(n406) );
  XNOR2_X1 U435 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n497) );
  XOR2_X1 U436 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n498) );
  XNOR2_X1 U437 ( .A(G113), .B(G143), .ZN(n503) );
  XOR2_X1 U438 ( .A(G122), .B(G104), .Z(n502) );
  XNOR2_X1 U439 ( .A(n435), .B(n515), .ZN(n473) );
  XNOR2_X1 U440 ( .A(KEYINPUT4), .B(G137), .ZN(n434) );
  NAND2_X1 U441 ( .A1(n347), .A2(n379), .ZN(n609) );
  INV_X1 U442 ( .A(n600), .ZN(n379) );
  XNOR2_X1 U443 ( .A(n453), .B(KEYINPUT15), .ZN(n602) );
  XNOR2_X1 U444 ( .A(G902), .B(KEYINPUT86), .ZN(n453) );
  XNOR2_X1 U445 ( .A(KEYINPUT83), .B(KEYINPUT76), .ZN(n482) );
  XOR2_X1 U446 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n483) );
  NAND2_X1 U447 ( .A1(G234), .A2(G237), .ZN(n458) );
  INV_X1 U448 ( .A(n683), .ZN(n685) );
  INV_X1 U449 ( .A(KEYINPUT1), .ZN(n392) );
  NOR2_X1 U450 ( .A1(n397), .A2(n392), .ZN(n390) );
  NAND2_X1 U451 ( .A1(n378), .A2(n606), .ZN(n740) );
  INV_X1 U452 ( .A(n609), .ZN(n378) );
  XNOR2_X1 U453 ( .A(G140), .B(KEYINPUT10), .ZN(n414) );
  XNOR2_X1 U454 ( .A(KEYINPUT87), .B(G110), .ZN(n438) );
  XNOR2_X1 U455 ( .A(G104), .B(KEYINPUT73), .ZN(n436) );
  XNOR2_X1 U456 ( .A(n473), .B(n387), .ZN(n738) );
  INV_X1 U457 ( .A(KEYINPUT92), .ZN(n387) );
  XNOR2_X1 U458 ( .A(n576), .B(n385), .ZN(n716) );
  XNOR2_X1 U459 ( .A(KEYINPUT41), .B(KEYINPUT106), .ZN(n385) );
  NOR2_X2 U460 ( .A1(n373), .A2(n372), .ZN(n538) );
  INV_X1 U461 ( .A(n431), .ZN(n372) );
  NAND2_X1 U462 ( .A1(n677), .A2(n678), .ZN(n683) );
  XNOR2_X1 U463 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U464 ( .A(n516), .B(n515), .ZN(n517) );
  AND2_X1 U465 ( .A1(n674), .A2(G475), .ZN(n400) );
  XOR2_X1 U466 ( .A(KEYINPUT59), .B(n625), .Z(n626) );
  XNOR2_X1 U467 ( .A(n617), .B(n619), .ZN(n620) );
  INV_X1 U468 ( .A(KEYINPUT35), .ZN(n375) );
  NAND2_X1 U469 ( .A1(n376), .A2(n349), .ZN(n659) );
  XNOR2_X1 U470 ( .A(n377), .B(KEYINPUT28), .ZN(n376) );
  AND2_X1 U471 ( .A1(n577), .A2(n680), .ZN(n377) );
  XNOR2_X1 U472 ( .A(n417), .B(KEYINPUT104), .ZN(n551) );
  NAND2_X1 U473 ( .A1(n546), .A2(n528), .ZN(n417) );
  AND2_X1 U474 ( .A1(n367), .A2(n366), .ZN(n365) );
  NAND2_X1 U475 ( .A1(n364), .A2(n363), .ZN(n362) );
  XNOR2_X1 U476 ( .A(n724), .B(n723), .ZN(n386) );
  INV_X1 U477 ( .A(G125), .ZN(n669) );
  OR2_X1 U478 ( .A1(n537), .A2(n536), .ZN(n345) );
  AND2_X1 U479 ( .A1(n353), .A2(n556), .ZN(n346) );
  XOR2_X1 U480 ( .A(n599), .B(n598), .Z(n347) );
  AND2_X1 U481 ( .A1(n393), .A2(n392), .ZN(n348) );
  XOR2_X1 U482 ( .A(n578), .B(KEYINPUT105), .Z(n349) );
  AND2_X1 U483 ( .A1(G214), .A2(n499), .ZN(n350) );
  NOR2_X1 U484 ( .A1(n707), .A2(n715), .ZN(n351) );
  AND2_X1 U485 ( .A1(n593), .A2(n558), .ZN(n353) );
  INV_X1 U486 ( .A(n528), .ZN(n547) );
  AND2_X1 U487 ( .A1(n492), .A2(G210), .ZN(n354) );
  INV_X1 U488 ( .A(G902), .ZN(n395) );
  AND2_X1 U489 ( .A1(n578), .A2(n522), .ZN(n355) );
  NAND2_X1 U490 ( .A1(n365), .A2(n362), .ZN(n749) );
  NAND2_X1 U491 ( .A1(n542), .A2(n541), .ZN(n559) );
  NAND2_X1 U492 ( .A1(n356), .A2(n560), .ZN(n370) );
  XNOR2_X2 U493 ( .A(n357), .B(n375), .ZN(n560) );
  NAND2_X1 U494 ( .A1(n752), .A2(n559), .ZN(n572) );
  NAND2_X1 U495 ( .A1(n358), .A2(n555), .ZN(n357) );
  XNOR2_X1 U496 ( .A(n416), .B(KEYINPUT34), .ZN(n358) );
  NAND2_X1 U497 ( .A1(n428), .A2(n359), .ZN(n373) );
  XNOR2_X2 U498 ( .A(n590), .B(KEYINPUT19), .ZN(n585) );
  XNOR2_X2 U499 ( .A(n533), .B(KEYINPUT81), .ZN(n590) );
  INV_X1 U500 ( .A(n563), .ZN(n364) );
  NAND2_X1 U501 ( .A1(n562), .A2(n368), .ZN(n366) );
  NAND2_X1 U502 ( .A1(n563), .A2(n368), .ZN(n367) );
  INV_X1 U503 ( .A(KEYINPUT102), .ZN(n368) );
  NAND2_X1 U504 ( .A1(n369), .A2(n371), .ZN(n571) );
  NAND2_X1 U505 ( .A1(n370), .A2(KEYINPUT44), .ZN(n369) );
  NAND2_X1 U506 ( .A1(n431), .A2(n428), .ZN(n374) );
  NOR2_X1 U507 ( .A1(n374), .A2(n692), .ZN(n565) );
  NOR2_X1 U508 ( .A1(n374), .A2(n568), .ZN(n650) );
  XNOR2_X1 U509 ( .A(n560), .B(G122), .ZN(G24) );
  NAND2_X1 U510 ( .A1(n382), .A2(n670), .ZN(n595) );
  XNOR2_X1 U511 ( .A(n383), .B(n589), .ZN(n382) );
  XNOR2_X1 U512 ( .A(n587), .B(KEYINPUT47), .ZN(n384) );
  NAND2_X1 U513 ( .A1(n585), .A2(KEYINPUT0), .ZN(n427) );
  XNOR2_X1 U514 ( .A(n571), .B(n426), .ZN(n425) );
  NAND2_X1 U515 ( .A1(n425), .A2(n352), .ZN(n424) );
  NAND2_X2 U516 ( .A1(n726), .A2(n610), .ZN(n674) );
  NAND2_X2 U517 ( .A1(n408), .A2(n604), .ZN(n407) );
  NAND2_X1 U518 ( .A1(n400), .A2(n407), .ZN(n627) );
  NOR2_X1 U519 ( .A1(n386), .A2(n725), .ZN(G66) );
  NAND2_X1 U520 ( .A1(n397), .A2(n393), .ZN(n578) );
  NAND2_X1 U521 ( .A1(n552), .A2(n593), .ZN(n554) );
  OR2_X1 U522 ( .A1(n642), .A2(n394), .ZN(n393) );
  INV_X1 U523 ( .A(n445), .ZN(n396) );
  NAND2_X1 U524 ( .A1(n642), .A2(n445), .ZN(n399) );
  NAND2_X1 U525 ( .A1(n407), .A2(n401), .ZN(n613) );
  AND2_X1 U526 ( .A1(n674), .A2(G478), .ZN(n401) );
  NAND2_X1 U527 ( .A1(n407), .A2(n402), .ZN(n621) );
  AND2_X1 U528 ( .A1(n674), .A2(G210), .ZN(n402) );
  NAND2_X1 U529 ( .A1(n407), .A2(n403), .ZN(n634) );
  AND2_X1 U530 ( .A1(n674), .A2(G472), .ZN(n403) );
  NAND2_X1 U531 ( .A1(n409), .A2(n601), .ZN(n408) );
  XNOR2_X1 U532 ( .A(n575), .B(n574), .ZN(n409) );
  NAND2_X1 U533 ( .A1(n557), .A2(n346), .ZN(n410) );
  XNOR2_X2 U534 ( .A(n538), .B(KEYINPUT22), .ZN(n557) );
  NAND2_X1 U535 ( .A1(n625), .A2(n395), .ZN(n413) );
  NAND2_X1 U536 ( .A1(n685), .A2(n355), .ZN(n466) );
  XNOR2_X2 U537 ( .A(n420), .B(G472), .ZN(n680) );
  XNOR2_X2 U538 ( .A(G116), .B(KEYINPUT3), .ZN(n422) );
  NOR2_X2 U539 ( .A1(n605), .A2(n602), .ZN(n575) );
  NAND2_X1 U540 ( .A1(n557), .A2(n556), .ZN(n563) );
  AND2_X2 U541 ( .A1(n427), .A2(n432), .ZN(n431) );
  INV_X1 U542 ( .A(n345), .ZN(n433) );
  INV_X1 U543 ( .A(KEYINPUT71), .ZN(n589) );
  INV_X1 U544 ( .A(KEYINPUT79), .ZN(n574) );
  XNOR2_X1 U545 ( .A(n500), .B(n350), .ZN(n501) );
  XNOR2_X1 U546 ( .A(n518), .B(n517), .ZN(n611) );
  INV_X1 U547 ( .A(n749), .ZN(n750) );
  XNOR2_X1 U548 ( .A(n506), .B(n434), .ZN(n435) );
  XNOR2_X1 U549 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U550 ( .A(n439), .B(n438), .ZN(n480) );
  NAND2_X1 U551 ( .A1(n744), .A2(G227), .ZN(n440) );
  XNOR2_X1 U552 ( .A(n440), .B(G140), .ZN(n442) );
  XNOR2_X1 U553 ( .A(G146), .B(KEYINPUT75), .ZN(n441) );
  XNOR2_X1 U554 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U555 ( .A(n480), .B(n443), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n738), .B(n444), .ZN(n642) );
  XNOR2_X1 U557 ( .A(KEYINPUT68), .B(G469), .ZN(n445) );
  XNOR2_X1 U558 ( .A(G128), .B(G110), .ZN(n446) );
  XNOR2_X1 U559 ( .A(n446), .B(KEYINPUT93), .ZN(n450) );
  XOR2_X1 U560 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n448) );
  XNOR2_X1 U561 ( .A(G119), .B(G137), .ZN(n447) );
  XNOR2_X1 U562 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U563 ( .A(n450), .B(n449), .Z(n452) );
  NAND2_X1 U564 ( .A1(G221), .A2(n510), .ZN(n451) );
  NAND2_X1 U565 ( .A1(G217), .A2(n455), .ZN(n454) );
  NAND2_X1 U566 ( .A1(n455), .A2(G221), .ZN(n457) );
  INV_X1 U567 ( .A(KEYINPUT21), .ZN(n456) );
  XNOR2_X1 U568 ( .A(n457), .B(n456), .ZN(n678) );
  XNOR2_X1 U569 ( .A(n458), .B(KEYINPUT88), .ZN(n459) );
  XNOR2_X1 U570 ( .A(KEYINPUT14), .B(n459), .ZN(n461) );
  NAND2_X1 U571 ( .A1(n461), .A2(G952), .ZN(n460) );
  XOR2_X1 U572 ( .A(KEYINPUT89), .B(n460), .Z(n712) );
  NOR2_X1 U573 ( .A1(n712), .A2(G953), .ZN(n537) );
  INV_X1 U574 ( .A(n537), .ZN(n465) );
  NAND2_X1 U575 ( .A1(n461), .A2(G902), .ZN(n462) );
  XOR2_X1 U576 ( .A(KEYINPUT90), .B(n462), .Z(n534) );
  NAND2_X1 U577 ( .A1(G953), .A2(n534), .ZN(n463) );
  OR2_X1 U578 ( .A1(n463), .A2(G900), .ZN(n464) );
  NAND2_X1 U579 ( .A1(n465), .A2(n464), .ZN(n522) );
  XNOR2_X1 U580 ( .A(n466), .B(KEYINPUT74), .ZN(n477) );
  XNOR2_X2 U581 ( .A(n468), .B(n467), .ZN(n479) );
  NOR2_X1 U582 ( .A1(G953), .A2(G237), .ZN(n499) );
  NAND2_X1 U583 ( .A1(n499), .A2(G210), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n469), .B(G146), .ZN(n471) );
  XNOR2_X1 U585 ( .A(G101), .B(KEYINPUT5), .ZN(n470) );
  XNOR2_X1 U586 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U587 ( .A1(n395), .A2(n474), .ZN(n492) );
  NAND2_X1 U588 ( .A1(n680), .A2(n700), .ZN(n475) );
  XNOR2_X1 U589 ( .A(n475), .B(KEYINPUT30), .ZN(n476) );
  XNOR2_X2 U590 ( .A(n479), .B(n478), .ZN(n481) );
  XNOR2_X1 U591 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U592 ( .A(KEYINPUT4), .B(n484), .Z(n490) );
  NAND2_X1 U593 ( .A1(G224), .A2(n744), .ZN(n485) );
  XNOR2_X1 U594 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U595 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U596 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U597 ( .A1(n617), .A2(n602), .ZN(n493) );
  XNOR2_X2 U598 ( .A(n493), .B(n354), .ZN(n532) );
  BUF_X1 U599 ( .A(n532), .Z(n528) );
  XNOR2_X1 U600 ( .A(KEYINPUT72), .B(KEYINPUT38), .ZN(n494) );
  NAND2_X1 U601 ( .A1(n546), .A2(n701), .ZN(n496) );
  XOR2_X1 U602 ( .A(KEYINPUT70), .B(KEYINPUT39), .Z(n495) );
  XNOR2_X1 U603 ( .A(n496), .B(n495), .ZN(n544) );
  INV_X1 U604 ( .A(n544), .ZN(n520) );
  XNOR2_X1 U605 ( .A(n498), .B(n497), .ZN(n500) );
  XNOR2_X1 U606 ( .A(n737), .B(n501), .ZN(n508) );
  XNOR2_X1 U607 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U608 ( .A(KEYINPUT98), .B(n504), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n508), .B(n507), .ZN(n625) );
  XOR2_X1 U611 ( .A(KEYINPUT13), .B(G475), .Z(n509) );
  XOR2_X1 U612 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n512) );
  NAND2_X1 U613 ( .A1(G217), .A2(n510), .ZN(n511) );
  XNOR2_X1 U614 ( .A(n512), .B(n511), .ZN(n518) );
  XNOR2_X1 U615 ( .A(G116), .B(G107), .ZN(n513) );
  XNOR2_X1 U616 ( .A(n514), .B(n513), .ZN(n516) );
  NAND2_X1 U617 ( .A1(n611), .A2(n395), .ZN(n519) );
  XNOR2_X1 U618 ( .A(n519), .B(G478), .ZN(n548) );
  INV_X1 U619 ( .A(n548), .ZN(n521) );
  OR2_X1 U620 ( .A1(n549), .A2(n521), .ZN(n653) );
  INV_X1 U621 ( .A(n653), .ZN(n666) );
  NAND2_X1 U622 ( .A1(n520), .A2(n666), .ZN(n606) );
  XNOR2_X1 U623 ( .A(n606), .B(G134), .ZN(G36) );
  XOR2_X1 U624 ( .A(G140), .B(KEYINPUT113), .Z(n530) );
  XNOR2_X1 U625 ( .A(KEYINPUT103), .B(KEYINPUT43), .ZN(n527) );
  AND2_X1 U626 ( .A1(n549), .A2(n521), .ZN(n664) );
  INV_X1 U627 ( .A(n677), .ZN(n558) );
  NAND2_X1 U628 ( .A1(n522), .A2(n558), .ZN(n523) );
  INV_X1 U629 ( .A(n678), .ZN(n531) );
  NOR2_X1 U630 ( .A1(n523), .A2(n531), .ZN(n577) );
  NAND2_X1 U631 ( .A1(n664), .A2(n577), .ZN(n524) );
  XNOR2_X1 U632 ( .A(n680), .B(KEYINPUT6), .ZN(n556) );
  NOR2_X1 U633 ( .A1(n524), .A2(n556), .ZN(n591) );
  NAND2_X1 U634 ( .A1(n591), .A2(n700), .ZN(n525) );
  NOR2_X1 U635 ( .A1(n525), .A2(n593), .ZN(n526) );
  XOR2_X1 U636 ( .A(n527), .B(n526), .Z(n529) );
  NOR2_X1 U637 ( .A1(n529), .A2(n528), .ZN(n600) );
  XOR2_X1 U638 ( .A(n530), .B(n600), .Z(G42) );
  NOR2_X1 U639 ( .A1(G898), .A2(n744), .ZN(n732) );
  NAND2_X1 U640 ( .A1(n732), .A2(n534), .ZN(n535) );
  XNOR2_X1 U641 ( .A(n535), .B(KEYINPUT91), .ZN(n536) );
  BUF_X1 U642 ( .A(n557), .Z(n542) );
  INV_X1 U643 ( .A(n680), .ZN(n539) );
  NAND2_X1 U644 ( .A1(n558), .A2(n539), .ZN(n540) );
  NOR2_X1 U645 ( .A1(n593), .A2(n540), .ZN(n541) );
  XNOR2_X1 U646 ( .A(G110), .B(KEYINPUT110), .ZN(n543) );
  XNOR2_X1 U647 ( .A(n559), .B(n543), .ZN(G12) );
  INV_X1 U648 ( .A(n664), .ZN(n658) );
  NOR2_X1 U649 ( .A1(n544), .A2(n658), .ZN(n545) );
  XNOR2_X1 U650 ( .A(n545), .B(KEYINPUT40), .ZN(n581) );
  XOR2_X1 U651 ( .A(G131), .B(n581), .Z(G33) );
  AND2_X1 U652 ( .A1(n549), .A2(n548), .ZN(n555) );
  INV_X1 U653 ( .A(n555), .ZN(n550) );
  NOR2_X1 U654 ( .A1(n551), .A2(n550), .ZN(n588) );
  XOR2_X1 U655 ( .A(G143), .B(n588), .Z(G45) );
  NOR2_X1 U656 ( .A1(n556), .A2(n683), .ZN(n552) );
  INV_X1 U657 ( .A(KEYINPUT33), .ZN(n553) );
  XNOR2_X1 U658 ( .A(n554), .B(n553), .ZN(n715) );
  INV_X1 U659 ( .A(KEYINPUT44), .ZN(n561) );
  INV_X1 U660 ( .A(n593), .ZN(n687) );
  NAND2_X1 U661 ( .A1(n687), .A2(n677), .ZN(n562) );
  XOR2_X1 U662 ( .A(KEYINPUT95), .B(KEYINPUT31), .Z(n566) );
  AND2_X1 U663 ( .A1(n685), .A2(n680), .ZN(n564) );
  NAND2_X1 U664 ( .A1(n593), .A2(n564), .ZN(n692) );
  XOR2_X1 U665 ( .A(n566), .B(n565), .Z(n667) );
  NOR2_X1 U666 ( .A1(n683), .A2(n680), .ZN(n567) );
  NAND2_X1 U667 ( .A1(n578), .A2(n567), .ZN(n568) );
  NOR2_X1 U668 ( .A1(n667), .A2(n650), .ZN(n569) );
  AND2_X1 U669 ( .A1(n658), .A2(n653), .ZN(n698) );
  NOR2_X1 U670 ( .A1(n569), .A2(n698), .ZN(n570) );
  NAND2_X1 U671 ( .A1(n700), .A2(n701), .ZN(n697) );
  NOR2_X1 U672 ( .A1(n703), .A2(n697), .ZN(n576) );
  NOR2_X1 U673 ( .A1(n716), .A2(n659), .ZN(n580) );
  XOR2_X1 U674 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n579) );
  XNOR2_X1 U675 ( .A(n580), .B(n579), .ZN(n753) );
  XNOR2_X1 U676 ( .A(n582), .B(KEYINPUT46), .ZN(n597) );
  INV_X1 U677 ( .A(n698), .ZN(n583) );
  NAND2_X1 U678 ( .A1(n583), .A2(KEYINPUT64), .ZN(n584) );
  INV_X1 U679 ( .A(n585), .ZN(n661) );
  NAND2_X1 U680 ( .A1(n586), .A2(n661), .ZN(n587) );
  NAND2_X1 U681 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U682 ( .A(KEYINPUT36), .B(n592), .Z(n594) );
  NAND2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n670) );
  XNOR2_X1 U684 ( .A(n595), .B(KEYINPUT67), .ZN(n596) );
  NAND2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U686 ( .A(KEYINPUT66), .B(KEYINPUT48), .ZN(n598) );
  INV_X1 U687 ( .A(n740), .ZN(n601) );
  INV_X1 U688 ( .A(n602), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n603), .A2(KEYINPUT2), .ZN(n604) );
  INV_X1 U690 ( .A(n672), .ZN(n726) );
  NAND2_X1 U691 ( .A1(n606), .A2(KEYINPUT2), .ZN(n607) );
  XOR2_X1 U692 ( .A(KEYINPUT77), .B(n607), .Z(n608) );
  NOR2_X1 U693 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U694 ( .A(n613), .B(n612), .ZN(n615) );
  INV_X1 U695 ( .A(G952), .ZN(n614) );
  INV_X1 U696 ( .A(n725), .ZN(n635) );
  NAND2_X1 U697 ( .A1(n615), .A2(n635), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U699 ( .A(KEYINPUT78), .B(KEYINPUT54), .ZN(n618) );
  XOR2_X1 U700 ( .A(n618), .B(KEYINPUT55), .Z(n619) );
  XNOR2_X1 U701 ( .A(n621), .B(n620), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n622), .A2(n635), .ZN(n624) );
  INV_X1 U703 ( .A(KEYINPUT56), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n624), .B(n623), .ZN(G51) );
  XNOR2_X1 U705 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n628), .A2(n635), .ZN(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT121), .B(KEYINPUT60), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n630), .B(n629), .ZN(G60) );
  XOR2_X1 U709 ( .A(KEYINPUT84), .B(KEYINPUT62), .Z(n631) );
  XNOR2_X1 U710 ( .A(n634), .B(n633), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n639) );
  XNOR2_X1 U712 ( .A(KEYINPUT85), .B(KEYINPUT63), .ZN(n637) );
  XOR2_X1 U713 ( .A(n637), .B(KEYINPUT82), .Z(n638) );
  XNOR2_X1 U714 ( .A(n639), .B(n638), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n722), .A2(G469), .ZN(n644) );
  XOR2_X1 U716 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n640) );
  XNOR2_X1 U717 ( .A(n640), .B(KEYINPUT58), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U719 ( .A(n644), .B(n643), .ZN(n645) );
  NOR2_X1 U720 ( .A1(n645), .A2(n725), .ZN(G54) );
  NAND2_X1 U721 ( .A1(n650), .A2(n664), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n646), .B(G104), .ZN(G6) );
  XOR2_X1 U723 ( .A(KEYINPUT109), .B(KEYINPUT27), .Z(n648) );
  XNOR2_X1 U724 ( .A(G107), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U725 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U726 ( .A(KEYINPUT108), .B(n649), .Z(n652) );
  NAND2_X1 U727 ( .A1(n650), .A2(n666), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n652), .B(n651), .ZN(G9) );
  XOR2_X1 U729 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n656) );
  NOR2_X1 U730 ( .A1(n659), .A2(n653), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n661), .A2(n654), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U733 ( .A(G128), .B(n657), .Z(G30) );
  NOR2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U735 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(KEYINPUT112), .ZN(n663) );
  XNOR2_X1 U737 ( .A(G146), .B(n663), .ZN(G48) );
  NAND2_X1 U738 ( .A1(n667), .A2(n664), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n665), .B(G113), .ZN(G15) );
  NAND2_X1 U740 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n668), .B(G116), .ZN(G18) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U743 ( .A(n671), .B(KEYINPUT37), .ZN(G27) );
  NOR2_X1 U744 ( .A1(n672), .A2(n740), .ZN(n673) );
  NOR2_X1 U745 ( .A1(n673), .A2(KEYINPUT2), .ZN(n676) );
  INV_X1 U746 ( .A(n674), .ZN(n675) );
  NOR2_X1 U747 ( .A1(n676), .A2(n675), .ZN(n714) );
  XOR2_X1 U748 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n695) );
  NOR2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U750 ( .A(KEYINPUT49), .B(n679), .Z(n681) );
  NOR2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n682), .B(KEYINPUT114), .ZN(n691) );
  NAND2_X1 U753 ( .A1(n687), .A2(n683), .ZN(n684) );
  NAND2_X1 U754 ( .A1(n684), .A2(KEYINPUT50), .ZN(n689) );
  NOR2_X1 U755 ( .A1(n685), .A2(KEYINPUT50), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n693) );
  AND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U760 ( .A(n695), .B(n694), .Z(n696) );
  NOR2_X1 U761 ( .A1(n716), .A2(n696), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U763 ( .A(KEYINPUT117), .B(n699), .Z(n706) );
  NOR2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U766 ( .A(KEYINPUT116), .B(n704), .ZN(n705) );
  NOR2_X1 U767 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U768 ( .A1(n708), .A2(n351), .ZN(n709) );
  XNOR2_X1 U769 ( .A(n709), .B(KEYINPUT52), .ZN(n710) );
  XNOR2_X1 U770 ( .A(KEYINPUT118), .B(n710), .ZN(n711) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n714), .A2(n713), .ZN(n719) );
  NOR2_X1 U773 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n717), .B(KEYINPUT119), .ZN(n718) );
  NAND2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n721), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U777 ( .A1(n722), .A2(G217), .ZN(n724) );
  NAND2_X1 U778 ( .A1(n726), .A2(n744), .ZN(n730) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n727) );
  XNOR2_X1 U780 ( .A(KEYINPUT61), .B(n727), .ZN(n728) );
  NAND2_X1 U781 ( .A1(n728), .A2(G898), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n736) );
  XOR2_X1 U783 ( .A(KEYINPUT124), .B(n731), .Z(n733) );
  NOR2_X1 U784 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U785 ( .A(KEYINPUT125), .B(n734), .Z(n735) );
  XNOR2_X1 U786 ( .A(n736), .B(n735), .ZN(G69) );
  XNOR2_X1 U787 ( .A(n737), .B(KEYINPUT126), .ZN(n739) );
  XNOR2_X1 U788 ( .A(n739), .B(n738), .ZN(n742) );
  XOR2_X1 U789 ( .A(n742), .B(n740), .Z(n741) );
  NAND2_X1 U790 ( .A1(n741), .A2(n744), .ZN(n747) );
  XOR2_X1 U791 ( .A(G227), .B(n742), .Z(n743) );
  NOR2_X1 U792 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U793 ( .A1(G900), .A2(n745), .ZN(n746) );
  NAND2_X1 U794 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U795 ( .A(KEYINPUT127), .B(n748), .ZN(G72) );
  XNOR2_X1 U796 ( .A(G101), .B(n750), .ZN(G3) );
  BUF_X1 U797 ( .A(n751), .Z(n752) );
  XNOR2_X1 U798 ( .A(n752), .B(G119), .ZN(G21) );
  XOR2_X1 U799 ( .A(G137), .B(n753), .Z(G39) );
endmodule

