//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n459), .A2(new_n461), .A3(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n460), .A2(KEYINPUT66), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n464), .A2(G2105), .B1(G101), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n470), .A2(G137), .A3(new_n471), .A4(new_n459), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n459), .ZN(new_n475));
  OR3_X1    g050(.A1(new_n475), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT67), .B1(new_n475), .B2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n471), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n471), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n481), .A2(G124), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n480), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  AND2_X1   g062(.A1(new_n471), .A2(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n470), .A2(new_n459), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n459), .A2(new_n461), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n492), .A2(new_n471), .A3(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n470), .A2(G126), .A3(G2105), .A4(new_n459), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT68), .A2(G114), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT68), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(G2104), .A3(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n496), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n494), .B1(new_n489), .B2(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n497), .A2(new_n502), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT69), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT71), .B1(new_n514), .B2(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n515), .B1(G75), .B2(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n514), .A2(KEYINPUT71), .A3(G62), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n520), .B1(new_n511), .B2(KEYINPUT6), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n522), .A2(KEYINPUT70), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n511), .A2(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(G543), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n524), .A2(new_n514), .A3(new_n525), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n519), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n518), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AND2_X1   g106(.A1(G63), .A2(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n535), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n514), .A2(new_n532), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G89), .ZN(new_n538));
  INV_X1    g113(.A(G51), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n537), .B1(new_n527), .B2(new_n538), .C1(new_n539), .C2(new_n526), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  INV_X1    g118(.A(new_n527), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n511), .ZN(new_n547));
  INV_X1    g122(.A(new_n526), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G52), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(new_n544), .A2(G81), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n511), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n548), .A2(G43), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND4_X1  g137(.A1(new_n524), .A2(G53), .A3(G543), .A4(new_n525), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n544), .A2(G91), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT73), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n514), .A2(G65), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n566), .A3(new_n568), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n564), .B(new_n565), .C1(new_n569), .C2(new_n571), .ZN(G299));
  XNOR2_X1  g147(.A(G168), .B(KEYINPUT74), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G286));
  NAND2_X1  g149(.A1(new_n548), .A2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n544), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT75), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n512), .B2(new_n513), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n524), .A2(G48), .A3(G543), .A4(new_n525), .ZN(new_n584));
  INV_X1    g159(.A(G86), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n527), .ZN(G305));
  NAND2_X1  g161(.A1(new_n544), .A2(G85), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n548), .A2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n587), .B(new_n588), .C1(new_n511), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n544), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n514), .A2(G66), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n511), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(G54), .B2(new_n548), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G321));
  NOR2_X1   g177(.A1(G299), .A2(G868), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n573), .B2(G868), .ZN(G297));
  AOI21_X1  g179(.A(new_n603), .B1(new_n573), .B2(G868), .ZN(G280));
  XNOR2_X1  g180(.A(KEYINPUT76), .B(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n600), .B1(G860), .B2(new_n606), .ZN(G148));
  OAI21_X1  g182(.A(KEYINPUT77), .B1(new_n557), .B2(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n606), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  MUX2_X1   g185(.A(KEYINPUT77), .B(new_n608), .S(new_n610), .Z(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g187(.A(new_n491), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n468), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT13), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n479), .A2(G135), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n471), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n481), .A2(G123), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n624), .A2(G2096), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(G2096), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n618), .A2(new_n625), .A3(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT79), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT80), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n638), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n639), .A2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n645), .B2(new_n641), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n644), .A2(new_n646), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT82), .ZN(new_n670));
  OR3_X1    g245(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1981), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G229));
  XOR2_X1   g253(.A(KEYINPUT84), .B(G16), .Z(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n680), .A2(G22), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G166), .B2(new_n680), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT87), .B(G1971), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  MUX2_X1   g259(.A(G6), .B(G305), .S(G16), .Z(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT86), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT32), .B(G1981), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G23), .ZN(new_n692));
  INV_X1    g267(.A(G288), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT33), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n684), .A2(new_n689), .A3(new_n690), .A4(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT88), .Z(new_n698));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n479), .A2(G131), .ZN(new_n704));
  OR2_X1    g279(.A1(G95), .A2(G2105), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n705), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT83), .Z(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G119), .B2(new_n481), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n703), .B1(new_n710), .B2(new_n702), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(new_n680), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT85), .B(G1986), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  NAND4_X1  g291(.A1(new_n700), .A2(new_n701), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n691), .A2(G5), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G171), .B2(new_n691), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT96), .ZN(new_n722));
  INV_X1    g297(.A(G1961), .ZN(new_n723));
  INV_X1    g298(.A(G2084), .ZN(new_n724));
  INV_X1    g299(.A(G34), .ZN(new_n725));
  AOI21_X1  g300(.A(G29), .B1(new_n725), .B2(KEYINPUT24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(KEYINPUT24), .B2(new_n725), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n473), .B2(new_n702), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n722), .A2(new_n723), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n702), .A2(G32), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n479), .A2(G141), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT26), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n468), .A2(G105), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n733), .B(new_n734), .C1(new_n481), .C2(G129), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(new_n702), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT93), .Z(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n729), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT97), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n702), .A2(G35), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G162), .B2(new_n702), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT29), .Z(new_n745));
  INV_X1    g320(.A(G2090), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT98), .Z(new_n748));
  XOR2_X1   g323(.A(KEYINPUT31), .B(G11), .Z(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT94), .B(G28), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT95), .Z(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n750), .B2(KEYINPUT30), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI221_X1 g329(.A(new_n754), .B1(new_n724), .B2(new_n728), .C1(new_n624), .C2(new_n702), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n691), .A2(G4), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n600), .B2(new_n691), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1348), .ZN(new_n758));
  NOR2_X1   g333(.A1(G27), .A2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G164), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2078), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n680), .A2(G19), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n557), .B2(new_n680), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1341), .ZN(new_n764));
  OR4_X1    g339(.A1(new_n755), .A2(new_n758), .A3(new_n761), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n702), .A2(G26), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n471), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n481), .A2(G128), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(G140), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n478), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT89), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n767), .B1(new_n774), .B2(new_n702), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2067), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n691), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n691), .ZN(new_n778));
  INV_X1    g353(.A(G1966), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n679), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT99), .B(G1956), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n780), .B(new_n785), .C1(new_n723), .C2(new_n722), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n765), .A2(new_n776), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n702), .A2(G33), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n479), .A2(G139), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT91), .Z(new_n790));
  XOR2_X1   g365(.A(KEYINPUT90), .B(KEYINPUT25), .Z(new_n791));
  NAND3_X1  g366(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n613), .A2(G127), .ZN(new_n794));
  NAND2_X1  g369(.A1(G115), .A2(G2104), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n471), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT92), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n788), .B1(new_n801), .B2(new_n702), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n746), .A2(new_n745), .B1(new_n802), .B2(G2072), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(G2072), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n739), .A2(new_n740), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n803), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n742), .A2(new_n748), .A3(new_n787), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n719), .A2(new_n807), .ZN(G311));
  OR2_X1    g383(.A1(new_n719), .A2(new_n807), .ZN(G150));
  NAND2_X1  g384(.A1(new_n544), .A2(G93), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n548), .A2(G55), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n810), .B(new_n811), .C1(new_n511), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT100), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(new_n557), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n813), .A2(new_n556), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n600), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT101), .B(G860), .Z(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n815), .A2(new_n824), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT102), .Z(G145));
  NOR2_X1   g404(.A1(new_n506), .A2(new_n507), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n774), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n774), .A2(new_n830), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n801), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n774), .B(new_n830), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(new_n800), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(new_n737), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n471), .A2(G118), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n481), .A2(G130), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G142), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n478), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n616), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(new_n709), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n833), .A2(new_n736), .A3(new_n835), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n837), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n845), .B(KEYINPUT103), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n837), .B2(new_n847), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n624), .B(new_n473), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n486), .ZN(new_n853));
  AOI21_X1  g428(.A(G37), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n848), .B2(new_n850), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g433(.A1(new_n600), .A2(G299), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n600), .A2(G299), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT105), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n865), .A3(new_n862), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT104), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n859), .A2(new_n867), .A3(new_n860), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n600), .A2(KEYINPUT104), .A3(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n864), .B(new_n866), .C1(new_n871), .C2(new_n862), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n818), .B(new_n609), .Z(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n870), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n877));
  XNOR2_X1  g452(.A(G303), .B(new_n693), .ZN(new_n878));
  XOR2_X1   g453(.A(G290), .B(G305), .Z(new_n879));
  XOR2_X1   g454(.A(new_n878), .B(new_n879), .Z(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(KEYINPUT42), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n877), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(G868), .B2(new_n815), .ZN(G295));
  OAI21_X1  g460(.A(new_n884), .B1(G868), .B2(new_n815), .ZN(G331));
  NAND2_X1  g461(.A1(new_n573), .A2(G171), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n541), .A2(new_n542), .A3(G301), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n818), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n818), .A2(new_n887), .A3(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n861), .A2(new_n862), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT107), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(KEYINPUT107), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n898), .B(new_n899), .C1(KEYINPUT41), .C2(new_n870), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n889), .A2(new_n890), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n871), .A2(new_n895), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n896), .A2(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n880), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  INV_X1    g481(.A(new_n893), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n902), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n901), .A2(new_n895), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n872), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n911), .A3(new_n904), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n905), .A2(new_n906), .A3(new_n914), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n894), .A2(new_n902), .B1(new_n872), .B2(new_n910), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(new_n904), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT44), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n916), .B2(new_n904), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(new_n906), .C1(new_n904), .C2(new_n903), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n914), .B2(new_n917), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n920), .B1(KEYINPUT44), .B2(new_n925), .ZN(G397));
  XNOR2_X1  g501(.A(new_n774), .B(G2067), .ZN(new_n927));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n736), .B(new_n928), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n710), .A2(new_n712), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n710), .A2(new_n712), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n927), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n464), .A2(G2105), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n468), .A2(G101), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n933), .A2(G40), .A3(new_n472), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n469), .A2(KEYINPUT109), .A3(G40), .A4(new_n472), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(KEYINPUT108), .B(G1384), .Z(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n506), .B2(new_n507), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n932), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(G290), .A2(G1986), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  NAND2_X1  g523(.A1(G290), .A2(G1986), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n950), .B(new_n944), .C1(new_n948), .C2(new_n949), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT111), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT112), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(new_n506), .B2(new_n507), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT113), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n955), .C1(new_n506), .C2(new_n507), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n942), .A3(new_n959), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n937), .A2(new_n938), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(KEYINPUT115), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(G1384), .B1(new_n505), .B2(new_n508), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT115), .B1(new_n960), .B2(new_n961), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n779), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n968), .B1(new_n509), .B2(new_n955), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT50), .B1(new_n957), .B2(new_n959), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(new_n939), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n724), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(G168), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(G8), .ZN(new_n974));
  AOI21_X1  g549(.A(G168), .B1(new_n967), .B2(new_n972), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT51), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n977), .A3(G8), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT62), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n976), .B2(new_n978), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n957), .A2(new_n959), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n961), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n693), .A2(G1976), .ZN(new_n984));
  INV_X1    g559(.A(G1976), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(G288), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n983), .A2(G8), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(G305), .A2(G1981), .ZN(new_n988));
  NOR2_X1   g563(.A1(G305), .A2(G1981), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n990));
  OR3_X1    g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n988), .B2(new_n989), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n991), .A2(new_n983), .A3(G8), .A4(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n983), .A2(G8), .A3(new_n984), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n995));
  OAI211_X1 g570(.A(new_n987), .B(new_n993), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G8), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT55), .Z(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n939), .B1(new_n982), .B2(new_n968), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n504), .B1(new_n496), .B2(new_n503), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT69), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n955), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT50), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1000), .A2(new_n746), .A3(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT45), .B(new_n940), .C1(new_n506), .C2(new_n507), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1006), .A2(new_n937), .A3(new_n938), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(KEYINPUT45), .B2(new_n963), .ZN(new_n1008));
  INV_X1    g583(.A(G1971), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n999), .B1(new_n1005), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n996), .B1(new_n998), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n997), .B(KEYINPUT55), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n968), .B(new_n955), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n957), .A2(KEYINPUT50), .A3(new_n959), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n961), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  AOI21_X1  g592(.A(G2090), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n939), .B1(new_n963), .B2(new_n968), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1019), .A2(KEYINPUT114), .A3(new_n1015), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1018), .A2(new_n1020), .B1(new_n1009), .B2(new_n1008), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1013), .B1(new_n1021), .B2(new_n999), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n982), .A2(new_n968), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1004), .A2(new_n1023), .A3(new_n961), .ZN(new_n1024));
  INV_X1    g599(.A(G2078), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1007), .B(new_n1025), .C1(KEYINPUT45), .C2(new_n963), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1024), .A2(new_n723), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n960), .A2(new_n961), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1027), .A2(G2078), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1031), .A2(new_n964), .A3(new_n962), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G301), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1012), .A2(new_n1022), .A3(new_n1034), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n980), .A2(new_n981), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1024), .A2(new_n723), .ZN(new_n1038));
  INV_X1    g613(.A(new_n935), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n943), .A2(KEYINPUT121), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT121), .B1(new_n943), .B2(new_n1039), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1006), .B(new_n1032), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1043));
  AND4_X1   g618(.A1(G301), .A2(new_n1038), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1037), .B1(new_n1044), .B2(new_n1034), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT122), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n1037), .C1(new_n1044), .C2(new_n1034), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n976), .A2(new_n978), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT117), .B(G1956), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1019), .B2(new_n1015), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT45), .B1(new_n509), .B2(new_n955), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1006), .A2(new_n937), .A3(new_n938), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(G299), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n565), .B1(new_n571), .B2(new_n569), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT9), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n563), .B(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1058), .A2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1052), .A2(new_n1057), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1051), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1054), .B1(new_n1003), .B2(new_n942), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1016), .A2(new_n1068), .B1(new_n1069), .B2(new_n1055), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1058), .A2(new_n1064), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT119), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1065), .C1(new_n1052), .C2(new_n1057), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G1348), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1076));
  INV_X1    g651(.A(G2067), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n982), .A2(new_n961), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(new_n599), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1067), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1016), .A2(new_n1068), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1069), .A2(new_n1055), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1071), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1083), .B1(new_n1066), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT60), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT60), .B(new_n1078), .C1(new_n971), .C2(G1348), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(new_n600), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(G1341), .Z(new_n1093));
  AOI22_X1  g668(.A1(new_n1069), .A2(new_n928), .B1(new_n983), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT59), .B1(new_n1094), .B2(new_n556), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1008), .A2(G1996), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1093), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n982), .B2(new_n961), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1096), .B(new_n557), .C1(new_n1097), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1087), .A2(new_n1091), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1083), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1104));
  AND3_X1   g679(.A1(new_n1072), .A2(new_n1104), .A3(new_n1074), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1082), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1028), .A2(G301), .A3(new_n1033), .ZN(new_n1107));
  AOI21_X1  g682(.A(G301), .B1(new_n1028), .B2(new_n1042), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1037), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1012), .A2(new_n1022), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1049), .A2(new_n1050), .A3(new_n1106), .A4(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n993), .A2(new_n985), .A3(new_n693), .ZN(new_n1113));
  OAI211_X1 g688(.A(G8), .B(new_n983), .C1(new_n1113), .C2(new_n989), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1011), .A2(new_n998), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1114), .B1(new_n1115), .B2(new_n996), .ZN(new_n1116));
  NOR2_X1   g691(.A1(G286), .A2(new_n999), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n967), .A2(new_n972), .ZN(new_n1118));
  AND4_X1   g693(.A1(KEYINPUT63), .A2(new_n1115), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(G8), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n996), .B1(new_n1121), .B2(new_n1013), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(KEYINPUT116), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1011), .A2(new_n998), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1124), .A2(new_n1125), .A3(new_n996), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1119), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1128), .B1(new_n1110), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1116), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1112), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1036), .B1(new_n1132), .B2(KEYINPUT123), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1112), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n954), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n927), .A2(new_n737), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n944), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n944), .A2(new_n928), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT46), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT124), .B(KEYINPUT47), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1146));
  INV_X1    g721(.A(new_n945), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n944), .A2(new_n946), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT48), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n774), .A2(new_n1077), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n927), .A2(new_n929), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n931), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1147), .A2(new_n1149), .B1(new_n944), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1145), .A2(new_n1146), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT126), .B1(new_n1136), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1154), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1112), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1134), .B1(new_n1112), .B2(new_n1131), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1036), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1156), .B(new_n1157), .C1(new_n1160), .C2(new_n954), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1155), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g737(.A(G319), .ZN(new_n1164));
  NOR3_X1   g738(.A1(G229), .A2(new_n1164), .A3(G227), .ZN(new_n1165));
  OAI21_X1  g739(.A(new_n1165), .B1(new_n644), .B2(new_n646), .ZN(new_n1166));
  AOI21_X1  g740(.A(new_n1166), .B1(new_n854), .B2(new_n856), .ZN(new_n1167));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n1168));
  AND3_X1   g742(.A1(new_n924), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g743(.A(new_n1168), .B1(new_n924), .B2(new_n1167), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1169), .A2(new_n1170), .ZN(G308));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n1167), .ZN(G225));
endmodule


