//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT64), .A2(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OR2_X1    g011(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT66), .A2(KEYINPUT1), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  INV_X1    g016(.A(new_n199), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT64), .B(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G146), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n206), .B1(new_n198), .B2(new_n200), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n197), .A2(new_n202), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n209), .B1(new_n210), .B2(G137), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT65), .A3(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT11), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n210), .B2(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n212), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n189), .B1(new_n208), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n219), .A3(new_n212), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n221), .ZN(new_n226));
  INV_X1    g040(.A(new_n194), .ZN(new_n227));
  NOR2_X1   g041(.A1(KEYINPUT64), .A2(G143), .ZN(new_n228));
  OAI21_X1  g042(.A(G146), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n199), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n197), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n226), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n202), .A2(new_n197), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n207), .A2(new_n229), .A3(new_n199), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n216), .A2(new_n221), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT67), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n223), .A2(new_n235), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT2), .B(G113), .Z(new_n248));
  OR2_X1    g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n248), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n241), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n238), .A2(new_n239), .ZN(new_n253));
  INV_X1    g067(.A(new_n251), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n235), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT28), .A4(new_n235), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G237), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(G210), .ZN(new_n262));
  INV_X1    g076(.A(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n265));
  XOR2_X1   g079(.A(new_n264), .B(new_n265), .Z(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n188), .B1(new_n259), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n241), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n253), .A2(new_n235), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT30), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n251), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n266), .B1(new_n273), .B2(new_n255), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n187), .B1(new_n268), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G902), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n257), .A2(new_n258), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n271), .A2(new_n254), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n275), .B(new_n276), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n268), .A2(new_n274), .A3(new_n187), .ZN(new_n282));
  OAI21_X1  g096(.A(G472), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(new_n255), .A3(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT31), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n273), .A2(new_n286), .A3(new_n255), .A4(new_n266), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n234), .A2(new_n231), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n253), .A2(new_n189), .B1(new_n289), .B2(new_n226), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n254), .B1(new_n290), .B2(new_n240), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n267), .B1(new_n277), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT68), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n259), .A2(new_n294), .A3(new_n267), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n285), .A2(new_n287), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G472), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n296), .A2(new_n297), .A3(new_n276), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n298), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n299));
  AOI21_X1  g113(.A(KEYINPUT32), .B1(new_n298), .B2(KEYINPUT69), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n283), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  OAI21_X1  g116(.A(G221), .B1(new_n302), .B2(G902), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n303), .B(KEYINPUT77), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n261), .A2(G227), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT78), .ZN(new_n307));
  XNOR2_X1  g121(.A(G110), .B(G140), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n311));
  INV_X1    g125(.A(G107), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(G104), .ZN(new_n313));
  INV_X1    g127(.A(G104), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT3), .B1(new_n314), .B2(G107), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(G107), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n263), .B(new_n313), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n312), .A2(G104), .ZN(new_n318));
  OAI21_X1  g132(.A(G101), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n236), .A2(new_n237), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n206), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n237), .B1(new_n323), .B2(new_n205), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n317), .A2(new_n319), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n236), .A2(new_n320), .A3(new_n327), .A4(new_n237), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT12), .A3(new_n226), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n329), .A2(KEYINPUT81), .A3(KEYINPUT12), .A4(new_n226), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n226), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT12), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n237), .ZN(new_n338));
  AOI22_X1  g152(.A1(G128), .A2(new_n201), .B1(new_n195), .B2(new_n196), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n325), .B(KEYINPUT10), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT79), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n238), .A2(new_n342), .A3(KEYINPUT10), .A4(new_n325), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n317), .A2(KEYINPUT4), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n348), .A2(new_n289), .B1(new_n326), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n226), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n344), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n310), .B1(new_n337), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n310), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n344), .A2(new_n350), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n351), .B1(new_n355), .B2(KEYINPUT82), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n350), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n276), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G469), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n344), .A2(new_n350), .A3(new_n357), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n357), .B1(new_n344), .B2(new_n350), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n362), .A2(new_n363), .A3(new_n351), .ZN(new_n364));
  INV_X1    g178(.A(new_n352), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n309), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n354), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n337), .ZN(new_n368));
  AOI21_X1  g182(.A(G902), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G469), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n361), .A2(KEYINPUT83), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n360), .A2(G469), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT83), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n305), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT74), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G137), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n380), .A2(KEYINPUT16), .A3(G140), .ZN(new_n381));
  XNOR2_X1  g195(.A(G125), .B(G140), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(new_n382), .B2(KEYINPUT16), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G146), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G125), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n380), .A2(G140), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT16), .ZN(new_n388));
  OR3_X1    g202(.A1(new_n380), .A2(KEYINPUT16), .A3(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n193), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n242), .A2(KEYINPUT23), .A3(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n242), .A2(G128), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT23), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(G119), .B2(new_n206), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n384), .A2(new_n391), .B1(G110), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g211(.A(KEYINPUT24), .B(G110), .Z(new_n398));
  INV_X1    g212(.A(KEYINPUT71), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n206), .B2(G119), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n242), .A2(KEYINPUT71), .A3(G128), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n206), .A2(G119), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT72), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n400), .A2(new_n401), .B1(G119), .B2(new_n206), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT72), .A3(new_n398), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n397), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n382), .A2(new_n193), .ZN(new_n411));
  OAI22_X1  g225(.A1(new_n396), .A2(G110), .B1(new_n407), .B2(new_n398), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT73), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n413), .B1(new_n383), .B2(G146), .ZN(new_n414));
  AND4_X1   g228(.A1(new_n413), .A2(new_n388), .A3(G146), .A4(new_n389), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n411), .B(new_n412), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n379), .B1(new_n417), .B2(KEYINPUT75), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT75), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n410), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  AND4_X1   g235(.A1(new_n419), .A2(new_n410), .A3(new_n416), .A4(new_n379), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G217), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n425), .B1(G234), .B2(new_n276), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G902), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n410), .A2(new_n419), .A3(new_n416), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n419), .B1(new_n410), .B2(new_n416), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n429), .A2(new_n430), .A3(new_n379), .ZN(new_n431));
  OAI211_X1 g245(.A(KEYINPUT25), .B(new_n276), .C1(new_n431), .C2(new_n422), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT76), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT25), .B1(new_n424), .B2(new_n276), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n276), .B1(new_n431), .B2(new_n422), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n426), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n428), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n382), .B(new_n193), .ZN(new_n443));
  INV_X1    g257(.A(G214), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n444), .A2(G237), .A3(G953), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G143), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n227), .A2(new_n228), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n446), .B(new_n447), .C1(new_n448), .C2(new_n445), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n446), .B(new_n220), .C1(new_n448), .C2(new_n445), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n443), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n448), .A2(new_n445), .ZN(new_n452));
  INV_X1    g266(.A(new_n446), .ZN(new_n453));
  OAI21_X1  g267(.A(G131), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n447), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n454), .ZN(new_n456));
  INV_X1    g270(.A(new_n450), .ZN(new_n457));
  NOR3_X1   g271(.A1(new_n456), .A2(KEYINPUT17), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n391), .B(new_n384), .C1(new_n454), .C2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n455), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G113), .B(G122), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(new_n314), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n463), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n382), .B(KEYINPUT19), .Z(new_n466));
  OAI22_X1  g280(.A1(new_n456), .A2(new_n457), .B1(G146), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n414), .A2(new_n415), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n455), .B(new_n465), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(G475), .A2(G902), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n464), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT20), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT20), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n464), .A2(new_n473), .A3(new_n469), .A4(new_n470), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n463), .A2(KEYINPUT87), .ZN(new_n475));
  AOI21_X1  g289(.A(G902), .B1(new_n461), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n476), .B1(new_n475), .B2(new_n461), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n472), .A2(new_n474), .B1(new_n477), .B2(G475), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(G234), .A2(G237), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n480), .A2(G952), .A3(new_n261), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT21), .B(G898), .Z(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n480), .A2(G902), .A3(G953), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G214), .B1(G237), .B2(G902), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT5), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n242), .A3(G116), .ZN(new_n490));
  OAI211_X1 g304(.A(G113), .B(new_n490), .C1(new_n246), .C2(new_n489), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n250), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(new_n320), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n345), .A2(G101), .A3(new_n346), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n347), .A2(KEYINPUT4), .A3(new_n317), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n251), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G110), .B(G122), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n288), .A2(G125), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n236), .A2(new_n380), .A3(new_n237), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT85), .B(G224), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(new_n504), .B2(G953), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n505), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n501), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n498), .B(KEYINPUT8), .ZN(new_n509));
  AND2_X1   g323(.A1(new_n492), .A2(new_n320), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n493), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n500), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n506), .A2(new_n511), .A3(new_n508), .A4(KEYINPUT86), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n494), .A2(new_n497), .ZN(new_n517));
  INV_X1    g331(.A(new_n498), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT6), .A4(new_n499), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n504), .A2(G953), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n503), .B(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n516), .A2(new_n276), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G210), .B1(G237), .B2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n514), .B2(new_n515), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n528), .A3(new_n526), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n488), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n244), .A2(G122), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n535));
  INV_X1    g349(.A(G122), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G116), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n244), .A2(G122), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(KEYINPUT89), .A3(KEYINPUT14), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n537), .B2(new_n535), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n538), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G107), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n191), .B2(G128), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n206), .A2(KEYINPUT88), .A3(G143), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(G134), .C1(new_n448), .C2(new_n206), .ZN(new_n549));
  OR3_X1    g363(.A1(new_n537), .A2(new_n534), .A3(G107), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n448), .B2(new_n206), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n210), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n544), .A2(new_n549), .A3(new_n550), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n210), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n551), .ZN(new_n556));
  OAI221_X1 g370(.A(new_n548), .B1(new_n554), .B2(new_n210), .C1(new_n448), .C2(new_n206), .ZN(new_n557));
  OAI21_X1  g371(.A(G107), .B1(new_n537), .B2(new_n534), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n302), .A2(new_n425), .A3(G953), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n553), .A2(new_n560), .A3(new_n562), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n564), .A2(KEYINPUT90), .A3(new_n565), .ZN(new_n566));
  OR3_X1    g380(.A1(new_n561), .A2(KEYINPUT90), .A3(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n276), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT91), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n566), .A2(new_n567), .A3(new_n572), .A4(new_n276), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n568), .B(KEYINPUT91), .C1(KEYINPUT15), .C2(new_n570), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(KEYINPUT92), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT92), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n574), .B2(new_n575), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n486), .B(new_n533), .C1(new_n577), .C2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n301), .A2(new_n375), .A3(new_n442), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  XOR2_X1   g397(.A(KEYINPUT93), .B(KEYINPUT33), .Z(new_n584));
  NAND3_X1  g398(.A1(new_n566), .A2(new_n567), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT94), .A4(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n565), .ZN(new_n590));
  OR3_X1    g404(.A1(new_n590), .A2(new_n564), .A3(KEYINPUT95), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n564), .B1(new_n590), .B2(KEYINPUT95), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(KEYINPUT33), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n570), .A2(G902), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT96), .B(G478), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n568), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n479), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n485), .ZN(new_n600));
  INV_X1    g414(.A(new_n532), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n528), .B1(new_n531), .B2(new_n526), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n487), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT97), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n488), .B(new_n485), .C1(new_n530), .C2(new_n532), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n478), .B1(new_n607), .B2(new_n597), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n605), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n298), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n297), .B1(new_n296), .B2(new_n276), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n611), .A2(new_n441), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n375), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT98), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  NAND3_X1  g431(.A1(new_n375), .A2(new_n605), .A3(new_n613), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n576), .B(KEYINPUT92), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n618), .A2(new_n619), .A3(new_n479), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G107), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NOR2_X1   g436(.A1(new_n611), .A2(new_n612), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n417), .B(KEYINPUT99), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n379), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n427), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n627), .B1(new_n435), .B2(new_n440), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n375), .A2(new_n581), .A3(new_n623), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT37), .B(G110), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G12));
  INV_X1    g445(.A(new_n628), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n298), .A2(KEYINPUT69), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT32), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n298), .A2(KEYINPUT69), .A3(KEYINPUT32), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n632), .B1(new_n637), .B2(new_n283), .ZN(new_n638));
  INV_X1    g452(.A(G900), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n484), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n481), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n619), .A2(new_n479), .A3(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n638), .A2(new_n375), .A3(new_n533), .A4(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  NOR2_X1   g460(.A1(new_n577), .A2(new_n579), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n479), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n648), .A2(new_n488), .A3(new_n628), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(KEYINPUT100), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(KEYINPUT100), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n530), .A2(new_n532), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT38), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n651), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n642), .B(KEYINPUT39), .Z(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n375), .A2(new_n658), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(KEYINPUT40), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n273), .A2(new_n255), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n267), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n267), .A2(new_n255), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n276), .B1(new_n278), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n637), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n656), .A2(new_n660), .A3(new_n661), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n448), .B(KEYINPUT101), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G45));
  AOI211_X1 g485(.A(new_n643), .B(new_n478), .C1(new_n607), .C2(new_n597), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n638), .A2(new_n375), .A3(new_n533), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  NAND2_X1  g488(.A1(new_n356), .A2(new_n358), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n310), .B1(new_n675), .B2(new_n352), .ZN(new_n676));
  INV_X1    g490(.A(new_n368), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(G469), .B1(new_n678), .B2(G902), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n370), .B(new_n276), .C1(new_n676), .C2(new_n677), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n303), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n610), .A2(new_n301), .A3(new_n442), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NOR3_X1   g500(.A1(new_n619), .A2(new_n479), .A3(new_n603), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n301), .A2(new_n687), .A3(new_n683), .A4(new_n442), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NAND4_X1  g503(.A1(new_n679), .A2(new_n303), .A3(new_n680), .A4(new_n533), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n486), .B1(new_n577), .B2(new_n579), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n301), .A3(new_n628), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  XNOR2_X1  g508(.A(new_n441), .B(KEYINPUT104), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n603), .A2(new_n577), .A3(new_n579), .A4(new_n478), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n296), .A2(new_n276), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT103), .B(G472), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n279), .A2(new_n267), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n285), .A2(new_n287), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(G472), .A2(G902), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n701), .A2(KEYINPUT102), .A3(new_n702), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n699), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n695), .A2(new_n683), .A3(new_n696), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  INV_X1    g523(.A(new_n672), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n699), .A2(new_n628), .A3(new_n705), .A4(new_n706), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n701), .A2(KEYINPUT102), .A3(new_n702), .ZN(new_n714));
  AOI21_X1  g528(.A(KEYINPUT102), .B1(new_n701), .B2(new_n702), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(KEYINPUT105), .A3(new_n628), .A4(new_n699), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n710), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n690), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  AOI21_X1  g535(.A(new_n441), .B1(new_n637), .B2(new_n283), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n682), .B1(new_n361), .B2(new_n680), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n653), .A2(new_n488), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n722), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n298), .A2(new_n634), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n611), .A2(KEYINPUT32), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n298), .A2(KEYINPUT106), .A3(new_n634), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n733), .A3(new_n283), .A4(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n723), .A2(new_n672), .A3(new_n725), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n695), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n729), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n220), .ZN(G33));
  NAND4_X1  g554(.A1(new_n727), .A2(new_n301), .A3(new_n644), .A4(new_n442), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G134), .ZN(G36));
  OR2_X1    g556(.A1(new_n353), .A2(new_n359), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n744), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(G469), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(G469), .A2(G902), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT46), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n680), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n749), .A2(KEYINPUT46), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n303), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(new_n657), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n479), .B1(new_n607), .B2(new_n597), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(KEYINPUT107), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT43), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n758), .A2(new_n623), .A3(new_n632), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n726), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n755), .B(new_n761), .C1(new_n760), .C2(new_n759), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT108), .B(G137), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G39));
  XNOR2_X1  g578(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n753), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n725), .A2(new_n642), .ZN(new_n767));
  OR4_X1    g581(.A1(new_n301), .A2(new_n442), .A3(new_n599), .A4(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  XOR2_X1   g584(.A(new_n681), .B(KEYINPUT49), .Z(new_n771));
  NOR3_X1   g585(.A1(new_n654), .A2(new_n305), .A3(new_n488), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n756), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n695), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n773), .A2(new_n668), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n766), .B1(new_n304), .B2(new_n681), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n758), .A2(new_n641), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n695), .A2(new_n707), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(new_n725), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n654), .A2(new_n487), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n683), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n777), .A2(new_n781), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n683), .A2(new_n725), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n790), .A2(new_n668), .A3(new_n441), .A4(new_n641), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n595), .A2(new_n479), .A3(new_n598), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n758), .A2(new_n641), .A3(new_n790), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n713), .A2(new_n717), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n789), .A2(KEYINPUT51), .B1(new_n787), .B2(new_n795), .ZN(new_n796));
  AND4_X1   g610(.A1(KEYINPUT112), .A2(new_n787), .A3(KEYINPUT51), .A4(new_n795), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n735), .A2(new_n695), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT48), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n780), .A2(new_n533), .A3(new_n683), .ZN(new_n801));
  INV_X1    g615(.A(G952), .ZN(new_n802));
  AOI211_X1 g616(.A(new_n802), .B(G953), .C1(new_n791), .C2(new_n608), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n796), .A2(new_n797), .A3(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n724), .A2(new_n628), .A3(new_n643), .ZN(new_n806));
  INV_X1    g620(.A(new_n533), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n648), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n668), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n645), .A2(new_n673), .A3(new_n720), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n301), .A2(new_n375), .A3(new_n533), .A4(new_n628), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n812), .A2(new_n644), .B1(new_n719), .B2(new_n718), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n673), .A4(new_n809), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n582), .A2(new_n693), .A3(new_n708), .A4(new_n629), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n608), .A2(KEYINPUT110), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n574), .A2(new_n575), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n820), .B1(new_n821), .B2(new_n478), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n822), .B2(new_n608), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n375), .A2(new_n823), .A3(new_n605), .A4(new_n613), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n684), .A2(new_n688), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n729), .A2(new_n738), .A3(new_n741), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n301), .A2(new_n375), .A3(new_n628), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n767), .A2(new_n821), .A3(new_n479), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n828), .A2(new_n829), .B1(new_n718), .B2(new_n727), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n826), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n816), .A2(new_n817), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n816), .A2(KEYINPUT111), .ZN(new_n833));
  INV_X1    g647(.A(new_n831), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n811), .A2(new_n815), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(KEYINPUT54), .B(new_n832), .C1(new_n837), .C2(new_n817), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n817), .B1(new_n816), .B2(new_n831), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n839), .B1(new_n837), .B2(new_n817), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n838), .B1(KEYINPUT54), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n805), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(G952), .A2(G953), .ZN(new_n843));
  OAI211_X1 g657(.A(KEYINPUT113), .B(new_n776), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n843), .B1(new_n805), .B2(new_n841), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(new_n775), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n847), .ZN(G75));
  NAND2_X1  g662(.A1(new_n521), .A2(new_n523), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(new_n525), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n831), .B1(new_n816), .B2(KEYINPUT111), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT53), .B1(new_n852), .B2(new_n836), .ZN(new_n853));
  OAI211_X1 g667(.A(G210), .B(G902), .C1(new_n853), .C2(new_n832), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n855), .B1(new_n854), .B2(new_n857), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n860), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n850), .A3(new_n858), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n261), .A2(G952), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n861), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n861), .A2(new_n863), .A3(KEYINPUT115), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(G51));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n837), .A2(new_n817), .ZN(new_n872));
  INV_X1    g686(.A(new_n832), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n747), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(G902), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT117), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n874), .A2(KEYINPUT117), .A3(G902), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n748), .B(KEYINPUT57), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n872), .B2(new_n873), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n884), .B2(new_n838), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n678), .B1(new_n885), .B2(KEYINPUT116), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n872), .A2(new_n883), .A3(new_n873), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT54), .B1(new_n853), .B2(new_n832), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n880), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n871), .B1(new_n892), .B2(new_n864), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n878), .A2(new_n879), .ZN(new_n894));
  INV_X1    g708(.A(new_n891), .ZN(new_n895));
  INV_X1    g709(.A(new_n678), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n889), .B2(new_n890), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n898), .A2(KEYINPUT118), .A3(new_n865), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n893), .A2(new_n899), .ZN(G54));
  NAND4_X1  g714(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n464), .A2(new_n469), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n901), .A2(KEYINPUT119), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT119), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n864), .B1(new_n901), .B2(new_n902), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT120), .ZN(G60));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT59), .Z(new_n909));
  NOR2_X1   g723(.A1(new_n841), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n589), .A2(new_n593), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n865), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n909), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n911), .B(new_n913), .C1(new_n884), .C2(new_n838), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(KEYINPUT121), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(KEYINPUT121), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(G63));
  INV_X1    g731(.A(KEYINPUT61), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n919));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT60), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n872), .B2(new_n873), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(new_n424), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n864), .B1(new_n922), .B2(new_n626), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n918), .A2(KEYINPUT122), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n925), .B(new_n926), .Z(G66));
  OAI21_X1  g741(.A(G953), .B1(new_n483), .B2(new_n504), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n826), .B2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n849), .B1(G898), .B2(new_n261), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  AOI21_X1  g745(.A(new_n261), .B1(G227), .B2(G900), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT124), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n270), .A2(new_n272), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n466), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n639), .A2(new_n261), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n755), .A2(new_n798), .A3(new_n808), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n769), .A2(new_n827), .A3(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n813), .A2(new_n673), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n762), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT126), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n762), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  AOI211_X1 g758(.A(new_n935), .B(new_n936), .C1(new_n944), .C2(new_n261), .ZN(new_n945));
  INV_X1    g759(.A(new_n935), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n669), .A2(new_n939), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  INV_X1    g762(.A(new_n659), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n722), .A3(new_n725), .A4(new_n823), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n769), .A2(new_n762), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n946), .B1(new_n953), .B2(new_n261), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n933), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n954), .B(KEYINPUT123), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n933), .B(KEYINPUT125), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n945), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n955), .B1(new_n956), .B2(new_n958), .ZN(G72));
  NAND2_X1  g773(.A1(G472), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT63), .Z(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n274), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n284), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n840), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n952), .B2(new_n826), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n966), .A2(new_n663), .A3(new_n267), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n962), .B1(new_n944), .B2(new_n826), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n663), .A2(new_n267), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n865), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(KEYINPUT127), .B(new_n865), .C1(new_n968), .C2(new_n969), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n965), .B(new_n967), .C1(new_n972), .C2(new_n973), .ZN(G57));
endmodule


