

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U326 ( .A(n395), .B(KEYINPUT98), .ZN(n396) );
  XNOR2_X1 U327 ( .A(n454), .B(n453), .ZN(n487) );
  XNOR2_X1 U328 ( .A(n397), .B(n396), .ZN(n401) );
  XNOR2_X1 U329 ( .A(n334), .B(n312), .ZN(n313) );
  XNOR2_X1 U330 ( .A(n319), .B(n318), .ZN(n386) );
  XOR2_X1 U331 ( .A(n404), .B(KEYINPUT28), .Z(n512) );
  XNOR2_X1 U332 ( .A(n489), .B(n488), .ZN(n511) );
  NOR2_X1 U333 ( .A1(n566), .A2(n570), .ZN(n568) );
  XOR2_X1 U334 ( .A(n321), .B(n320), .Z(n294) );
  XOR2_X1 U335 ( .A(KEYINPUT10), .B(G36GAT), .Z(n295) );
  XOR2_X1 U336 ( .A(n437), .B(n436), .Z(n296) );
  XNOR2_X1 U337 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n465) );
  XNOR2_X1 U338 ( .A(n466), .B(n465), .ZN(n468) );
  INV_X1 U339 ( .A(G148GAT), .ZN(n316) );
  XNOR2_X1 U340 ( .A(n311), .B(KEYINPUT71), .ZN(n312) );
  NOR2_X1 U341 ( .A1(n495), .A2(n584), .ZN(n434) );
  XNOR2_X1 U342 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n363) );
  XNOR2_X1 U343 ( .A(n317), .B(n316), .ZN(n319) );
  INV_X1 U344 ( .A(KEYINPUT37), .ZN(n452) );
  XNOR2_X1 U345 ( .A(n452), .B(KEYINPUT105), .ZN(n453) );
  XNOR2_X1 U346 ( .A(n386), .B(n294), .ZN(n322) );
  XNOR2_X1 U347 ( .A(n478), .B(KEYINPUT122), .ZN(n479) );
  XNOR2_X1 U348 ( .A(n472), .B(KEYINPUT48), .ZN(n534) );
  XOR2_X1 U349 ( .A(n393), .B(n392), .Z(n477) );
  XNOR2_X1 U350 ( .A(n323), .B(n322), .ZN(n459) );
  XNOR2_X1 U351 ( .A(n399), .B(n398), .ZN(n575) );
  XNOR2_X1 U352 ( .A(n450), .B(n449), .ZN(n548) );
  XNOR2_X1 U353 ( .A(KEYINPUT110), .B(n455), .ZN(n532) );
  INV_X1 U354 ( .A(G29GAT), .ZN(n490) );
  XNOR2_X1 U355 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U356 ( .A(n456), .B(G106GAT), .ZN(n457) );
  XNOR2_X1 U357 ( .A(n490), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U358 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U359 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  XOR2_X1 U360 ( .A(G36GAT), .B(G8GAT), .Z(n369) );
  XOR2_X1 U361 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n298) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(G169GAT), .ZN(n297) );
  XNOR2_X1 U363 ( .A(n298), .B(n297), .ZN(n301) );
  XOR2_X1 U364 ( .A(G1GAT), .B(G22GAT), .Z(n414) );
  XNOR2_X1 U365 ( .A(G29GAT), .B(n414), .ZN(n299) );
  XNOR2_X1 U366 ( .A(n299), .B(G197GAT), .ZN(n300) );
  XOR2_X1 U367 ( .A(n301), .B(n300), .Z(n305) );
  XNOR2_X1 U368 ( .A(G50GAT), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U369 ( .A(n302), .B(KEYINPUT8), .ZN(n440) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(G43GAT), .ZN(n303) );
  XNOR2_X1 U371 ( .A(n303), .B(G15GAT), .ZN(n356) );
  XNOR2_X1 U372 ( .A(n440), .B(n356), .ZN(n304) );
  XNOR2_X1 U373 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U374 ( .A(n369), .B(n306), .Z(n308) );
  NAND2_X1 U375 ( .A1(G229GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U376 ( .A(n308), .B(n307), .ZN(n576) );
  XNOR2_X1 U377 ( .A(G99GAT), .B(G71GAT), .ZN(n309) );
  XNOR2_X1 U378 ( .A(n309), .B(G176GAT), .ZN(n358) );
  XNOR2_X1 U379 ( .A(G85GAT), .B(G57GAT), .ZN(n310) );
  XNOR2_X1 U380 ( .A(n310), .B(G120GAT), .ZN(n334) );
  AND2_X1 U381 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XOR2_X1 U382 ( .A(n358), .B(n313), .Z(n315) );
  XOR2_X1 U383 ( .A(KEYINPUT13), .B(KEYINPUT68), .Z(n415) );
  XOR2_X1 U384 ( .A(G92GAT), .B(G64GAT), .Z(n371) );
  XNOR2_X1 U385 ( .A(n415), .B(n371), .ZN(n314) );
  XNOR2_X1 U386 ( .A(n315), .B(n314), .ZN(n323) );
  XNOR2_X1 U387 ( .A(G106GAT), .B(G78GAT), .ZN(n317) );
  XOR2_X1 U388 ( .A(KEYINPUT69), .B(G204GAT), .Z(n318) );
  XOR2_X1 U389 ( .A(KEYINPUT33), .B(KEYINPUT70), .Z(n321) );
  XNOR2_X1 U390 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n320) );
  XOR2_X1 U391 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n324) );
  XNOR2_X1 U392 ( .A(n459), .B(n324), .ZN(n464) );
  XNOR2_X1 U393 ( .A(n464), .B(KEYINPUT107), .ZN(n566) );
  NOR2_X1 U394 ( .A1(n576), .A2(n566), .ZN(n515) );
  XOR2_X1 U395 ( .A(G155GAT), .B(G141GAT), .Z(n326) );
  XNOR2_X1 U396 ( .A(KEYINPUT89), .B(KEYINPUT2), .ZN(n325) );
  XNOR2_X1 U397 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U398 ( .A(KEYINPUT3), .B(n327), .ZN(n391) );
  XOR2_X1 U399 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n329) );
  XNOR2_X1 U400 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n328) );
  XNOR2_X1 U401 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U402 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n331) );
  XNOR2_X1 U403 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n330) );
  XNOR2_X1 U404 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U405 ( .A(n333), .B(n332), .Z(n344) );
  XOR2_X1 U406 ( .A(n334), .B(KEYINPUT93), .Z(n336) );
  NAND2_X1 U407 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U408 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U409 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n338) );
  XNOR2_X1 U410 ( .A(G134GAT), .B(G127GAT), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n338), .B(n337), .ZN(n353) );
  XOR2_X1 U412 ( .A(n353), .B(G113GAT), .Z(n340) );
  XOR2_X1 U413 ( .A(G29GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U414 ( .A(n437), .B(G148GAT), .ZN(n339) );
  XNOR2_X1 U415 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U416 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U417 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U418 ( .A(n391), .B(n345), .Z(n406) );
  XOR2_X1 U419 ( .A(G169GAT), .B(KEYINPUT82), .Z(n347) );
  XNOR2_X1 U420 ( .A(G183GAT), .B(KEYINPUT81), .ZN(n346) );
  XNOR2_X1 U421 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U422 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n349) );
  XNOR2_X1 U423 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n348) );
  XNOR2_X1 U424 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U425 ( .A(n351), .B(n350), .Z(n375) );
  INV_X1 U426 ( .A(n375), .ZN(n352) );
  XOR2_X1 U427 ( .A(n353), .B(n352), .Z(n362) );
  XOR2_X1 U428 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n355) );
  NAND2_X1 U429 ( .A1(G227GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U430 ( .A(n355), .B(n354), .ZN(n357) );
  XOR2_X1 U431 ( .A(n357), .B(n356), .Z(n360) );
  XNOR2_X1 U432 ( .A(G120GAT), .B(n358), .ZN(n359) );
  XNOR2_X1 U433 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U434 ( .A(n362), .B(n361), .Z(n531) );
  XNOR2_X1 U435 ( .A(n363), .B(KEYINPUT87), .ZN(n364) );
  XOR2_X1 U436 ( .A(n364), .B(KEYINPUT21), .Z(n366) );
  XNOR2_X1 U437 ( .A(G218GAT), .B(G211GAT), .ZN(n365) );
  XNOR2_X1 U438 ( .A(n366), .B(n365), .ZN(n388) );
  XOR2_X1 U439 ( .A(G176GAT), .B(G204GAT), .Z(n368) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U441 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U442 ( .A(n370), .B(n369), .Z(n373) );
  XNOR2_X1 U443 ( .A(KEYINPUT74), .B(n371), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U445 ( .A(n388), .B(n374), .ZN(n376) );
  XOR2_X1 U446 ( .A(n376), .B(n375), .Z(n520) );
  INV_X1 U447 ( .A(n520), .ZN(n529) );
  NAND2_X1 U448 ( .A1(n531), .A2(n529), .ZN(n394) );
  XOR2_X1 U449 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n378) );
  XNOR2_X1 U450 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n377) );
  XNOR2_X1 U451 ( .A(n378), .B(n377), .ZN(n385) );
  XOR2_X1 U452 ( .A(KEYINPUT85), .B(G22GAT), .Z(n380) );
  XNOR2_X1 U453 ( .A(G162GAT), .B(G50GAT), .ZN(n379) );
  XNOR2_X1 U454 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U455 ( .A(KEYINPUT23), .B(n381), .Z(n383) );
  NAND2_X1 U456 ( .A1(G228GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U457 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U458 ( .A(n385), .B(n384), .Z(n390) );
  INV_X1 U459 ( .A(n386), .ZN(n387) );
  XOR2_X1 U460 ( .A(n388), .B(n387), .Z(n389) );
  XNOR2_X1 U461 ( .A(n390), .B(n389), .ZN(n393) );
  INV_X1 U462 ( .A(n391), .ZN(n392) );
  INV_X1 U463 ( .A(n477), .ZN(n404) );
  NAND2_X1 U464 ( .A1(n394), .A2(n404), .ZN(n397) );
  XOR2_X1 U465 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n395) );
  XOR2_X1 U466 ( .A(KEYINPUT27), .B(n529), .Z(n407) );
  XNOR2_X1 U467 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n399) );
  INV_X1 U468 ( .A(n531), .ZN(n536) );
  NAND2_X1 U469 ( .A1(n477), .A2(n536), .ZN(n398) );
  NOR2_X1 U470 ( .A1(n407), .A2(n575), .ZN(n400) );
  NOR2_X1 U471 ( .A1(n401), .A2(n400), .ZN(n402) );
  NOR2_X1 U472 ( .A1(n406), .A2(n402), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n403), .B(KEYINPUT99), .ZN(n410) );
  XOR2_X1 U474 ( .A(KEYINPUT84), .B(n536), .Z(n405) );
  NOR2_X1 U475 ( .A1(n512), .A2(n405), .ZN(n408) );
  XOR2_X1 U476 ( .A(KEYINPUT95), .B(n406), .Z(n527) );
  INV_X1 U477 ( .A(n527), .ZN(n516) );
  NOR2_X1 U478 ( .A1(n516), .A2(n407), .ZN(n535) );
  NAND2_X1 U479 ( .A1(n408), .A2(n535), .ZN(n409) );
  NAND2_X1 U480 ( .A1(n410), .A2(n409), .ZN(n411) );
  XOR2_X1 U481 ( .A(KEYINPUT100), .B(n411), .Z(n495) );
  XOR2_X1 U482 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n413) );
  XNOR2_X1 U483 ( .A(G127GAT), .B(KEYINPUT14), .ZN(n412) );
  XNOR2_X1 U484 ( .A(n413), .B(n412), .ZN(n419) );
  XOR2_X1 U485 ( .A(G183GAT), .B(G211GAT), .Z(n417) );
  XNOR2_X1 U486 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U487 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U488 ( .A(n419), .B(n418), .Z(n421) );
  NAND2_X1 U489 ( .A1(G231GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U491 ( .A(G8GAT), .B(G64GAT), .Z(n423) );
  XNOR2_X1 U492 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n422) );
  XNOR2_X1 U493 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U494 ( .A(n425), .B(n424), .Z(n433) );
  XOR2_X1 U495 ( .A(KEYINPUT78), .B(KEYINPUT76), .Z(n427) );
  XNOR2_X1 U496 ( .A(G155GAT), .B(KEYINPUT77), .ZN(n426) );
  XNOR2_X1 U497 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U498 ( .A(KEYINPUT75), .B(G15GAT), .Z(n429) );
  XNOR2_X1 U499 ( .A(G78GAT), .B(G71GAT), .ZN(n428) );
  XNOR2_X1 U500 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U501 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U502 ( .A(n433), .B(n432), .Z(n571) );
  INV_X1 U503 ( .A(n571), .ZN(n584) );
  XNOR2_X1 U504 ( .A(n434), .B(KEYINPUT104), .ZN(n451) );
  XNOR2_X1 U505 ( .A(G134GAT), .B(G218GAT), .ZN(n435) );
  XNOR2_X1 U506 ( .A(n295), .B(n435), .ZN(n436) );
  NAND2_X1 U507 ( .A1(G232GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U508 ( .A(n296), .B(n438), .ZN(n439) );
  XNOR2_X1 U509 ( .A(n439), .B(G92GAT), .ZN(n442) );
  XOR2_X1 U510 ( .A(n440), .B(G99GAT), .Z(n441) );
  XNOR2_X1 U511 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U512 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n444) );
  XNOR2_X1 U513 ( .A(G85GAT), .B(G43GAT), .ZN(n443) );
  XNOR2_X1 U514 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U515 ( .A(G106GAT), .B(G190GAT), .Z(n446) );
  XNOR2_X1 U516 ( .A(KEYINPUT66), .B(KEYINPUT73), .ZN(n445) );
  XNOR2_X1 U517 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U518 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U519 ( .A(KEYINPUT36), .B(n548), .Z(n586) );
  NAND2_X1 U520 ( .A1(n451), .A2(n586), .ZN(n454) );
  AND2_X1 U521 ( .A1(n515), .A2(n487), .ZN(n455) );
  NAND2_X1 U522 ( .A1(n532), .A2(n512), .ZN(n458) );
  XOR2_X1 U523 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n456) );
  XNOR2_X1 U524 ( .A(n458), .B(n457), .ZN(G1339GAT) );
  NAND2_X1 U525 ( .A1(n584), .A2(n586), .ZN(n460) );
  XNOR2_X1 U526 ( .A(n460), .B(KEYINPUT113), .ZN(n461) );
  XNOR2_X1 U527 ( .A(n461), .B(KEYINPUT45), .ZN(n462) );
  XNOR2_X1 U528 ( .A(n576), .B(KEYINPUT67), .ZN(n564) );
  NAND2_X1 U529 ( .A1(n462), .A2(n564), .ZN(n463) );
  NOR2_X1 U530 ( .A1(n459), .A2(n463), .ZN(n471) );
  NAND2_X1 U531 ( .A1(n464), .A2(n576), .ZN(n466) );
  INV_X1 U532 ( .A(n548), .ZN(n562) );
  NOR2_X1 U533 ( .A1(n584), .A2(n562), .ZN(n467) );
  NAND2_X1 U534 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U535 ( .A(n469), .B(KEYINPUT47), .ZN(n470) );
  OR2_X1 U536 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U537 ( .A1(n534), .A2(n529), .ZN(n474) );
  XOR2_X1 U538 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n473) );
  XNOR2_X1 U539 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U540 ( .A1(n475), .A2(n527), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n476), .B(KEYINPUT65), .ZN(n574) );
  NOR2_X1 U542 ( .A1(n477), .A2(n574), .ZN(n480) );
  INV_X1 U543 ( .A(KEYINPUT55), .ZN(n478) );
  XNOR2_X1 U544 ( .A(n480), .B(n479), .ZN(n481) );
  NAND2_X1 U545 ( .A1(n481), .A2(n531), .ZN(n570) );
  NOR2_X1 U546 ( .A1(n548), .A2(n570), .ZN(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n483) );
  INV_X1 U548 ( .A(G190GAT), .ZN(n482) );
  XOR2_X1 U549 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n489) );
  NOR2_X1 U550 ( .A1(n459), .A2(n564), .ZN(n486) );
  XNOR2_X1 U551 ( .A(KEYINPUT72), .B(n486), .ZN(n497) );
  NAND2_X1 U552 ( .A1(n487), .A2(n497), .ZN(n488) );
  NAND2_X1 U553 ( .A1(n527), .A2(n511), .ZN(n492) );
  XOR2_X1 U554 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n494) );
  NAND2_X1 U555 ( .A1(n584), .A2(n548), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(n496) );
  NOR2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n514) );
  NAND2_X1 U558 ( .A1(n514), .A2(n497), .ZN(n505) );
  NOR2_X1 U559 ( .A1(n516), .A2(n505), .ZN(n498) );
  XOR2_X1 U560 ( .A(KEYINPUT34), .B(n498), .Z(n499) );
  XNOR2_X1 U561 ( .A(G1GAT), .B(n499), .ZN(G1324GAT) );
  NOR2_X1 U562 ( .A1(n520), .A2(n505), .ZN(n500) );
  XOR2_X1 U563 ( .A(G8GAT), .B(n500), .Z(G1325GAT) );
  NOR2_X1 U564 ( .A1(n505), .A2(n536), .ZN(n504) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n502) );
  XNOR2_X1 U566 ( .A(G15GAT), .B(KEYINPUT102), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1326GAT) );
  INV_X1 U569 ( .A(n512), .ZN(n538) );
  NOR2_X1 U570 ( .A1(n538), .A2(n505), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1327GAT) );
  NAND2_X1 U573 ( .A1(n511), .A2(n529), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U575 ( .A1(n531), .A2(n511), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(KEYINPUT40), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G43GAT), .B(n510), .ZN(G1330GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U580 ( .A1(n515), .A2(n514), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n516), .A2(n524), .ZN(n518) );
  XNOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT42), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U584 ( .A(G57GAT), .B(n519), .Z(G1332GAT) );
  NOR2_X1 U585 ( .A1(n520), .A2(n524), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G64GAT), .B(KEYINPUT109), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n522), .B(n521), .ZN(G1333GAT) );
  NOR2_X1 U588 ( .A1(n536), .A2(n524), .ZN(n523) );
  XOR2_X1 U589 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U590 ( .A1(n538), .A2(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n532), .ZN(n528) );
  XNOR2_X1 U594 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n533), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n552) );
  NOR2_X1 U600 ( .A1(n536), .A2(n552), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(n547) );
  NOR2_X1 U602 ( .A1(n564), .A2(n547), .ZN(n539) );
  XOR2_X1 U603 ( .A(n539), .B(KEYINPUT114), .Z(n540) );
  XNOR2_X1 U604 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  NOR2_X1 U605 ( .A1(n566), .A2(n547), .ZN(n542) );
  XNOR2_X1 U606 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  NOR2_X1 U609 ( .A1(n571), .A2(n547), .ZN(n545) );
  XNOR2_X1 U610 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  NOR2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n550) );
  XNOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U616 ( .A(G134GAT), .B(n551), .Z(G1343GAT) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n554) );
  NOR2_X1 U618 ( .A1(n575), .A2(n552), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n576), .A2(n561), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n556) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U624 ( .A(KEYINPUT52), .B(n557), .Z(n559) );
  NAND2_X1 U625 ( .A1(n561), .A2(n464), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n584), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U631 ( .A1(n564), .A2(n570), .ZN(n565) );
  XOR2_X1 U632 ( .A(G169GAT), .B(n565), .Z(G1348GAT) );
  XNOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G176GAT), .ZN(G1349GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n578) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n587) );
  NAND2_X1 U641 ( .A1(n587), .A2(n576), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(n579), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n587), .A2(n459), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

