

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n540), .A2(n539), .ZN(G160) );
  OR2_X2 U550 ( .A1(G164), .A2(G1384), .ZN(n598) );
  XNOR2_X2 U551 ( .A(n531), .B(KEYINPUT89), .ZN(G164) );
  NOR2_X1 U552 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U553 ( .A(n691), .ZN(n676) );
  AND2_X2 U554 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  INV_X1 U555 ( .A(n536), .ZN(n518) );
  INV_X2 U556 ( .A(n518), .ZN(n519) );
  NOR2_X1 U557 ( .A1(n521), .A2(n520), .ZN(n536) );
  XNOR2_X1 U558 ( .A(KEYINPUT23), .B(KEYINPUT67), .ZN(n532) );
  INV_X1 U559 ( .A(KEYINPUT31), .ZN(n642) );
  XNOR2_X1 U560 ( .A(n642), .B(KEYINPUT100), .ZN(n643) );
  NOR2_X1 U561 ( .A1(G1966), .A2(n716), .ZN(n711) );
  NAND2_X1 U562 ( .A1(n631), .A2(n630), .ZN(n664) );
  AND2_X1 U563 ( .A1(n713), .A2(n712), .ZN(n722) );
  NAND2_X1 U564 ( .A1(n888), .A2(G138), .ZN(n524) );
  INV_X1 U565 ( .A(KEYINPUT17), .ZN(n522) );
  AND2_X1 U566 ( .A1(n521), .A2(n520), .ZN(n889) );
  NOR2_X1 U567 ( .A1(G651), .A2(n578), .ZN(n795) );
  XNOR2_X1 U568 ( .A(n533), .B(n532), .ZN(n535) );
  INV_X1 U569 ( .A(G2105), .ZN(n521) );
  XNOR2_X1 U570 ( .A(G2104), .B(KEYINPUT66), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n889), .A2(G102), .ZN(n530) );
  NAND2_X1 U572 ( .A1(G126), .A2(n519), .ZN(n525) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XNOR2_X2 U574 ( .A(n523), .B(n522), .ZN(n888) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n528) );
  NAND2_X1 U576 ( .A1(G114), .A2(n892), .ZN(n526) );
  XOR2_X1 U577 ( .A(KEYINPUT88), .B(n526), .Z(n527) );
  NOR2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G101), .A2(n889), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G137), .A2(n888), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n540) );
  NAND2_X1 U583 ( .A1(G113), .A2(n892), .ZN(n538) );
  NAND2_X1 U584 ( .A1(G125), .A2(n519), .ZN(n537) );
  NAND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n539) );
  INV_X1 U586 ( .A(G651), .ZN(n547) );
  NOR2_X1 U587 ( .A1(G543), .A2(n547), .ZN(n541) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n541), .Z(n799) );
  NAND2_X1 U589 ( .A1(G63), .A2(n799), .ZN(n543) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n578) );
  NAND2_X1 U591 ( .A1(G51), .A2(n795), .ZN(n542) );
  NAND2_X1 U592 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U593 ( .A(KEYINPUT6), .B(n544), .ZN(n552) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n791) );
  NAND2_X1 U595 ( .A1(G89), .A2(n791), .ZN(n545) );
  XNOR2_X1 U596 ( .A(n545), .B(KEYINPUT4), .ZN(n546) );
  XNOR2_X1 U597 ( .A(n546), .B(KEYINPUT74), .ZN(n549) );
  NOR2_X1 U598 ( .A1(n578), .A2(n547), .ZN(n792) );
  NAND2_X1 U599 ( .A1(G76), .A2(n792), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U601 ( .A(n550), .B(KEYINPUT5), .Z(n551) );
  NOR2_X1 U602 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U603 ( .A(KEYINPUT7), .B(n553), .Z(n555) );
  XOR2_X1 U604 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n554) );
  XNOR2_X1 U605 ( .A(n555), .B(n554), .ZN(G168) );
  NAND2_X1 U606 ( .A1(G90), .A2(n791), .ZN(n557) );
  NAND2_X1 U607 ( .A1(G77), .A2(n792), .ZN(n556) );
  NAND2_X1 U608 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U609 ( .A(n558), .B(KEYINPUT9), .ZN(n560) );
  NAND2_X1 U610 ( .A1(G52), .A2(n795), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n560), .A2(n559), .ZN(n563) );
  NAND2_X1 U612 ( .A1(n799), .A2(G64), .ZN(n561) );
  XOR2_X1 U613 ( .A(KEYINPUT68), .B(n561), .Z(n562) );
  NOR2_X1 U614 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U615 ( .A(KEYINPUT69), .B(n564), .Z(G171) );
  NAND2_X1 U616 ( .A1(G91), .A2(n791), .ZN(n566) );
  NAND2_X1 U617 ( .A1(G78), .A2(n792), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U619 ( .A(KEYINPUT70), .B(n567), .Z(n571) );
  NAND2_X1 U620 ( .A1(G65), .A2(n799), .ZN(n569) );
  NAND2_X1 U621 ( .A1(G53), .A2(n795), .ZN(n568) );
  AND2_X1 U622 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U623 ( .A1(n571), .A2(n570), .ZN(G299) );
  NAND2_X1 U624 ( .A1(G88), .A2(n791), .ZN(n573) );
  NAND2_X1 U625 ( .A1(G75), .A2(n792), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U627 ( .A1(G62), .A2(n799), .ZN(n575) );
  NAND2_X1 U628 ( .A1(G50), .A2(n795), .ZN(n574) );
  NAND2_X1 U629 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U630 ( .A1(n577), .A2(n576), .ZN(G166) );
  INV_X1 U631 ( .A(G166), .ZN(G303) );
  XOR2_X1 U632 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U633 ( .A1(G49), .A2(n795), .ZN(n580) );
  NAND2_X1 U634 ( .A1(G87), .A2(n578), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U636 ( .A1(n799), .A2(n581), .ZN(n584) );
  NAND2_X1 U637 ( .A1(G74), .A2(G651), .ZN(n582) );
  XOR2_X1 U638 ( .A(KEYINPUT83), .B(n582), .Z(n583) );
  NAND2_X1 U639 ( .A1(n584), .A2(n583), .ZN(G288) );
  NAND2_X1 U640 ( .A1(G61), .A2(n799), .ZN(n586) );
  NAND2_X1 U641 ( .A1(G86), .A2(n791), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U643 ( .A1(n792), .A2(G73), .ZN(n587) );
  XOR2_X1 U644 ( .A(KEYINPUT2), .B(n587), .Z(n588) );
  NOR2_X1 U645 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U646 ( .A1(n795), .A2(G48), .ZN(n590) );
  NAND2_X1 U647 ( .A1(n591), .A2(n590), .ZN(G305) );
  NAND2_X1 U648 ( .A1(G85), .A2(n791), .ZN(n593) );
  NAND2_X1 U649 ( .A1(G72), .A2(n792), .ZN(n592) );
  NAND2_X1 U650 ( .A1(n593), .A2(n592), .ZN(n597) );
  NAND2_X1 U651 ( .A1(G60), .A2(n799), .ZN(n595) );
  NAND2_X1 U652 ( .A1(G47), .A2(n795), .ZN(n594) );
  NAND2_X1 U653 ( .A1(n595), .A2(n594), .ZN(n596) );
  OR2_X1 U654 ( .A1(n597), .A2(n596), .ZN(G290) );
  NAND2_X1 U655 ( .A1(n598), .A2(KEYINPUT65), .ZN(n601) );
  OR2_X1 U656 ( .A1(G1384), .A2(KEYINPUT65), .ZN(n599) );
  OR2_X1 U657 ( .A1(G164), .A2(n599), .ZN(n600) );
  NAND2_X1 U658 ( .A1(n601), .A2(n600), .ZN(n631) );
  NAND2_X1 U659 ( .A1(G160), .A2(G40), .ZN(n629) );
  NOR2_X1 U660 ( .A1(n631), .A2(n629), .ZN(n758) );
  XNOR2_X1 U661 ( .A(KEYINPUT37), .B(G2067), .ZN(n756) );
  NAND2_X1 U662 ( .A1(G140), .A2(n888), .ZN(n603) );
  NAND2_X1 U663 ( .A1(G104), .A2(n889), .ZN(n602) );
  NAND2_X1 U664 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U665 ( .A(KEYINPUT34), .B(n604), .ZN(n609) );
  NAND2_X1 U666 ( .A1(G116), .A2(n892), .ZN(n606) );
  NAND2_X1 U667 ( .A1(G128), .A2(n519), .ZN(n605) );
  NAND2_X1 U668 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U669 ( .A(KEYINPUT35), .B(n607), .Z(n608) );
  NOR2_X1 U670 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U671 ( .A(KEYINPUT36), .B(n610), .ZN(n885) );
  NOR2_X1 U672 ( .A1(n756), .A2(n885), .ZN(n1009) );
  NAND2_X1 U673 ( .A1(n758), .A2(n1009), .ZN(n754) );
  NAND2_X1 U674 ( .A1(G107), .A2(n892), .ZN(n612) );
  NAND2_X1 U675 ( .A1(G131), .A2(n888), .ZN(n611) );
  NAND2_X1 U676 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U677 ( .A1(n889), .A2(G95), .ZN(n613) );
  XOR2_X1 U678 ( .A(KEYINPUT90), .B(n613), .Z(n614) );
  NOR2_X1 U679 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U680 ( .A1(n519), .A2(G119), .ZN(n616) );
  NAND2_X1 U681 ( .A1(n617), .A2(n616), .ZN(n901) );
  NAND2_X1 U682 ( .A1(G1991), .A2(n901), .ZN(n627) );
  NAND2_X1 U683 ( .A1(G105), .A2(n889), .ZN(n618) );
  XNOR2_X1 U684 ( .A(n618), .B(KEYINPUT38), .ZN(n625) );
  NAND2_X1 U685 ( .A1(G117), .A2(n892), .ZN(n620) );
  NAND2_X1 U686 ( .A1(G129), .A2(n519), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U688 ( .A1(G141), .A2(n888), .ZN(n621) );
  XNOR2_X1 U689 ( .A(KEYINPUT91), .B(n621), .ZN(n622) );
  NOR2_X1 U690 ( .A1(n623), .A2(n622), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n625), .A2(n624), .ZN(n880) );
  NAND2_X1 U692 ( .A1(G1996), .A2(n880), .ZN(n626) );
  NAND2_X1 U693 ( .A1(n627), .A2(n626), .ZN(n1017) );
  NAND2_X1 U694 ( .A1(n758), .A2(n1017), .ZN(n749) );
  NAND2_X1 U695 ( .A1(n754), .A2(n749), .ZN(n628) );
  XNOR2_X1 U696 ( .A(KEYINPUT92), .B(n628), .ZN(n742) );
  INV_X1 U697 ( .A(n629), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n664), .A2(G8), .ZN(n632) );
  XNOR2_X1 U699 ( .A(KEYINPUT93), .B(n632), .ZN(n734) );
  INV_X1 U700 ( .A(n734), .ZN(n716) );
  NOR2_X1 U701 ( .A1(n664), .A2(G2084), .ZN(n633) );
  XOR2_X1 U702 ( .A(n633), .B(KEYINPUT95), .Z(n707) );
  INV_X1 U703 ( .A(n707), .ZN(n634) );
  NAND2_X1 U704 ( .A1(G8), .A2(n634), .ZN(n635) );
  NOR2_X1 U705 ( .A1(n711), .A2(n635), .ZN(n636) );
  XOR2_X1 U706 ( .A(n636), .B(KEYINPUT30), .Z(n637) );
  NOR2_X1 U707 ( .A1(G168), .A2(n637), .ZN(n641) );
  BUF_X2 U708 ( .A(n664), .Z(n691) );
  INV_X1 U709 ( .A(G1961), .ZN(n941) );
  NAND2_X1 U710 ( .A1(n691), .A2(n941), .ZN(n639) );
  XNOR2_X1 U711 ( .A(G2078), .B(KEYINPUT25), .ZN(n982) );
  NAND2_X1 U712 ( .A1(n676), .A2(n982), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n688) );
  NOR2_X1 U714 ( .A1(G171), .A2(n688), .ZN(n640) );
  NOR2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n644) );
  XNOR2_X1 U716 ( .A(n644), .B(n643), .ZN(n706) );
  NAND2_X1 U717 ( .A1(G66), .A2(n799), .ZN(n646) );
  NAND2_X1 U718 ( .A1(G92), .A2(n791), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U720 ( .A1(G79), .A2(n792), .ZN(n648) );
  NAND2_X1 U721 ( .A1(G54), .A2(n795), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n652) );
  XNOR2_X1 U724 ( .A(KEYINPUT73), .B(KEYINPUT15), .ZN(n651) );
  XOR2_X1 U725 ( .A(n652), .B(n651), .Z(n925) );
  NOR2_X1 U726 ( .A1(n676), .A2(G1348), .ZN(n654) );
  NOR2_X1 U727 ( .A1(G2067), .A2(n691), .ZN(n653) );
  NOR2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n671) );
  NAND2_X1 U729 ( .A1(n925), .A2(n671), .ZN(n670) );
  NAND2_X1 U730 ( .A1(G56), .A2(n799), .ZN(n655) );
  XOR2_X1 U731 ( .A(KEYINPUT14), .B(n655), .Z(n661) );
  NAND2_X1 U732 ( .A1(n791), .A2(G81), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n656), .B(KEYINPUT12), .ZN(n658) );
  NAND2_X1 U734 ( .A1(G68), .A2(n792), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U736 ( .A(KEYINPUT13), .B(n659), .Z(n660) );
  NOR2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n795), .A2(G43), .ZN(n662) );
  NAND2_X1 U739 ( .A1(n663), .A2(n662), .ZN(n926) );
  INV_X1 U740 ( .A(G1996), .ZN(n840) );
  NOR2_X1 U741 ( .A1(n664), .A2(n840), .ZN(n665) );
  XOR2_X1 U742 ( .A(n665), .B(KEYINPUT26), .Z(n667) );
  NAND2_X1 U743 ( .A1(n691), .A2(G1341), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U745 ( .A1(n926), .A2(n668), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n670), .A2(n669), .ZN(n673) );
  OR2_X1 U747 ( .A1(n671), .A2(n925), .ZN(n672) );
  NAND2_X1 U748 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U749 ( .A(KEYINPUT97), .B(n674), .ZN(n680) );
  NAND2_X1 U750 ( .A1(n676), .A2(G2072), .ZN(n675) );
  XNOR2_X1 U751 ( .A(n675), .B(KEYINPUT27), .ZN(n678) );
  XOR2_X1 U752 ( .A(G1956), .B(KEYINPUT96), .Z(n948) );
  NOR2_X1 U753 ( .A1(n676), .A2(n948), .ZN(n677) );
  NOR2_X1 U754 ( .A1(n678), .A2(n677), .ZN(n681) );
  INV_X1 U755 ( .A(G299), .ZN(n931) );
  NAND2_X1 U756 ( .A1(n681), .A2(n931), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n680), .A2(n679), .ZN(n684) );
  NOR2_X1 U758 ( .A1(n681), .A2(n931), .ZN(n682) );
  XOR2_X1 U759 ( .A(n682), .B(KEYINPUT28), .Z(n683) );
  NAND2_X1 U760 ( .A1(n684), .A2(n683), .ZN(n687) );
  XNOR2_X1 U761 ( .A(KEYINPUT29), .B(KEYINPUT98), .ZN(n685) );
  XNOR2_X1 U762 ( .A(n685), .B(KEYINPUT99), .ZN(n686) );
  XNOR2_X1 U763 ( .A(n687), .B(n686), .ZN(n690) );
  NAND2_X1 U764 ( .A1(n688), .A2(G171), .ZN(n689) );
  NAND2_X1 U765 ( .A1(n690), .A2(n689), .ZN(n705) );
  INV_X1 U766 ( .A(G8), .ZN(n697) );
  NOR2_X1 U767 ( .A1(G1971), .A2(n716), .ZN(n693) );
  NOR2_X1 U768 ( .A1(G2090), .A2(n691), .ZN(n692) );
  NOR2_X1 U769 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U770 ( .A(KEYINPUT101), .B(n694), .Z(n695) );
  NAND2_X1 U771 ( .A1(n695), .A2(G303), .ZN(n696) );
  OR2_X1 U772 ( .A1(n697), .A2(n696), .ZN(n699) );
  AND2_X1 U773 ( .A1(n705), .A2(n699), .ZN(n698) );
  NAND2_X1 U774 ( .A1(n706), .A2(n698), .ZN(n703) );
  INV_X1 U775 ( .A(n699), .ZN(n701) );
  AND2_X1 U776 ( .A1(G286), .A2(G8), .ZN(n700) );
  OR2_X1 U777 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U778 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U779 ( .A(n704), .B(KEYINPUT32), .ZN(n713) );
  NAND2_X1 U780 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U781 ( .A1(G8), .A2(n707), .ZN(n708) );
  NAND2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n710) );
  OR2_X1 U783 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U784 ( .A1(G1976), .A2(G288), .ZN(n733) );
  NOR2_X1 U785 ( .A1(G1971), .A2(G303), .ZN(n714) );
  NOR2_X1 U786 ( .A1(n733), .A2(n714), .ZN(n935) );
  INV_X1 U787 ( .A(n935), .ZN(n715) );
  NOR2_X1 U788 ( .A1(n722), .A2(n715), .ZN(n718) );
  NAND2_X1 U789 ( .A1(G1976), .A2(G288), .ZN(n930) );
  NAND2_X1 U790 ( .A1(n734), .A2(n930), .ZN(n717) );
  NOR2_X1 U791 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U792 ( .A(n719), .B(KEYINPUT64), .ZN(n729) );
  NAND2_X1 U793 ( .A1(G166), .A2(G8), .ZN(n720) );
  NOR2_X1 U794 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U795 ( .A1(n722), .A2(n721), .ZN(n723) );
  OR2_X1 U796 ( .A1(n723), .A2(n734), .ZN(n731) );
  NOR2_X1 U797 ( .A1(G1981), .A2(G305), .ZN(n724) );
  XNOR2_X1 U798 ( .A(n724), .B(KEYINPUT94), .ZN(n725) );
  XNOR2_X1 U799 ( .A(n725), .B(KEYINPUT24), .ZN(n726) );
  AND2_X1 U800 ( .A1(n726), .A2(n734), .ZN(n730) );
  NOR2_X1 U801 ( .A1(n730), .A2(KEYINPUT33), .ZN(n727) );
  NAND2_X1 U802 ( .A1(n731), .A2(n727), .ZN(n728) );
  OR2_X1 U803 ( .A1(n729), .A2(n728), .ZN(n740) );
  INV_X1 U804 ( .A(n730), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n732), .A2(n731), .ZN(n738) );
  XNOR2_X1 U806 ( .A(G1981), .B(G305), .ZN(n923) );
  AND2_X1 U807 ( .A1(n733), .A2(KEYINPUT33), .ZN(n735) );
  AND2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U809 ( .A1(n923), .A2(n736), .ZN(n737) );
  OR2_X1 U810 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U811 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U812 ( .A(n743), .B(KEYINPUT102), .ZN(n745) );
  XNOR2_X1 U813 ( .A(G1986), .B(G290), .ZN(n937) );
  NAND2_X1 U814 ( .A1(n937), .A2(n758), .ZN(n744) );
  NAND2_X1 U815 ( .A1(n745), .A2(n744), .ZN(n761) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n880), .ZN(n746) );
  XOR2_X1 U817 ( .A(KEYINPUT103), .B(n746), .Z(n1014) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n901), .ZN(n1008) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n747) );
  NOR2_X1 U820 ( .A1(n1008), .A2(n747), .ZN(n748) );
  XOR2_X1 U821 ( .A(KEYINPUT104), .B(n748), .Z(n750) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U823 ( .A(KEYINPUT105), .B(n751), .ZN(n752) );
  NOR2_X1 U824 ( .A1(n1014), .A2(n752), .ZN(n753) );
  XNOR2_X1 U825 ( .A(n753), .B(KEYINPUT39), .ZN(n755) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n757) );
  NAND2_X1 U827 ( .A1(n756), .A2(n885), .ZN(n1016) );
  NAND2_X1 U828 ( .A1(n757), .A2(n1016), .ZN(n759) );
  NAND2_X1 U829 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U831 ( .A(n762), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U832 ( .A(G171), .ZN(G301) );
  AND2_X1 U833 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U834 ( .A(G57), .ZN(G237) );
  INV_X1 U835 ( .A(G69), .ZN(G235) );
  INV_X1 U836 ( .A(G108), .ZN(G238) );
  INV_X1 U837 ( .A(G120), .ZN(G236) );
  INV_X1 U838 ( .A(G132), .ZN(G219) );
  INV_X1 U839 ( .A(G82), .ZN(G220) );
  XOR2_X1 U840 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n764) );
  NAND2_X1 U841 ( .A1(G7), .A2(G661), .ZN(n763) );
  XOR2_X1 U842 ( .A(n764), .B(n763), .Z(n831) );
  AND2_X1 U843 ( .A1(G567), .A2(n831), .ZN(n765) );
  XNOR2_X1 U844 ( .A(n765), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U845 ( .A(G860), .ZN(n790) );
  NOR2_X1 U846 ( .A1(n926), .A2(n790), .ZN(n766) );
  XOR2_X1 U847 ( .A(KEYINPUT72), .B(n766), .Z(G153) );
  NAND2_X1 U848 ( .A1(G868), .A2(G301), .ZN(n768) );
  INV_X1 U849 ( .A(G868), .ZN(n811) );
  NAND2_X1 U850 ( .A1(n925), .A2(n811), .ZN(n767) );
  NAND2_X1 U851 ( .A1(n768), .A2(n767), .ZN(G284) );
  NAND2_X1 U852 ( .A1(G868), .A2(G286), .ZN(n770) );
  NAND2_X1 U853 ( .A1(G299), .A2(n811), .ZN(n769) );
  NAND2_X1 U854 ( .A1(n770), .A2(n769), .ZN(G297) );
  NAND2_X1 U855 ( .A1(n790), .A2(G559), .ZN(n771) );
  INV_X1 U856 ( .A(n925), .ZN(n859) );
  NAND2_X1 U857 ( .A1(n771), .A2(n859), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U859 ( .A1(G559), .A2(n811), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n859), .A2(n773), .ZN(n774) );
  XNOR2_X1 U861 ( .A(n774), .B(KEYINPUT77), .ZN(n776) );
  NOR2_X1 U862 ( .A1(n926), .A2(G868), .ZN(n775) );
  NOR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(G282) );
  XNOR2_X1 U864 ( .A(G2100), .B(KEYINPUT81), .ZN(n788) );
  NAND2_X1 U865 ( .A1(n888), .A2(G135), .ZN(n777) );
  XNOR2_X1 U866 ( .A(KEYINPUT78), .B(n777), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n519), .A2(G123), .ZN(n778) );
  XNOR2_X1 U868 ( .A(KEYINPUT18), .B(n778), .ZN(n779) );
  NAND2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(KEYINPUT79), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G111), .A2(n892), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n889), .A2(G99), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT80), .B(n784), .Z(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n1007) );
  XNOR2_X1 U876 ( .A(n1007), .B(G2096), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(G156) );
  NAND2_X1 U878 ( .A1(G559), .A2(n859), .ZN(n789) );
  XOR2_X1 U879 ( .A(n926), .B(n789), .Z(n808) );
  NAND2_X1 U880 ( .A1(n790), .A2(n808), .ZN(n802) );
  NAND2_X1 U881 ( .A1(G93), .A2(n791), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G80), .A2(n792), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n795), .A2(G55), .ZN(n796) );
  XOR2_X1 U885 ( .A(KEYINPUT82), .B(n796), .Z(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n799), .A2(G67), .ZN(n800) );
  NAND2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n810) );
  XNOR2_X1 U889 ( .A(n802), .B(n810), .ZN(G145) );
  XOR2_X1 U890 ( .A(G303), .B(KEYINPUT19), .Z(n807) );
  XOR2_X1 U891 ( .A(G299), .B(G305), .Z(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(n810), .ZN(n804) );
  XNOR2_X1 U893 ( .A(n804), .B(G290), .ZN(n805) );
  XNOR2_X1 U894 ( .A(n805), .B(G288), .ZN(n806) );
  XNOR2_X1 U895 ( .A(n807), .B(n806), .ZN(n858) );
  XNOR2_X1 U896 ( .A(n808), .B(n858), .ZN(n809) );
  NAND2_X1 U897 ( .A1(n809), .A2(G868), .ZN(n813) );
  NAND2_X1 U898 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U899 ( .A1(n813), .A2(n812), .ZN(G295) );
  XOR2_X1 U900 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n815) );
  NAND2_X1 U901 ( .A1(G2078), .A2(G2084), .ZN(n814) );
  XNOR2_X1 U902 ( .A(n815), .B(n814), .ZN(n816) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n816), .ZN(n817) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n817), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n818), .A2(G2072), .ZN(n819) );
  XOR2_X1 U906 ( .A(KEYINPUT85), .B(n819), .Z(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U908 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U909 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U910 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U911 ( .A1(G96), .A2(n822), .ZN(n835) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n835), .ZN(n823) );
  XOR2_X1 U913 ( .A(KEYINPUT86), .B(n823), .Z(n828) );
  NOR2_X1 U914 ( .A1(G236), .A2(G238), .ZN(n825) );
  NOR2_X1 U915 ( .A1(G235), .A2(G237), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n826) );
  XOR2_X1 U917 ( .A(KEYINPUT87), .B(n826), .Z(n836) );
  AND2_X1 U918 ( .A1(n836), .A2(G567), .ZN(n827) );
  NOR2_X1 U919 ( .A1(n828), .A2(n827), .ZN(G319) );
  INV_X1 U920 ( .A(G319), .ZN(n830) );
  NAND2_X1 U921 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n834) );
  NAND2_X1 U923 ( .A1(n834), .A2(G36), .ZN(G176) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  INV_X1 U925 ( .A(n831), .ZN(G223) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U927 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U929 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U933 ( .A(KEYINPUT106), .B(n837), .Z(G261) );
  INV_X1 U934 ( .A(G261), .ZN(G325) );
  XNOR2_X1 U935 ( .A(G1966), .B(KEYINPUT41), .ZN(n848) );
  XOR2_X1 U936 ( .A(G1981), .B(G1956), .Z(n839) );
  XOR2_X1 U937 ( .A(G1986), .B(n941), .Z(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n844) );
  XOR2_X1 U939 ( .A(G1976), .B(G1971), .Z(n842) );
  XOR2_X1 U940 ( .A(n840), .B(G1991), .Z(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U943 ( .A(KEYINPUT108), .B(G2474), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2090), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2078), .B(G2072), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n851), .B(G2096), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2084), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U952 ( .A(G2100), .B(KEYINPUT43), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT107), .B(G2678), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(G227) );
  XNOR2_X1 U956 ( .A(n926), .B(n858), .ZN(n861) );
  XOR2_X1 U957 ( .A(G301), .B(n859), .Z(n860) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n862), .B(G286), .ZN(n863) );
  NOR2_X1 U960 ( .A1(G37), .A2(n863), .ZN(G397) );
  NAND2_X1 U961 ( .A1(G112), .A2(n892), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G136), .A2(n888), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n870) );
  NAND2_X1 U964 ( .A1(n519), .A2(G124), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U966 ( .A1(G100), .A2(n889), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U968 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U969 ( .A1(G118), .A2(n892), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G130), .A2(n519), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n879) );
  XNOR2_X1 U972 ( .A(KEYINPUT110), .B(KEYINPUT45), .ZN(n877) );
  NAND2_X1 U973 ( .A1(n889), .A2(G106), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n888), .A2(G142), .ZN(n873) );
  XOR2_X1 U975 ( .A(KEYINPUT109), .B(n873), .Z(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n877), .B(n876), .Z(n878) );
  NOR2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n884) );
  XNOR2_X1 U979 ( .A(n880), .B(G162), .ZN(n882) );
  XNOR2_X1 U980 ( .A(G164), .B(G160), .ZN(n881) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n885), .B(n1007), .ZN(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n903) );
  XOR2_X1 U985 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n899) );
  NAND2_X1 U986 ( .A1(G139), .A2(n888), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G103), .A2(n889), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n897) );
  NAND2_X1 U989 ( .A1(G115), .A2(n892), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G127), .A2(n519), .ZN(n893) );
  NAND2_X1 U991 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U992 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n999) );
  XNOR2_X1 U994 ( .A(n999), .B(KEYINPUT111), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(n905) );
  XNOR2_X1 U999 ( .A(KEYINPUT112), .B(n905), .ZN(G395) );
  XOR2_X1 U1000 ( .A(G2451), .B(G2430), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2443), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n913) );
  XOR2_X1 U1003 ( .A(G2435), .B(G2454), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G2446), .B(G2427), .Z(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1009 ( .A1(G14), .A2(n914), .ZN(n920) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G397), .A2(G395), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(n920), .ZN(G401) );
  XNOR2_X1 U1018 ( .A(KEYINPUT56), .B(KEYINPUT121), .ZN(n921) );
  XOR2_X1 U1019 ( .A(G16), .B(n921), .Z(n947) );
  XOR2_X1 U1020 ( .A(G168), .B(G1966), .Z(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1022 ( .A(KEYINPUT57), .B(n924), .Z(n945) );
  XNOR2_X1 U1023 ( .A(G1348), .B(n925), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n926), .B(G1341), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n940) );
  NAND2_X1 U1026 ( .A1(G1971), .A2(G303), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1028 ( .A(G1956), .B(n931), .Z(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(n938), .B(KEYINPUT122), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n943) );
  XOR2_X1 U1034 ( .A(n941), .B(G301), .Z(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1037 ( .A1(n947), .A2(n946), .ZN(n974) );
  INV_X1 U1038 ( .A(G16), .ZN(n972) );
  XOR2_X1 U1039 ( .A(G5), .B(G1961), .Z(n962) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G21), .ZN(n960) );
  XNOR2_X1 U1041 ( .A(n948), .B(G20), .ZN(n956) );
  XNOR2_X1 U1042 ( .A(KEYINPUT59), .B(G1348), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n949), .B(G4), .ZN(n951) );
  XOR2_X1 U1044 ( .A(G1341), .B(G19), .Z(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1046 ( .A(KEYINPUT123), .B(G1981), .Z(n952) );
  XNOR2_X1 U1047 ( .A(G6), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(n957), .B(KEYINPUT60), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(KEYINPUT124), .B(n958), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1053 ( .A1(n962), .A2(n961), .ZN(n969) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n966) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n965) );
  NAND2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n967), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(KEYINPUT61), .B(n970), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(KEYINPUT125), .B(n975), .ZN(n976) );
  NAND2_X1 U1065 ( .A1(n976), .A2(G11), .ZN(n1030) );
  XOR2_X1 U1066 ( .A(KEYINPUT119), .B(G34), .Z(n978) );
  XNOR2_X1 U1067 ( .A(G2084), .B(KEYINPUT54), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n978), .B(n977), .ZN(n995) );
  XNOR2_X1 U1069 ( .A(G2090), .B(G35), .ZN(n992) );
  XOR2_X1 U1070 ( .A(G1991), .B(G25), .Z(n979) );
  NAND2_X1 U1071 ( .A1(n979), .A2(G28), .ZN(n988) );
  XNOR2_X1 U1072 ( .A(G2067), .B(G26), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G33), .B(G2072), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n986) );
  XOR2_X1 U1075 ( .A(n982), .B(G27), .Z(n984) );
  XNOR2_X1 U1076 ( .A(G1996), .B(G32), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1080 ( .A(KEYINPUT53), .B(n989), .Z(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(KEYINPUT117), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1083 ( .A(KEYINPUT118), .B(n993), .Z(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1085 ( .A(KEYINPUT120), .B(n996), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(G29), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1087 ( .A(n998), .B(KEYINPUT55), .ZN(n1028) );
  XOR2_X1 U1088 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n1004) );
  XOR2_X1 U1089 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1090 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT50), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1004), .B(n1003), .ZN(n1024) );
  XNOR2_X1 U1094 ( .A(G2084), .B(G160), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(KEYINPUT113), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(KEYINPUT114), .B(n1012), .ZN(n1022) );
  XOR2_X1 U1100 ( .A(G2090), .B(G162), .Z(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT51), .B(n1015), .Z(n1020) );
  INV_X1 U1103 ( .A(n1016), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1025), .ZN(n1026) );
  NAND2_X1 U1109 ( .A1(G29), .A2(n1026), .ZN(n1027) );
  NAND2_X1 U1110 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1111 ( .A1(n1030), .A2(n1029), .ZN(n1032) );
  XNOR2_X1 U1112 ( .A(KEYINPUT126), .B(KEYINPUT62), .ZN(n1031) );
  XNOR2_X1 U1113 ( .A(n1032), .B(n1031), .ZN(G311) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

