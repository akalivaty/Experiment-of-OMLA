//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n205), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n208), .B(new_n214), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n216), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n239), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G179), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT66), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(KEYINPUT66), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g0059(.A1(new_n251), .A2(new_n256), .A3(G232), .A4(new_n259), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n251), .A2(new_n256), .A3(G238), .A4(G1698), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n249), .A2(new_n250), .A3(new_n248), .ZN(new_n262));
  AOI21_X1  g0062(.A(KEYINPUT66), .B1(new_n254), .B2(new_n255), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G107), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n260), .B(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(G1), .A3(G13), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G1), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(G274), .C1(G41), .C2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(G41), .B2(G45), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n268), .A2(KEYINPUT65), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT65), .B1(new_n268), .B2(new_n274), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n277), .B2(G244), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(KEYINPUT71), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n270), .B2(new_n278), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n247), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n284), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n285));
  AOI21_X1  g0085(.A(KEYINPUT69), .B1(new_n284), .B2(new_n211), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G13), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n288), .A2(new_n212), .A3(G1), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n271), .A2(G20), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(G77), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n288), .A2(G1), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n286), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n284), .A2(KEYINPUT69), .A3(new_n211), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT15), .B(G87), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n212), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(G77), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n298), .A2(new_n299), .B1(new_n212), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT8), .B(G58), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n301), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n292), .B1(G77), .B2(new_n294), .C1(new_n297), .C2(new_n305), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n279), .B(KEYINPUT71), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n283), .B(new_n306), .C1(new_n307), .C2(G169), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n291), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n290), .A2(new_n311), .B1(new_n289), .B2(new_n303), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G58), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n241), .ZN(new_n315));
  OAI21_X1  g0115(.A(G20), .B1(new_n315), .B2(new_n201), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n302), .A2(G159), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n249), .A2(new_n250), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n212), .B1(new_n262), .B2(new_n263), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT7), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n319), .B1(new_n325), .B2(new_n241), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT16), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n254), .A2(new_n255), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n324), .B1(new_n329), .B2(G20), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n321), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n318), .B1(new_n331), .B2(G68), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n297), .B1(new_n332), .B2(KEYINPUT16), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n313), .B1(new_n328), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G223), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G226), .A2(G1698), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n320), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G33), .A2(G87), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n269), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n268), .A2(new_n274), .ZN(new_n343));
  INV_X1    g0143(.A(G232), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n272), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n342), .A2(new_n247), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(KEYINPUT80), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT80), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n259), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n340), .B1(new_n350), .B2(new_n320), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n345), .B1(new_n351), .B2(new_n269), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(new_n247), .ZN(new_n353));
  AOI21_X1  g0153(.A(G169), .B1(new_n342), .B2(new_n346), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n348), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(KEYINPUT18), .B1(new_n334), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(G20), .B1(new_n251), .B2(new_n256), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n321), .B1(new_n358), .B2(KEYINPUT7), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n318), .B1(new_n359), .B2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n333), .B1(KEYINPUT16), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n312), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT18), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n352), .A2(new_n349), .A3(new_n247), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n347), .A2(KEYINPUT80), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n354), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n368), .B1(new_n342), .B2(new_n346), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(G190), .B2(new_n352), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n361), .A2(new_n370), .A3(new_n312), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n334), .A2(KEYINPUT17), .A3(new_n370), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n357), .A2(new_n367), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n280), .A2(new_n282), .ZN(new_n376));
  INV_X1    g0176(.A(G190), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT72), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT72), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(G190), .C1(new_n280), .C2(new_n282), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n306), .B1(new_n376), .B2(G200), .ZN(new_n382));
  AOI211_X1 g0182(.A(new_n309), .B(new_n375), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n310), .A2(new_n241), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n297), .A2(new_n294), .A3(new_n384), .ZN(new_n385));
  XOR2_X1   g0185(.A(new_n385), .B(KEYINPUT76), .Z(new_n386));
  INV_X1    g0186(.A(KEYINPUT12), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n289), .B(new_n241), .C1(KEYINPUT77), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n388), .B(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n241), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n300), .B2(new_n299), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n287), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n287), .A2(new_n392), .ZN(new_n395));
  INV_X1    g0195(.A(new_n393), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n390), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT78), .B1(new_n386), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n398), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT78), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n385), .B(KEYINPUT76), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n251), .A2(new_n256), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n259), .A2(G226), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT73), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(G33), .A2(G97), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n251), .A2(new_n256), .A3(G232), .A4(G1698), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n257), .A2(new_n258), .A3(new_n217), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT73), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(new_n251), .A3(new_n256), .A4(new_n411), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n407), .A2(new_n408), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n269), .ZN(new_n414));
  OAI21_X1  g0214(.A(G238), .B1(new_n275), .B2(new_n276), .ZN(new_n415));
  XNOR2_X1  g0215(.A(new_n272), .B(KEYINPUT74), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n414), .A2(new_n421), .A3(new_n418), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(G190), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n414), .B2(new_n418), .ZN(new_n424));
  AOI211_X1 g0224(.A(KEYINPUT13), .B(new_n417), .C1(new_n413), .C2(new_n269), .ZN(new_n425));
  OAI21_X1  g0225(.A(G200), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n404), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n424), .A2(new_n425), .ZN(new_n428));
  INV_X1    g0228(.A(G169), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT14), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT14), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n431), .B(G169), .C1(new_n424), .C2(new_n425), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT79), .B1(new_n428), .B2(G179), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT79), .ZN(new_n434));
  NOR4_X1   g0234(.A1(new_n424), .A2(new_n425), .A3(new_n434), .A4(new_n247), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n430), .B(new_n432), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n404), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n427), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n264), .A2(G222), .A3(new_n259), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n264), .A2(G223), .A3(G1698), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n300), .C2(new_n264), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n269), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT68), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n273), .B1(new_n277), .B2(G226), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n443), .B1(new_n442), .B2(new_n444), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n247), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n447), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(new_n429), .A3(new_n445), .ZN(new_n450));
  OAI21_X1  g0250(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n451));
  INV_X1    g0251(.A(G150), .ZN(new_n452));
  INV_X1    g0252(.A(new_n302), .ZN(new_n453));
  OAI221_X1 g0253(.A(new_n451), .B1(new_n452), .B2(new_n453), .C1(new_n299), .C2(new_n303), .ZN(new_n454));
  AOI22_X1  g0254(.A1(new_n454), .A2(new_n287), .B1(new_n216), .B2(new_n289), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n291), .A2(G50), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT70), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n290), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n448), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(G190), .B1(new_n446), .B2(new_n447), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n449), .A2(G200), .A3(new_n445), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n459), .B(KEYINPUT9), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT10), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT10), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n462), .A2(new_n463), .A3(new_n467), .A4(new_n464), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n461), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AND3_X1   g0269(.A1(new_n383), .A2(new_n438), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n298), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n294), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n271), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n297), .A2(new_n294), .A3(new_n471), .A4(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(G20), .B1(new_n254), .B2(new_n255), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n476), .A2(G68), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G87), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n480), .A2(new_n481), .A3(new_n265), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT19), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT19), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n408), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n482), .B1(new_n487), .B2(G20), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n473), .B(new_n475), .C1(new_n489), .C2(new_n297), .ZN(new_n490));
  OAI211_X1 g0290(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n329), .A2(KEYINPUT83), .A3(G244), .A4(G1698), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n329), .A2(new_n259), .A3(G238), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G116), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n269), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n271), .A2(G45), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n499), .A2(G250), .ZN(new_n500));
  INV_X1    g0300(.A(G45), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G1), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n500), .A2(new_n268), .B1(G274), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n247), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n503), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n497), .B2(new_n269), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n490), .B(new_n504), .C1(G169), .C2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n498), .A2(G190), .A3(new_n503), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n297), .B1(new_n479), .B2(new_n488), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n294), .B(new_n474), .C1(new_n285), .C2(new_n286), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n480), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n509), .A2(new_n511), .A3(new_n472), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n508), .B(new_n512), .C1(new_n368), .C2(new_n506), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT5), .A2(G41), .ZN(new_n515));
  NOR2_X1   g0315(.A1(KEYINPUT5), .A2(G41), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n502), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(G257), .A3(new_n268), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT81), .ZN(new_n519));
  XNOR2_X1  g0319(.A(KEYINPUT5), .B(G41), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n520), .A2(G274), .A3(new_n268), .A4(new_n502), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n519), .B1(new_n518), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n251), .A2(new_n256), .A3(G250), .A4(G1698), .ZN(new_n525));
  AND2_X1   g0325(.A1(KEYINPUT4), .A2(G244), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n251), .A2(new_n256), .A3(new_n259), .A4(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT4), .ZN(new_n528));
  OAI21_X1  g0328(.A(G244), .B1(new_n249), .B2(new_n250), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n335), .A2(new_n336), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n525), .A2(new_n527), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n269), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n524), .A2(new_n534), .A3(new_n247), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT82), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n510), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n289), .A2(new_n481), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n481), .A3(G107), .ZN(new_n542));
  XNOR2_X1  g0342(.A(G97), .B(G107), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  OAI22_X1  g0344(.A1(new_n544), .A2(new_n212), .B1(new_n300), .B2(new_n453), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n359), .B2(G107), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n539), .B(new_n540), .C1(new_n546), .C2(new_n297), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n524), .A2(new_n534), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n429), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n524), .A2(new_n534), .A3(KEYINPUT82), .A4(new_n247), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n537), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n539), .A2(new_n540), .ZN(new_n552));
  INV_X1    g0352(.A(new_n545), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n325), .B2(new_n265), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n552), .B1(new_n554), .B2(new_n287), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n548), .A2(G200), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n555), .B(new_n556), .C1(new_n377), .C2(new_n548), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n514), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n405), .A2(G303), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n335), .A2(G257), .A3(new_n336), .ZN(new_n560));
  AND2_X1   g0360(.A1(G264), .A2(G1698), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n329), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n268), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n517), .A2(new_n268), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n521), .B1(new_n564), .B2(new_n219), .ZN(new_n565));
  OAI21_X1  g0365(.A(G169), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n284), .A2(new_n211), .B1(G20), .B2(new_n218), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n532), .B(new_n212), .C1(G33), .C2(new_n481), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g0370(.A(new_n570), .B(KEYINPUT20), .Z(new_n571));
  NAND2_X1  g0371(.A1(new_n538), .A2(G116), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n293), .A2(G20), .A3(new_n218), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n567), .A2(KEYINPUT21), .A3(new_n574), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n559), .A2(new_n562), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n565), .B1(new_n577), .B2(new_n269), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n576), .B(new_n579), .C1(new_n368), .C2(new_n578), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT21), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n576), .B2(new_n566), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n563), .A2(new_n247), .A3(new_n565), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n574), .ZN(new_n584));
  AND4_X1   g0384(.A1(new_n575), .A2(new_n580), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT86), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n289), .A2(new_n265), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT25), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n510), .A2(new_n265), .ZN(new_n589));
  OR2_X1    g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n480), .A2(KEYINPUT22), .A3(G20), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n251), .A2(new_n256), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n212), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT22), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n496), .A2(G20), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT23), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n212), .B2(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n265), .A2(KEYINPUT23), .A3(G20), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n595), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n590), .B1(new_n605), .B2(new_n287), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n517), .A2(G264), .A3(new_n268), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n329), .A2(new_n259), .A3(G250), .ZN(new_n609));
  AND2_X1   g0409(.A1(G257), .A2(G1698), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n249), .B2(new_n250), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT85), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n329), .A2(new_n613), .A3(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(G33), .A2(G294), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n609), .A2(new_n612), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n608), .B1(new_n616), .B2(new_n269), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n247), .A3(new_n521), .ZN(new_n618));
  INV_X1    g0418(.A(new_n521), .ZN(new_n619));
  AOI211_X1 g0419(.A(new_n619), .B(new_n608), .C1(new_n616), .C2(new_n269), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(G169), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n586), .B1(new_n606), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n604), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n603), .B1(new_n595), .B2(new_n600), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n287), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n590), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n617), .A2(new_n521), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n429), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n627), .A2(KEYINPUT86), .A3(new_n618), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n616), .A2(new_n269), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(new_n377), .A3(new_n521), .A4(new_n607), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT87), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n632), .B(KEYINPUT87), .C1(new_n620), .C2(G200), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(new_n606), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n622), .A2(new_n630), .A3(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n470), .A2(new_n558), .A3(new_n585), .A4(new_n636), .ZN(G372));
  NAND2_X1  g0437(.A1(new_n357), .A2(new_n367), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n436), .A2(new_n437), .ZN(new_n640));
  INV_X1    g0440(.A(new_n427), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n309), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n373), .A2(new_n374), .ZN(new_n644));
  OAI211_X1 g0444(.A(KEYINPUT91), .B(new_n639), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n466), .A2(new_n468), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT91), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n644), .B1(new_n640), .B2(new_n642), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n647), .B1(new_n648), .B2(new_n638), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n460), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n383), .A2(new_n438), .A3(new_n469), .ZN(new_n653));
  INV_X1    g0453(.A(new_n621), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(new_n627), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT88), .B1(new_n606), .B2(new_n621), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n582), .A2(new_n575), .A3(new_n584), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n551), .A2(new_n514), .A3(new_n635), .A4(new_n557), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT89), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n659), .B1(new_n656), .B2(new_n657), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n514), .A2(new_n635), .A3(new_n557), .A4(new_n551), .ZN(new_n666));
  OAI21_X1  g0466(.A(KEYINPUT89), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n537), .A2(new_n549), .A3(new_n547), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n669), .A2(new_n514), .A3(KEYINPUT26), .A4(new_n550), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n507), .A2(new_n513), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n671), .B1(new_n551), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n668), .B1(new_n674), .B2(new_n507), .ZN(new_n675));
  INV_X1    g0475(.A(new_n507), .ZN(new_n676));
  AOI211_X1 g0476(.A(KEYINPUT90), .B(new_n676), .C1(new_n670), .C2(new_n673), .ZN(new_n677));
  OAI211_X1 g0477(.A(new_n664), .B(new_n667), .C1(new_n675), .C2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n652), .B1(new_n653), .B2(new_n679), .ZN(G369));
  INV_X1    g0480(.A(KEYINPUT27), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n293), .A2(new_n681), .A3(new_n212), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT92), .ZN(new_n683));
  INV_X1    g0483(.A(G213), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n293), .A2(new_n212), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(KEYINPUT27), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G343), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT93), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT94), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n690), .A2(new_n691), .A3(new_n576), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT94), .B1(new_n689), .B2(new_n574), .ZN(new_n693));
  OR3_X1    g0493(.A1(new_n692), .A2(new_n585), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n660), .B1(new_n692), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n696), .B(KEYINPUT95), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n636), .B1(new_n606), .B2(new_n690), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n689), .A2(new_n654), .A3(new_n627), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n656), .A2(new_n657), .A3(new_n690), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n660), .A2(new_n689), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n636), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n206), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n482), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n209), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n622), .A2(new_n630), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n558), .B(new_n635), .C1(new_n659), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n676), .B1(new_n670), .B2(new_n673), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n689), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n675), .A2(new_n677), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n664), .A2(new_n667), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n690), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n578), .A2(new_n506), .A3(new_n617), .A4(G179), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT96), .B(new_n725), .C1(new_n726), .C2(new_n548), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n578), .A2(new_n506), .A3(G179), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n548), .A3(new_n628), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n725), .B1(new_n726), .B2(new_n548), .ZN(new_n731));
  INV_X1    g0531(.A(new_n548), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n506), .A2(new_n617), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT30), .A4(new_n583), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(KEYINPUT96), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n730), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n724), .B1(new_n736), .B2(new_n690), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n636), .A2(new_n558), .A3(new_n585), .A4(new_n690), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n729), .A3(new_n731), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n723), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n713), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n288), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n271), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OR3_X1    g0548(.A1(new_n708), .A2(new_n748), .A3(KEYINPUT97), .ZN(new_n749));
  OAI21_X1  g0549(.A(KEYINPUT97), .B1(new_n708), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n698), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G330), .B2(new_n697), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT98), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n211), .B1(G20), .B2(new_n429), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n212), .A2(new_n377), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n368), .A2(G179), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G303), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n247), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G322), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n212), .A2(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n765), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n247), .A2(new_n368), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n760), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n764), .B(new_n771), .C1(G326), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n761), .A2(new_n768), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G283), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n772), .A2(new_n768), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n768), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n780), .A2(new_n781), .B1(new_n784), .B2(G329), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n212), .B1(new_n782), .B2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n264), .B1(G294), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n775), .A2(new_n778), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n776), .A2(new_n265), .ZN(new_n790));
  INV_X1    g0590(.A(new_n766), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n405), .B(new_n790), .C1(G58), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(G97), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n773), .A2(new_n216), .B1(new_n762), .B2(new_n480), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n779), .A2(new_n241), .B1(new_n769), .B2(new_n300), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n792), .A2(new_n793), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n759), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n758), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT99), .Z(new_n806));
  NOR2_X1   g0606(.A1(new_n707), .A2(new_n329), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n501), .B2(new_n210), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n245), .B2(new_n501), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n405), .A2(new_n707), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n811), .A2(G355), .B1(new_n218), .B2(new_n707), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n806), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n801), .A2(new_n751), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n804), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n697), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n756), .A2(new_n757), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n308), .A2(new_n689), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n381), .A2(new_n382), .B1(new_n306), .B2(new_n689), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n821), .B2(new_n309), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n721), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n379), .B1(new_n307), .B2(G190), .ZN(new_n824));
  INV_X1    g0624(.A(new_n380), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n382), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n689), .A2(new_n306), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n819), .B1(new_n828), .B2(new_n308), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n678), .A2(new_n690), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n823), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n752), .B1(new_n831), .B2(new_n742), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n742), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n779), .A2(new_n452), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT101), .B(G143), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n766), .A2(new_n835), .B1(new_n769), .B2(new_n794), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(G137), .C2(new_n774), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  INV_X1    g0638(.A(G132), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n329), .B1(new_n783), .B2(new_n839), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n762), .A2(new_n216), .B1(new_n776), .B2(new_n241), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(G58), .C2(new_n787), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(KEYINPUT34), .B2(new_n837), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n773), .A2(new_n763), .B1(new_n762), .B2(new_n265), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(G294), .B2(new_n791), .ZN(new_n846));
  INV_X1    g0646(.A(G283), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n779), .A2(new_n847), .B1(new_n776), .B2(new_n480), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n769), .A2(new_n218), .B1(new_n783), .B2(new_n770), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n846), .A2(new_n405), .A3(new_n793), .A4(new_n850), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n851), .B(KEYINPUT100), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n758), .B1(new_n844), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n758), .A2(new_n802), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n751), .B1(new_n300), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n853), .B(new_n855), .C1(new_n829), .C2(new_n803), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n833), .A2(new_n856), .ZN(G384));
  INV_X1    g0657(.A(new_n544), .ZN(new_n858));
  OR2_X1    g0658(.A1(new_n858), .A2(KEYINPUT35), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(KEYINPUT35), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n859), .A2(G116), .A3(new_n213), .A4(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT36), .Z(new_n862));
  OR3_X1    g0662(.A1(new_n209), .A2(new_n300), .A3(new_n315), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n271), .B(G13), .C1(new_n863), .C2(new_n240), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n717), .A2(KEYINPUT29), .ZN(new_n866));
  AND4_X1   g0666(.A1(new_n550), .A2(new_n537), .A3(new_n549), .A4(new_n547), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT26), .B1(new_n867), .B2(new_n514), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n551), .A2(new_n672), .A3(new_n671), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n507), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT90), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n716), .A2(new_n668), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n664), .A2(new_n667), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n689), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n470), .B(new_n866), .C1(new_n875), .C2(KEYINPUT29), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT102), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n721), .A2(new_n722), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n878), .A2(new_n879), .A3(new_n470), .A4(new_n866), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n651), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n690), .A2(new_n404), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n427), .B(new_n882), .C1(new_n436), .C2(new_n437), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n436), .A2(new_n437), .A3(new_n689), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n830), .B2(new_n820), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n331), .A2(G68), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(KEYINPUT16), .A3(new_n319), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n241), .B1(new_n330), .B2(new_n321), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n327), .B1(new_n890), .B2(new_n318), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n891), .A3(new_n287), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n312), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n687), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n375), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n366), .A2(new_n893), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n371), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(KEYINPUT37), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n362), .A2(new_n366), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n362), .A2(new_n687), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n371), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n896), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n887), .A2(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n896), .A2(KEYINPUT38), .A3(new_n904), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n371), .B1(new_n334), .B2(new_n356), .ZN(new_n913));
  INV_X1    g0713(.A(new_n687), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n334), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT37), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n903), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n375), .A2(new_n915), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n920), .A2(KEYINPUT39), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n640), .A2(new_n689), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n638), .A2(new_n914), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n911), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(new_n881), .B(new_n926), .Z(new_n927));
  INV_X1    g0727(.A(G330), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n735), .A2(new_n731), .ZN(new_n929));
  OAI211_X1 g0729(.A(KEYINPUT31), .B(new_n689), .C1(new_n929), .C2(new_n730), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n737), .A2(new_n930), .A3(new_n738), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n829), .B(new_n931), .C1(new_n883), .C2(new_n885), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT40), .B1(new_n932), .B2(new_n920), .ZN(new_n933));
  INV_X1    g0733(.A(new_n882), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n640), .A2(new_n641), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n822), .B1(new_n935), .B2(new_n884), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT40), .B1(new_n907), .B2(new_n908), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n936), .A2(new_n937), .A3(new_n931), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n470), .A2(new_n931), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n928), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n940), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n927), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n271), .B2(new_n746), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n927), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n865), .B1(new_n944), .B2(new_n945), .ZN(G367));
  INV_X1    g0746(.A(new_n806), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n206), .B2(new_n298), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n235), .A2(new_n808), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n752), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n773), .A2(new_n835), .B1(new_n779), .B2(new_n794), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(G137), .B2(new_n784), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n314), .A2(new_n762), .B1(new_n766), .B2(new_n452), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n216), .A2(new_n769), .B1(new_n776), .B2(new_n300), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n787), .A2(G68), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n952), .A2(new_n264), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n762), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(G116), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT46), .ZN(new_n960));
  AOI22_X1  g0760(.A1(G294), .A2(new_n780), .B1(new_n791), .B2(G303), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n960), .B(new_n961), .C1(new_n847), .C2(new_n769), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n774), .A2(G311), .B1(new_n777), .B2(G97), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n329), .B1(new_n784), .B2(G317), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n265), .C2(new_n786), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n957), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n950), .B1(new_n967), .B2(new_n758), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n690), .A2(new_n512), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(new_n514), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n968), .B1(new_n971), .B2(new_n815), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n705), .A2(new_n703), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n551), .B(new_n557), .C1(new_n690), .C2(new_n555), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n867), .A2(new_n689), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n973), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT44), .Z(new_n979));
  NOR2_X1   g0779(.A1(new_n973), .A2(new_n977), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(new_n698), .A3(new_n701), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n705), .B1(new_n701), .B2(new_n704), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n698), .B(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n702), .A2(new_n981), .A3(new_n979), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n983), .A2(new_n985), .A3(new_n744), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n744), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n708), .B(KEYINPUT41), .Z(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n748), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n977), .A2(new_n705), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT42), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n714), .A2(new_n557), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n689), .B1(new_n995), .B2(new_n551), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n993), .B2(KEYINPUT42), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n994), .A2(new_n997), .B1(KEYINPUT43), .B2(new_n971), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n702), .A2(new_n977), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1000), .B(new_n1001), .Z(new_n1002));
  OAI21_X1  g0802(.A(new_n972), .B1(new_n991), .B2(new_n1002), .ZN(G387));
  OR2_X1    g0803(.A1(new_n698), .A2(new_n984), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n698), .A2(new_n984), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n747), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT103), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(KEYINPUT103), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n699), .A2(new_n700), .A3(new_n804), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n304), .A2(new_n216), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT50), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n710), .B(new_n501), .C1(new_n241), .C2(new_n300), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n807), .B1(new_n1011), .B2(new_n1012), .C1(new_n232), .C2(new_n501), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n710), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n811), .A2(new_n1014), .B1(new_n265), .B2(new_n707), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(KEYINPUT104), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n947), .ZN(new_n1017));
  AOI21_X1  g0817(.A(KEYINPUT104), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n752), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n786), .A2(new_n298), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n320), .B(new_n1020), .C1(G97), .C2(new_n777), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n774), .A2(KEYINPUT106), .A3(G159), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT106), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n773), .B2(new_n794), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n762), .A2(new_n300), .B1(new_n783), .B2(new_n452), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n1022), .A2(new_n1024), .B1(new_n1025), .B2(KEYINPUT105), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n779), .A2(new_n303), .B1(new_n769), .B2(new_n241), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G50), .B2(new_n791), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1025), .A2(KEYINPUT105), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1021), .A2(new_n1026), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n329), .B1(new_n784), .B2(G326), .ZN(new_n1031));
  INV_X1    g0831(.A(G294), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n762), .A2(new_n1032), .B1(new_n786), .B2(new_n847), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT107), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n769), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G317), .A2(new_n791), .B1(new_n1035), .B2(G303), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n770), .B2(new_n779), .C1(new_n767), .C2(new_n773), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT108), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1034), .B1(new_n1038), .B2(KEYINPUT48), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(KEYINPUT48), .B2(new_n1038), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT49), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1031), .B1(new_n218), .B2(new_n776), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1030), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1019), .B1(new_n1044), .B2(new_n758), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1007), .A2(new_n1008), .B1(new_n1009), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n985), .A2(new_n744), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n985), .A2(new_n744), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n708), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1046), .B1(new_n1047), .B2(new_n1049), .ZN(G393));
  INV_X1    g0850(.A(KEYINPUT109), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n986), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n986), .A2(new_n1051), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n983), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n747), .B1(new_n1054), .B2(KEYINPUT110), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(KEYINPUT110), .B2(new_n1054), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1048), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1057), .A2(new_n708), .A3(new_n987), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n947), .B1(new_n481), .B2(new_n206), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n239), .A2(new_n808), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n752), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT111), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n762), .A2(new_n241), .B1(new_n783), .B2(new_n835), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n320), .B(new_n1063), .C1(G87), .C2(new_n777), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT112), .Z(new_n1065));
  OAI22_X1  g0865(.A1(new_n773), .A2(new_n452), .B1(new_n766), .B2(new_n794), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT51), .Z(new_n1067));
  NAND2_X1  g0867(.A1(new_n787), .A2(G77), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n216), .B2(new_n779), .C1(new_n303), .C2(new_n769), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1070), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1071), .A2(KEYINPUT113), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(KEYINPUT113), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G317), .A2(new_n774), .B1(new_n791), .B2(G311), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  AOI211_X1 g0875(.A(new_n790), .B(new_n264), .C1(G303), .C2(new_n780), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n769), .A2(new_n1032), .B1(new_n783), .B2(new_n767), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G283), .B2(new_n958), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n787), .A2(G116), .ZN(new_n1079));
  AND4_X1   g0879(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1072), .A2(new_n1073), .A3(new_n1080), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1062), .B1(new_n815), .B2(new_n976), .C1(new_n1081), .C2(new_n759), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1056), .A2(new_n1058), .A3(new_n1082), .ZN(G390));
  NAND2_X1  g0883(.A1(new_n921), .A2(new_n923), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n887), .B2(new_n922), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n936), .A2(new_n743), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n828), .A2(new_n308), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n717), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n820), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n935), .A2(new_n884), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n922), .B(new_n920), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n1085), .A2(new_n1086), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n931), .A2(G330), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n936), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n470), .A2(new_n1095), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n879), .B1(new_n723), .B2(new_n470), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT29), .B1(new_n678), .B2(new_n690), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1101), .A2(KEYINPUT102), .A3(new_n718), .A4(new_n653), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n652), .B(new_n1099), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n886), .B1(new_n742), .B2(new_n822), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n830), .A2(new_n820), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n886), .B1(new_n1094), .B2(new_n822), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1086), .A2(new_n1108), .A3(new_n820), .A4(new_n1088), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT114), .B1(new_n1098), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n709), .B1(new_n1098), .B2(new_n1111), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1085), .A2(new_n1092), .A3(new_n1086), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n922), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n819), .B1(new_n875), .B2(new_n829), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n886), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1091), .B1(new_n1117), .B2(new_n1084), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1114), .B1(new_n1118), .B2(new_n1096), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n881), .A2(new_n1099), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1112), .A2(new_n1113), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n854), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n958), .A2(G150), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT53), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n769), .A2(new_n1128), .B1(new_n783), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(G128), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n773), .A2(new_n1131), .B1(new_n766), .B2(new_n839), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1127), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(G137), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n779), .A2(new_n1134), .B1(new_n776), .B2(new_n216), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n405), .B(new_n1135), .C1(G159), .C2(new_n787), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n405), .B1(new_n480), .B2(new_n762), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT116), .Z(new_n1138));
  OAI221_X1 g0938(.A(new_n1068), .B1(new_n241), .B2(new_n776), .C1(new_n1032), .C2(new_n783), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n779), .A2(new_n265), .B1(new_n769), .B2(new_n481), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n773), .A2(new_n847), .B1(new_n766), .B2(new_n218), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1133), .A2(new_n1136), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n752), .B1(new_n304), .B2(new_n1125), .C1(new_n1143), .C2(new_n759), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n1084), .B2(new_n802), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1098), .A2(KEYINPUT115), .A3(new_n748), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT115), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n1119), .B2(new_n747), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1145), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1124), .A2(new_n1149), .ZN(G378));
  INV_X1    g0950(.A(new_n1103), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1119), .B2(new_n1110), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT117), .B1(new_n939), .B2(G330), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT117), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1154), .B(new_n928), .C1(new_n933), .C2(new_n938), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n459), .A2(new_n687), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n469), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n469), .A2(new_n1157), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1156), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1156), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1162), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1153), .A2(new_n1155), .A3(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(KEYINPUT117), .B(new_n1165), .C1(G330), .C2(new_n939), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n926), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n932), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n903), .A2(new_n916), .B1(new_n375), .B2(new_n915), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n908), .B1(new_n1171), .B2(KEYINPUT38), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1090), .A2(new_n1172), .A3(new_n829), .A4(new_n931), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1170), .A2(new_n937), .B1(new_n1173), .B2(KEYINPUT40), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1154), .B1(new_n1174), .B2(new_n928), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n939), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n1176), .A3(new_n1165), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n926), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1154), .B(new_n1166), .C1(new_n1174), .C2(new_n928), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1152), .A2(new_n1169), .A3(KEYINPUT57), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT118), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1178), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT118), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(KEYINPUT57), .A4(new_n1152), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT57), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1169), .A2(new_n1180), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1103), .B1(new_n1098), .B2(new_n1111), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1182), .A2(new_n1187), .A3(new_n1191), .A4(new_n708), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1165), .A2(new_n802), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n752), .B1(G50), .B2(new_n1125), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n773), .A2(new_n1129), .B1(new_n779), .B2(new_n839), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1035), .A2(G137), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1196), .B1(new_n1131), .B2(new_n766), .C1(new_n762), .C2(new_n1128), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G150), .C2(new_n787), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT59), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n777), .A2(G159), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G33), .B(G41), .C1(new_n784), .C2(G124), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n776), .A2(new_n314), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G283), .B2(new_n784), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G41), .B(new_n329), .C1(new_n958), .C2(G77), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n956), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n773), .A2(new_n218), .B1(new_n769), .B2(new_n298), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n481), .A2(new_n779), .B1(new_n766), .B2(new_n265), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(KEYINPUT58), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(KEYINPUT58), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n216), .B1(new_n249), .B2(G41), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1204), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1194), .B1(new_n1215), .B2(new_n758), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1185), .A2(new_n748), .B1(new_n1193), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1192), .A2(new_n1217), .ZN(G375));
  AND3_X1   g1018(.A1(new_n1103), .A2(KEYINPUT119), .A3(new_n1110), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT119), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1221), .A2(new_n990), .A3(new_n1122), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1110), .A2(new_n747), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n886), .A2(new_n802), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT120), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n774), .A2(G132), .B1(new_n784), .B2(G128), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n1134), .B2(new_n766), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n794), .A2(new_n762), .B1(new_n779), .B2(new_n1128), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1227), .A2(new_n320), .A3(new_n1205), .A4(new_n1228), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n769), .A2(new_n452), .B1(new_n786), .B2(new_n216), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT121), .ZN(new_n1231));
  OAI22_X1  g1031(.A1(new_n766), .A2(new_n847), .B1(new_n783), .B2(new_n763), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G107), .B2(new_n1035), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n773), .A2(new_n1032), .B1(new_n776), .B2(new_n300), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n481), .A2(new_n762), .B1(new_n779), .B2(new_n218), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n264), .A4(new_n1020), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n1229), .A2(new_n1231), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n752), .B1(G68), .B2(new_n1125), .C1(new_n1237), .C2(new_n759), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1225), .A2(new_n1238), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1223), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1222), .A2(new_n1241), .ZN(G381));
  NOR3_X1   g1042(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT122), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1243), .B(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G378), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1192), .A2(new_n1246), .A3(new_n1217), .ZN(new_n1247));
  OR2_X1    g1047(.A1(G390), .A2(G387), .ZN(new_n1248));
  OR4_X1    g1048(.A1(G381), .A2(new_n1245), .A3(new_n1247), .A4(new_n1248), .ZN(G407));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(G343), .C2(new_n1247), .ZN(G409));
  XNOR2_X1  g1050(.A(G393), .B(G396), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G390), .A2(G387), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(G390), .A2(G387), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1248), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G375), .A2(G378), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1103), .A2(new_n1110), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT119), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1103), .A2(KEYINPUT119), .A3(new_n1110), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1122), .A2(KEYINPUT60), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1121), .B1(new_n881), .B2(new_n1099), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n709), .B1(new_n1266), .B2(KEYINPUT60), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G384), .B1(new_n1268), .B2(new_n1241), .ZN(new_n1269));
  INV_X1    g1069(.A(G384), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1270), .B(new_n1240), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(G343), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(G213), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1152), .A2(new_n1169), .A3(new_n990), .A4(new_n1180), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1193), .A2(new_n1216), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1275), .B(new_n1276), .C1(new_n747), .C2(new_n1189), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1274), .B1(new_n1277), .B2(G378), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1259), .A2(new_n1272), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(KEYINPUT62), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(G375), .B2(G378), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1273), .A2(G213), .A3(G2897), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n708), .B1(new_n1260), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1221), .B2(new_n1264), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1270), .B1(new_n1288), .B2(new_n1240), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1268), .A2(G384), .A3(new_n1241), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1284), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1285), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(KEYINPUT126), .B(new_n1282), .C1(new_n1283), .C2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT62), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1283), .A2(new_n1295), .A3(new_n1272), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1281), .A2(new_n1294), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1285), .A2(new_n1292), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1246), .B1(new_n1192), .B2(new_n1217), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1298), .B1(new_n1299), .B2(new_n1278), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT126), .B1(new_n1300), .B2(new_n1282), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1258), .B1(new_n1297), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1298), .B(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT124), .B1(new_n1299), .B2(new_n1278), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT124), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1283), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1280), .A2(KEYINPUT123), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(KEYINPUT63), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT63), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1280), .A2(KEYINPUT123), .A3(new_n1311), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1256), .A2(new_n1257), .A3(new_n1282), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1308), .A2(new_n1310), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1302), .A2(new_n1314), .ZN(G405));
  NAND3_X1  g1115(.A1(new_n1256), .A2(new_n1257), .A3(KEYINPUT127), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1259), .A2(new_n1247), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1259), .A2(new_n1247), .A3(new_n1272), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1316), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT127), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1320), .A2(new_n1321), .A3(new_n1258), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1258), .A2(new_n1321), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1323), .A2(new_n1318), .A3(new_n1319), .A4(new_n1316), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(G402));
endmodule


