

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n361) );
  XOR2_X1 U324 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n291) );
  XOR2_X1 U325 ( .A(n335), .B(n334), .Z(n292) );
  NOR2_X1 U326 ( .A1(n529), .A2(n366), .ZN(n367) );
  XNOR2_X1 U327 ( .A(n362), .B(n361), .ZN(n369) );
  XNOR2_X1 U328 ( .A(n296), .B(KEYINPUT73), .ZN(n297) );
  NAND2_X1 U329 ( .A1(n369), .A2(n368), .ZN(n370) );
  XNOR2_X1 U330 ( .A(n298), .B(n297), .ZN(n302) );
  XNOR2_X1 U331 ( .A(n370), .B(KEYINPUT48), .ZN(n541) );
  XOR2_X1 U332 ( .A(n340), .B(n339), .Z(n560) );
  XNOR2_X1 U333 ( .A(n451), .B(KEYINPUT120), .ZN(n452) );
  XNOR2_X1 U334 ( .A(n453), .B(n452), .ZN(G1350GAT) );
  XNOR2_X1 U335 ( .A(G120GAT), .B(G148GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n293), .B(G57GAT), .ZN(n393) );
  XOR2_X1 U337 ( .A(G99GAT), .B(G85GAT), .Z(n335) );
  XNOR2_X1 U338 ( .A(n393), .B(n335), .ZN(n295) );
  AND2_X1 U339 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n298) );
  XOR2_X1 U341 ( .A(G71GAT), .B(KEYINPUT13), .Z(n350) );
  XOR2_X1 U342 ( .A(n350), .B(KEYINPUT72), .Z(n296) );
  XOR2_X1 U343 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n300) );
  XNOR2_X1 U344 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U346 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U347 ( .A(G78GAT), .B(G204GAT), .Z(n304) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n419) );
  XNOR2_X1 U350 ( .A(G176GAT), .B(G92GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n305), .B(G64GAT), .ZN(n384) );
  XNOR2_X1 U352 ( .A(n419), .B(n384), .ZN(n306) );
  XNOR2_X1 U353 ( .A(n307), .B(n306), .ZN(n573) );
  XOR2_X1 U354 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n308) );
  XOR2_X1 U355 ( .A(n573), .B(n308), .Z(n501) );
  XOR2_X1 U356 ( .A(KEYINPUT8), .B(G50GAT), .Z(n310) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G36GAT), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U359 ( .A(KEYINPUT7), .B(n311), .Z(n340) );
  XOR2_X1 U360 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n313) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n340), .B(n314), .ZN(n324) );
  XOR2_X1 U364 ( .A(G169GAT), .B(G8GAT), .Z(n380) );
  XNOR2_X1 U365 ( .A(G22GAT), .B(G15GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n315), .B(KEYINPUT67), .ZN(n354) );
  XOR2_X1 U367 ( .A(n380), .B(n354), .Z(n317) );
  NAND2_X1 U368 ( .A1(G229GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n320) );
  XOR2_X1 U370 ( .A(G1GAT), .B(G113GAT), .Z(n319) );
  XNOR2_X1 U371 ( .A(G29GAT), .B(G141GAT), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n397) );
  XOR2_X1 U373 ( .A(n320), .B(n397), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT66), .B(KEYINPUT68), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U376 ( .A(n324), .B(n323), .Z(n544) );
  OR2_X1 U377 ( .A1(n501), .A2(n544), .ZN(n326) );
  XOR2_X1 U378 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n360) );
  XOR2_X1 U380 ( .A(G92GAT), .B(G162GAT), .Z(n328) );
  XNOR2_X1 U381 ( .A(G29GAT), .B(G106GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U383 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n330) );
  XNOR2_X1 U384 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n338) );
  XNOR2_X1 U387 ( .A(G190GAT), .B(G218GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n291), .B(n333), .ZN(n334) );
  NAND2_X1 U389 ( .A1(G232GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n292), .B(n336), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U392 ( .A(KEYINPUT76), .B(G64GAT), .Z(n342) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G127GAT), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U395 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n344) );
  XNOR2_X1 U396 ( .A(G1GAT), .B(G57GAT), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n358) );
  XOR2_X1 U399 ( .A(G155GAT), .B(G78GAT), .Z(n348) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G211GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U402 ( .A(n350), .B(n349), .Z(n352) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U405 ( .A(n353), .B(KEYINPUT12), .Z(n356) );
  XNOR2_X1 U406 ( .A(n354), .B(KEYINPUT77), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U408 ( .A(n358), .B(n357), .Z(n576) );
  INV_X1 U409 ( .A(n576), .ZN(n470) );
  NAND2_X1 U410 ( .A1(n560), .A2(n470), .ZN(n359) );
  OR2_X1 U411 ( .A1(n360), .A2(n359), .ZN(n362) );
  XOR2_X1 U412 ( .A(n544), .B(KEYINPUT69), .Z(n555) );
  INV_X1 U413 ( .A(n555), .ZN(n529) );
  INV_X1 U414 ( .A(n560), .ZN(n552) );
  XOR2_X1 U415 ( .A(n552), .B(KEYINPUT101), .Z(n363) );
  XNOR2_X1 U416 ( .A(n363), .B(KEYINPUT36), .ZN(n579) );
  NAND2_X1 U417 ( .A1(n579), .A2(n576), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n364), .B(KEYINPUT114), .ZN(n365) );
  XNOR2_X1 U419 ( .A(n365), .B(KEYINPUT45), .ZN(n366) );
  INV_X1 U420 ( .A(n573), .ZN(n456) );
  NAND2_X1 U421 ( .A1(n367), .A2(n456), .ZN(n368) );
  XOR2_X1 U422 ( .A(KEYINPUT18), .B(G190GAT), .Z(n372) );
  XNOR2_X1 U423 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U425 ( .A(KEYINPUT17), .B(n373), .Z(n446) );
  XOR2_X1 U426 ( .A(KEYINPUT82), .B(G218GAT), .Z(n375) );
  XNOR2_X1 U427 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U429 ( .A(G197GAT), .B(n376), .Z(n429) );
  XNOR2_X1 U430 ( .A(n446), .B(n429), .ZN(n388) );
  XOR2_X1 U431 ( .A(KEYINPUT76), .B(KEYINPUT92), .Z(n378) );
  XNOR2_X1 U432 ( .A(G36GAT), .B(G204GAT), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U434 ( .A(n380), .B(n379), .Z(n382) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U437 ( .A(n383), .B(KEYINPUT93), .Z(n386) );
  XNOR2_X1 U438 ( .A(n384), .B(KEYINPUT91), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n518) );
  NAND2_X1 U441 ( .A1(n541), .A2(n518), .ZN(n390) );
  XOR2_X1 U442 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n413) );
  XOR2_X1 U444 ( .A(KEYINPUT86), .B(KEYINPUT89), .Z(n392) );
  XNOR2_X1 U445 ( .A(G85GAT), .B(KEYINPUT6), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U447 ( .A(n394), .B(n393), .Z(n399) );
  XOR2_X1 U448 ( .A(G155GAT), .B(KEYINPUT2), .Z(n396) );
  XNOR2_X1 U449 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n395) );
  XNOR2_X1 U450 ( .A(n396), .B(n395), .ZN(n418) );
  XNOR2_X1 U451 ( .A(n397), .B(n418), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n412) );
  XOR2_X1 U453 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n401) );
  XNOR2_X1 U454 ( .A(KEYINPUT84), .B(KEYINPUT5), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(KEYINPUT87), .B(n402), .Z(n404) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U459 ( .A(n405), .B(KEYINPUT1), .Z(n410) );
  XOR2_X1 U460 ( .A(KEYINPUT79), .B(G134GAT), .Z(n407) );
  XNOR2_X1 U461 ( .A(KEYINPUT78), .B(G127GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(KEYINPUT0), .B(n408), .ZN(n432) );
  XOR2_X1 U464 ( .A(n432), .B(KEYINPUT85), .Z(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U466 ( .A(n412), .B(n411), .Z(n463) );
  XNOR2_X1 U467 ( .A(KEYINPUT90), .B(n463), .ZN(n516) );
  NOR2_X2 U468 ( .A1(n413), .A2(n516), .ZN(n565) );
  XOR2_X1 U469 ( .A(KEYINPUT23), .B(KEYINPUT81), .Z(n415) );
  XNOR2_X1 U470 ( .A(G22GAT), .B(KEYINPUT83), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U472 ( .A(G50GAT), .B(KEYINPUT74), .Z(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n425) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U475 ( .A(G148GAT), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(KEYINPUT22), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n427) );
  NAND2_X1 U480 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n464) );
  NAND2_X1 U483 ( .A1(n565), .A2(n464), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n430), .B(KEYINPUT55), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n431), .B(KEYINPUT118), .ZN(n447) );
  INV_X1 U486 ( .A(n432), .ZN(n440) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XOR2_X1 U488 ( .A(G71GAT), .B(G120GAT), .Z(n434) );
  XNOR2_X1 U489 ( .A(G113GAT), .B(G15GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U491 ( .A(G43GAT), .B(G99GAT), .Z(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n440), .B(n439), .Z(n444) );
  XOR2_X1 U495 ( .A(G176GAT), .B(KEYINPUT20), .Z(n442) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(KEYINPUT80), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n526) );
  NAND2_X1 U500 ( .A1(n447), .A2(n526), .ZN(n554) );
  NOR2_X1 U501 ( .A1(n501), .A2(n554), .ZN(n450) );
  XNOR2_X1 U502 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n448), .B(G176GAT), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(G1349GAT) );
  NOR2_X1 U505 ( .A1(n470), .A2(n554), .ZN(n453) );
  INV_X1 U506 ( .A(G183GAT), .ZN(n451) );
  XNOR2_X1 U507 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n454), .B(KEYINPUT97), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT96), .B(n455), .Z(n475) );
  NAND2_X1 U510 ( .A1(n529), .A2(n456), .ZN(n488) );
  NAND2_X1 U511 ( .A1(n518), .A2(n526), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n464), .A2(n457), .ZN(n458) );
  XNOR2_X1 U513 ( .A(n458), .B(KEYINPUT25), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n518), .B(KEYINPUT27), .ZN(n465) );
  NOR2_X1 U515 ( .A1(n526), .A2(n464), .ZN(n459) );
  XNOR2_X1 U516 ( .A(KEYINPUT26), .B(n459), .ZN(n566) );
  AND2_X1 U517 ( .A1(n465), .A2(n566), .ZN(n460) );
  NOR2_X1 U518 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n463), .A2(n462), .ZN(n469) );
  XOR2_X1 U520 ( .A(KEYINPUT28), .B(n464), .Z(n523) );
  INV_X1 U521 ( .A(n523), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n465), .A2(n516), .ZN(n466) );
  XOR2_X1 U523 ( .A(KEYINPUT94), .B(n466), .Z(n540) );
  NAND2_X1 U524 ( .A1(n467), .A2(n540), .ZN(n528) );
  NOR2_X1 U525 ( .A1(n528), .A2(n526), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n484) );
  NOR2_X1 U527 ( .A1(n470), .A2(n552), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  NOR2_X1 U529 ( .A1(n484), .A2(n472), .ZN(n473) );
  XNOR2_X1 U530 ( .A(KEYINPUT95), .B(n473), .ZN(n502) );
  NOR2_X1 U531 ( .A1(n488), .A2(n502), .ZN(n482) );
  NAND2_X1 U532 ( .A1(n482), .A2(n516), .ZN(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n482), .A2(n518), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT98), .ZN(n477) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n479) );
  NAND2_X1 U538 ( .A1(n482), .A2(n526), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n481) );
  XOR2_X1 U540 ( .A(G15GAT), .B(KEYINPUT99), .Z(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U542 ( .A1(n523), .A2(n482), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n491) );
  NOR2_X1 U545 ( .A1(n484), .A2(n576), .ZN(n485) );
  XNOR2_X1 U546 ( .A(KEYINPUT102), .B(n485), .ZN(n486) );
  NAND2_X1 U547 ( .A1(n486), .A2(n579), .ZN(n487) );
  XOR2_X1 U548 ( .A(KEYINPUT37), .B(n487), .Z(n515) );
  NOR2_X1 U549 ( .A1(n515), .A2(n488), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT38), .B(n489), .ZN(n497) );
  NAND2_X1 U551 ( .A1(n497), .A2(n516), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NAND2_X1 U554 ( .A1(n497), .A2(n518), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n495) );
  NAND2_X1 U557 ( .A1(n497), .A2(n526), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n496), .Z(G1330GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n499) );
  NAND2_X1 U561 ( .A1(n497), .A2(n523), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n505) );
  INV_X1 U565 ( .A(n501), .ZN(n546) );
  NAND2_X1 U566 ( .A1(n546), .A2(n544), .ZN(n514) );
  NOR2_X1 U567 ( .A1(n514), .A2(n502), .ZN(n503) );
  XOR2_X1 U568 ( .A(KEYINPUT107), .B(n503), .Z(n510) );
  NAND2_X1 U569 ( .A1(n510), .A2(n516), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n506), .Z(G1332GAT) );
  NAND2_X1 U572 ( .A1(n510), .A2(n518), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U574 ( .A(G71GAT), .B(KEYINPUT109), .Z(n509) );
  NAND2_X1 U575 ( .A1(n510), .A2(n526), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n509), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n512) );
  NAND2_X1 U578 ( .A1(n510), .A2(n523), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n522) );
  NAND2_X1 U582 ( .A1(n522), .A2(n516), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT111), .Z(n521) );
  NAND2_X1 U587 ( .A1(n522), .A2(n526), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT115), .Z(n531) );
  NAND2_X1 U593 ( .A1(n541), .A2(n526), .ZN(n527) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n537), .A2(n529), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U598 ( .A1(n537), .A2(n546), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U601 ( .A1(n537), .A2(n576), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U605 ( .A1(n537), .A2(n552), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  INV_X1 U607 ( .A(n566), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n551) );
  INV_X1 U610 ( .A(n544), .ZN(n568) );
  NAND2_X1 U611 ( .A1(n551), .A2(n568), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  NAND2_X1 U614 ( .A1(n551), .A2(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n576), .A2(n551), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G169GAT), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT119), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n559) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n562) );
  NOR2_X1 U627 ( .A1(n554), .A2(n560), .ZN(n561) );
  XOR2_X1 U628 ( .A(n562), .B(n561), .Z(G1351GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n572) );
  XOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .Z(n570) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT123), .ZN(n580) );
  NAND2_X1 U635 ( .A1(n580), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n575) );
  NAND2_X1 U639 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(G1353GAT) );
  XOR2_X1 U641 ( .A(G211GAT), .B(KEYINPUT127), .Z(n578) );
  NAND2_X1 U642 ( .A1(n580), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1354GAT) );
  NAND2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(KEYINPUT62), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

