//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT23), .B1(new_n187), .B2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT76), .B1(new_n189), .B2(G128), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n188), .B(new_n190), .Z(new_n191));
  XNOR2_X1  g005(.A(G119), .B(G128), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT24), .B(G110), .Z(new_n193));
  OAI22_X1  g007(.A1(new_n191), .A2(G110), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G125), .B(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT16), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  OR3_X1    g011(.A1(new_n197), .A2(KEYINPUT16), .A3(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(G146), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n194), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n196), .A2(new_n198), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n200), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n199), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n193), .A2(new_n192), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n191), .A2(G110), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G137), .ZN(new_n210));
  INV_X1    g024(.A(G953), .ZN(new_n211));
  AND3_X1   g025(.A1(new_n211), .A2(G221), .A3(G234), .ZN(new_n212));
  XOR2_X1   g026(.A(new_n210), .B(new_n212), .Z(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G902), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n202), .A2(new_n208), .A3(new_n213), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(new_n218), .B(KEYINPUT25), .Z(new_n219));
  INV_X1    g033(.A(G217), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(G234), .B2(new_n216), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n215), .A2(new_n217), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n221), .A2(G902), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT73), .ZN(new_n228));
  INV_X1    g042(.A(G472), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n216), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT2), .B(G113), .Z(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n200), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n238), .B(KEYINPUT1), .C1(new_n235), .C2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G128), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n237), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n234), .A3(new_n236), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n247), .A3(new_n244), .ZN(new_n248));
  INV_X1    g062(.A(G137), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT66), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G137), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT11), .A2(G134), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G131), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT11), .A2(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G137), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT11), .A2(G134), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n254), .A2(new_n255), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n250), .A2(new_n252), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n255), .B1(G134), .B2(G137), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n246), .A2(new_n248), .A3(new_n264), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n257), .B1(KEYINPUT11), .B2(G134), .ZN(new_n267));
  OAI21_X1  g081(.A(G131), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n259), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n234), .A2(new_n236), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G143), .B(G146), .ZN(new_n274));
  NOR3_X1   g088(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n265), .A2(KEYINPUT30), .A3(new_n278), .ZN(new_n279));
  OR3_X1    g093(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n237), .A2(new_n280), .B1(KEYINPUT0), .B2(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT65), .B1(new_n281), .B2(new_n272), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT65), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(new_n283), .A3(new_n276), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n269), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n264), .A2(new_n245), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n288));
  AOI21_X1  g102(.A(KEYINPUT68), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  AOI211_X1 g104(.A(new_n290), .B(KEYINPUT30), .C1(new_n285), .C2(new_n286), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n233), .B(new_n279), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n233), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n265), .A2(new_n293), .A3(new_n278), .ZN(new_n294));
  NOR2_X1   g108(.A1(G237), .A2(G953), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G210), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT27), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT26), .B(G101), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n294), .A2(KEYINPUT70), .A3(new_n299), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n292), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n292), .A2(new_n302), .A3(KEYINPUT31), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n294), .A2(KEYINPUT72), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n287), .A2(new_n233), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n294), .B2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT72), .B1(new_n294), .B2(new_n309), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(new_n299), .B(KEYINPUT71), .Z(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n230), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n228), .B1(new_n319), .B2(KEYINPUT32), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT32), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n306), .A2(new_n307), .B1(new_n316), .B2(new_n317), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT73), .B(new_n321), .C1(new_n322), .C2(new_n230), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n322), .A2(new_n321), .A3(new_n230), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n311), .B2(new_n314), .ZN(new_n327));
  INV_X1    g141(.A(new_n314), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(KEYINPUT75), .A3(new_n310), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n265), .A2(new_n278), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n233), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n294), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT28), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n299), .A2(KEYINPUT29), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n292), .A2(new_n294), .ZN(new_n337));
  INV_X1    g151(.A(new_n299), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n317), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n315), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n337), .A2(KEYINPUT74), .A3(new_n338), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n345), .A3(new_n216), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n325), .B1(G472), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n227), .B1(new_n324), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(G214), .B1(G237), .B2(G902), .ZN(new_n349));
  OAI21_X1  g163(.A(G210), .B1(G237), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT78), .B1(new_n352), .B2(G104), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  INV_X1    g168(.A(G104), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G107), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n352), .A2(KEYINPUT3), .A3(G104), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n352), .B2(G104), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n353), .B(new_n356), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n355), .B2(G107), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n352), .A2(KEYINPUT3), .A3(G104), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n353), .A4(new_n356), .ZN(new_n366));
  XOR2_X1   g180(.A(KEYINPUT80), .B(KEYINPUT4), .Z(new_n367));
  NAND4_X1  g181(.A1(new_n361), .A2(G101), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n233), .ZN(new_n369));
  INV_X1    g183(.A(G101), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n365), .A2(new_n370), .A3(new_n353), .A4(new_n356), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n359), .B2(new_n360), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n366), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT84), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n189), .A2(G116), .ZN(new_n376));
  OAI21_X1  g190(.A(G113), .B1(new_n376), .B2(KEYINPUT5), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(KEYINPUT5), .B2(new_n232), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(new_n232), .B2(new_n231), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n352), .A2(G104), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n355), .A2(G107), .ZN(new_n381));
  OAI21_X1  g195(.A(G101), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n361), .A2(G101), .A3(new_n366), .ZN(new_n386));
  AND2_X1   g200(.A1(new_n371), .A2(KEYINPUT4), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n368), .A4(new_n233), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n375), .A2(new_n385), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(G110), .B(G122), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n392), .B(KEYINPUT8), .ZN(new_n396));
  INV_X1    g210(.A(new_n385), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n379), .A2(new_n384), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n277), .A2(G125), .ZN(new_n400));
  INV_X1    g214(.A(new_n245), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n400), .B1(new_n401), .B2(G125), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n211), .A2(G224), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT7), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT7), .ZN(new_n405));
  AOI22_X1  g219(.A1(KEYINPUT87), .A2(new_n405), .B1(new_n211), .B2(G224), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(KEYINPUT87), .B2(new_n405), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n400), .B(new_n407), .C1(new_n401), .C2(G125), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n399), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(G902), .B1(new_n395), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n391), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n375), .A2(new_n390), .A3(KEYINPUT85), .A4(new_n385), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n392), .A2(KEYINPUT6), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n413), .A2(KEYINPUT86), .A3(new_n414), .A4(new_n415), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n414), .A3(new_n393), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n394), .A2(new_n421), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n418), .A2(new_n419), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n402), .B(new_n403), .ZN(new_n424));
  AOI211_X1 g238(.A(new_n351), .B(new_n411), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n418), .A2(new_n419), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n420), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n424), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n350), .B1(new_n428), .B2(new_n410), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n349), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G469), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n368), .A2(new_n277), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n187), .B1(new_n234), .B2(KEYINPUT1), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n244), .B1(new_n433), .B2(new_n274), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n371), .A3(new_n382), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n434), .A2(new_n371), .A3(KEYINPUT81), .A4(new_n382), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n388), .A2(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n269), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n246), .A2(KEYINPUT10), .A3(new_n248), .A4(new_n384), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n441), .A2(KEYINPUT82), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n440), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n388), .A2(new_n277), .A3(new_n368), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n445), .A2(new_n442), .A3(new_n446), .A4(new_n443), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n211), .A2(G227), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT77), .ZN(new_n452));
  XNOR2_X1  g266(.A(G110), .B(G140), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n445), .A2(new_n443), .A3(new_n446), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n269), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n450), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n401), .A2(new_n383), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n439), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT12), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n460), .A3(new_n269), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n437), .A2(new_n438), .B1(new_n401), .B2(new_n383), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT12), .B1(new_n462), .B2(new_n442), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n464), .B1(new_n444), .B2(new_n449), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n457), .B1(new_n465), .B2(new_n454), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n431), .B1(new_n466), .B2(new_n216), .ZN(new_n467));
  INV_X1    g281(.A(new_n454), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n468), .B(new_n464), .C1(new_n449), .C2(new_n444), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n454), .B1(new_n450), .B2(new_n456), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n431), .B(new_n216), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n465), .A2(new_n454), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n444), .A2(new_n449), .B1(new_n269), .B2(new_n455), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n454), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n476), .A2(KEYINPUT83), .A3(new_n431), .A4(new_n216), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n467), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G221), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT9), .B(G234), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n481), .B2(new_n216), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n430), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(G113), .B(G122), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(new_n355), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n295), .A2(G143), .A3(G214), .ZN(new_n486));
  AOI21_X1  g300(.A(G143), .B1(new_n295), .B2(G214), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G131), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n255), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n195), .B(KEYINPUT19), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n200), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n199), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT18), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n488), .B1(new_n496), .B2(new_n255), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n195), .B(new_n200), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(KEYINPUT18), .A3(G131), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n485), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n489), .A2(KEYINPUT17), .A3(G131), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n503), .A2(new_n204), .A3(new_n199), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n490), .A2(new_n491), .A3(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n504), .A2(new_n506), .B1(new_n500), .B2(new_n499), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n502), .B1(new_n507), .B2(new_n485), .ZN(new_n508));
  NOR2_X1   g322(.A1(G475), .A2(G902), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT20), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n504), .A2(new_n506), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n485), .A3(new_n501), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n512), .B(new_n509), .C1(new_n515), .C2(new_n502), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n507), .A2(new_n485), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n216), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n511), .A2(new_n516), .B1(new_n518), .B2(G475), .ZN(new_n519));
  INV_X1    g333(.A(G952), .ZN(new_n520));
  AOI211_X1 g334(.A(G953), .B(new_n520), .C1(G234), .C2(G237), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n216), .B(new_n211), .C1(G234), .C2(G237), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n235), .A2(G128), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT13), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n187), .A2(G143), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  OAI21_X1  g345(.A(G134), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(new_n529), .A3(new_n260), .ZN(new_n533));
  XNOR2_X1  g347(.A(G116), .B(G122), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(new_n352), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n534), .A2(new_n352), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n532), .B(new_n533), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n480), .A2(new_n220), .A3(G953), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n526), .A2(new_n529), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G134), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n540), .A2(KEYINPUT88), .A3(new_n533), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT88), .B1(new_n540), .B2(new_n533), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n536), .A2(KEYINPUT89), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT14), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G116), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT14), .A3(G122), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n546), .A2(G107), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n534), .A2(new_n352), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT89), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n544), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n537), .B(new_n538), .C1(new_n543), .C2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n537), .B1(new_n543), .B2(new_n553), .ZN(new_n558));
  INV_X1    g372(.A(new_n538), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n216), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT15), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(new_n563), .A3(G478), .ZN(new_n564));
  INV_X1    g378(.A(G478), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n561), .B(new_n216), .C1(KEYINPUT15), .C2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n519), .A2(new_n525), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT91), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n348), .A2(new_n483), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  INV_X1    g385(.A(new_n349), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n428), .A2(new_n410), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n351), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n428), .A2(new_n410), .A3(new_n350), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n558), .B2(new_n559), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n561), .A2(new_n577), .B1(new_n578), .B2(new_n554), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n565), .A2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT92), .B(G478), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n562), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n511), .A2(new_n516), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n518), .A2(G475), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n576), .A2(new_n525), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G472), .B1(new_n322), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n319), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR4_X1   g408(.A1(new_n478), .A2(new_n594), .A3(new_n482), .A4(new_n227), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT34), .B(G104), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G6));
  NAND2_X1  g412(.A1(new_n564), .A2(new_n566), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n519), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n576), .A2(new_n525), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n595), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  NOR2_X1   g419(.A1(new_n214), .A2(KEYINPUT36), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n209), .B(new_n606), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n219), .A2(new_n221), .B1(new_n224), .B2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n568), .A2(new_n594), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n483), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT93), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT37), .B(G110), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G12));
  XOR2_X1   g427(.A(KEYINPUT94), .B(G900), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n522), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n521), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n600), .A2(new_n617), .ZN(new_n618));
  NOR4_X1   g432(.A1(new_n430), .A2(new_n478), .A3(new_n482), .A4(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n608), .B1(new_n324), .B2(new_n347), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G128), .ZN(G30));
  NAND2_X1  g436(.A1(new_n574), .A2(new_n575), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT38), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n229), .B1(new_n332), .B2(new_n317), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n304), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(G472), .A2(G902), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n628), .B(KEYINPUT95), .Z(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n325), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n324), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n519), .B1(new_n564), .B2(new_n566), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n632), .A2(new_n349), .A3(new_n608), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n624), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n478), .A2(new_n482), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n617), .B(KEYINPUT39), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT40), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n634), .A2(KEYINPUT96), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n631), .A2(new_n633), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n642), .A2(new_n640), .A3(new_n638), .A4(new_n624), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n235), .ZN(G45));
  NAND2_X1  g461(.A1(new_n346), .A2(G472), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n319), .A2(KEYINPUT32), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n320), .A3(new_n323), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n617), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n588), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n608), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n650), .A2(new_n635), .A3(new_n576), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT97), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n654), .B1(new_n324), .B2(new_n347), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT97), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n483), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT98), .B(G146), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G48));
  OAI21_X1  g477(.A(new_n216), .B1(new_n469), .B2(new_n470), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n476), .A2(KEYINPUT99), .A3(new_n216), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(G469), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n473), .A2(new_n477), .ZN(new_n669));
  INV_X1    g483(.A(new_n482), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n650), .A3(new_n226), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n590), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT41), .B(G113), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  INV_X1    g490(.A(new_n673), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n602), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT100), .B(G116), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G18));
  NAND3_X1  g494(.A1(new_n650), .A2(new_n569), .A3(new_n653), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n671), .A2(new_n430), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G119), .ZN(G21));
  NAND2_X1  g499(.A1(new_n576), .A2(new_n525), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n334), .A2(new_n317), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n308), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n230), .B(KEYINPUT101), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n592), .A3(new_n226), .A4(new_n632), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n686), .A2(new_n671), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(G122), .Z(G24));
  AND2_X1   g507(.A1(new_n668), .A2(new_n669), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n592), .A2(new_n652), .A3(new_n690), .A4(new_n653), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n695), .A3(new_n670), .A4(new_n576), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G125), .ZN(G27));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  AOI221_X4 g512(.A(new_n468), .B1(new_n269), .B2(new_n455), .C1(new_n444), .C2(new_n449), .ZN(new_n699));
  INV_X1    g513(.A(new_n464), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n454), .B1(new_n450), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n698), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n457), .A2(KEYINPUT102), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(G469), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT103), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n431), .A2(new_n216), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n702), .A2(new_n708), .A3(G469), .A4(new_n703), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n669), .A2(new_n705), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT104), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n706), .B1(new_n473), .B2(new_n477), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n709), .A4(new_n705), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n670), .A2(new_n349), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n623), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n348), .A3(new_n652), .A4(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n719));
  NAND2_X1  g533(.A1(new_n593), .A2(new_n321), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n649), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n319), .A2(KEYINPUT32), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT106), .B1(new_n723), .B2(new_n325), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n724), .A3(new_n648), .ZN(new_n725));
  AND4_X1   g539(.A1(KEYINPUT42), .A2(new_n725), .A3(new_n226), .A4(new_n652), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n623), .A2(new_n716), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n714), .B2(new_n711), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n718), .A2(new_n719), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n255), .ZN(G33));
  INV_X1    g544(.A(new_n618), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n715), .A2(new_n348), .A3(new_n731), .A4(new_n717), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G134), .ZN(G36));
  AOI22_X1  g547(.A1(new_n579), .A2(new_n580), .B1(new_n562), .B2(new_n582), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n587), .A2(new_n734), .A3(KEYINPUT43), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n584), .B2(new_n519), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT108), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n587), .B2(new_n734), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n584), .A2(new_n519), .A3(new_n736), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT44), .A3(new_n594), .A4(new_n653), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n623), .A2(new_n572), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT109), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n744), .A2(new_n748), .A3(new_n745), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n743), .A2(new_n594), .A3(new_n653), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n747), .A2(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n702), .A2(KEYINPUT45), .A3(new_n703), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n431), .B1(new_n466), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n707), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n706), .B1(new_n753), .B2(new_n755), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n669), .B1(new_n760), .B2(KEYINPUT46), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n670), .B(new_n637), .C1(new_n759), .C2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n752), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  NAND2_X1  g581(.A1(new_n227), .A2(new_n652), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n650), .A2(new_n623), .A3(new_n768), .A4(new_n572), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT110), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n772));
  OAI221_X1 g586(.A(new_n670), .B1(new_n771), .B2(new_n772), .C1(new_n759), .C2(new_n761), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n759), .A2(new_n761), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n482), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n769), .B(new_n773), .C1(new_n775), .C2(new_n772), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NAND2_X1  g591(.A1(new_n668), .A2(new_n669), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT111), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT49), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n631), .A2(new_n227), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n624), .A2(new_n587), .A3(new_n734), .A4(new_n716), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n478), .A2(new_n599), .A3(new_n587), .A4(new_n651), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n620), .A2(new_n717), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n732), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n728), .A2(new_n695), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n728), .A2(KEYINPUT114), .A3(new_n695), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n729), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n619), .A2(new_n620), .B1(new_n683), .B2(new_n695), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n651), .A2(new_n482), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n632), .A2(new_n608), .A3(new_n796), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(new_n349), .C1(new_n425), .C2(new_n429), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n324), .B2(new_n630), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n715), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n661), .A2(new_n794), .A3(new_n795), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n656), .A2(KEYINPUT97), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n659), .B1(new_n658), .B2(new_n483), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n795), .B(new_n800), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n792), .A2(new_n793), .A3(new_n801), .A4(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n590), .A2(KEYINPUT113), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n590), .A2(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n595), .A3(new_n808), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n570), .A2(new_n809), .A3(new_n610), .A4(new_n603), .ZN(new_n810));
  INV_X1    g624(.A(new_n683), .ZN(new_n811));
  OAI22_X1  g625(.A1(new_n673), .A2(new_n601), .B1(new_n811), .B2(new_n681), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n671), .A2(new_n691), .ZN(new_n813));
  OAI22_X1  g627(.A1(new_n673), .A2(new_n590), .B1(new_n813), .B2(new_n686), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT112), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n812), .A2(new_n814), .A3(KEYINPUT112), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n810), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n784), .B1(new_n806), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n805), .A2(new_n801), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n728), .A2(KEYINPUT114), .A3(new_n695), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT114), .B1(new_n728), .B2(new_n695), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n824), .A2(new_n729), .A3(new_n787), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n812), .A2(new_n814), .A3(new_n784), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n635), .A2(new_n576), .A3(new_n731), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n650), .A2(new_n653), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n696), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT52), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n821), .A2(new_n825), .A3(new_n810), .A4(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n819), .A2(new_n820), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n809), .A2(new_n610), .A3(new_n570), .A4(new_n603), .ZN(new_n834));
  INV_X1    g648(.A(new_n814), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n836), .A3(new_n678), .A4(new_n684), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n834), .B1(new_n837), .B2(new_n815), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n830), .A2(new_n784), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n821), .A2(new_n825), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n820), .B1(new_n819), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n623), .B(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n592), .A2(new_n690), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n735), .A2(new_n737), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n226), .A2(new_n844), .A3(new_n521), .A4(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n843), .A2(new_n572), .A3(new_n846), .A4(new_n672), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(KEYINPUT50), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n727), .A2(new_n616), .A3(new_n778), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(new_n519), .A3(new_n734), .A4(new_n781), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n845), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n653), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n775), .A2(new_n772), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n773), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n779), .A2(new_n482), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n846), .A2(new_n745), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n854), .B(KEYINPUT51), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n848), .A2(new_n853), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n856), .B2(new_n857), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n725), .A2(new_n226), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n849), .A2(new_n865), .A3(new_n845), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT48), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n849), .A2(new_n589), .A3(new_n781), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n520), .B(G953), .C1(new_n846), .C2(new_n683), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n860), .A2(new_n864), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n833), .A2(new_n841), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n783), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT115), .B(new_n783), .C1(new_n872), .C2(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(G75));
  XNOR2_X1  g692(.A(new_n423), .B(new_n424), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT55), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n819), .A2(new_n832), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n881), .A2(G210), .A3(G902), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n882), .B2(KEYINPUT56), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n211), .A2(G952), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n882), .A2(KEYINPUT56), .A3(new_n880), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(G51));
  XNOR2_X1  g702(.A(new_n706), .B(KEYINPUT57), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n820), .B1(new_n819), .B2(new_n832), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n889), .B1(new_n833), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT116), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n893), .B(new_n889), .C1(new_n833), .C2(new_n890), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n476), .B(KEYINPUT117), .Z(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n881), .A2(G902), .A3(new_n753), .A4(new_n755), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n884), .B1(new_n896), .B2(new_n897), .ZN(G54));
  NAND4_X1  g712(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(new_n508), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n508), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n884), .ZN(G60));
  OR2_X1    g716(.A1(new_n833), .A2(new_n841), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n565), .A2(new_n216), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n579), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n579), .B(new_n906), .C1(new_n833), .C2(new_n890), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n885), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(G63));
  NAND2_X1  g724(.A1(G217), .A2(G902), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT119), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT60), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n881), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n223), .B(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n881), .A2(new_n607), .A3(new_n913), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n885), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G66));
  INV_X1    g734(.A(G224), .ZN(new_n921));
  OAI21_X1  g735(.A(G953), .B1(new_n523), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT121), .Z(new_n923));
  OAI21_X1  g737(.A(new_n923), .B1(new_n838), .B2(G953), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  INV_X1    g739(.A(G898), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n423), .B1(new_n926), .B2(G953), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n925), .B(new_n927), .ZN(G69));
  OAI21_X1  g742(.A(new_n279), .B1(new_n289), .B2(new_n291), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT123), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n493), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(G900), .B(G953), .C1(new_n932), .C2(G227), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(G227), .B2(new_n932), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n829), .B1(new_n660), .B2(new_n657), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n793), .A2(new_n732), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n766), .A2(new_n776), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n576), .A2(new_n632), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n865), .B(new_n938), .C1(new_n764), .C2(new_n765), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(G953), .B1(new_n940), .B2(new_n932), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n641), .A2(new_n645), .A3(new_n935), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  INV_X1    g757(.A(new_n639), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n589), .A2(new_n600), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n944), .A2(new_n348), .A3(new_n745), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n766), .A2(new_n776), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n942), .A2(new_n949), .A3(KEYINPUT62), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n949), .B1(new_n942), .B2(KEYINPUT62), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n931), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n934), .B1(new_n941), .B2(new_n953), .ZN(G72));
  XNOR2_X1  g768(.A(new_n627), .B(KEYINPUT63), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n337), .B(KEYINPUT125), .Z(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n299), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n299), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n955), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n885), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n948), .B(new_n957), .C1(new_n950), .C2(new_n951), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n936), .A2(new_n937), .A3(new_n939), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n963), .B2(new_n838), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n819), .A2(new_n840), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n341), .A2(new_n344), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n955), .B1(new_n966), .B2(new_n304), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT126), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n965), .A2(KEYINPUT126), .A3(new_n967), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n964), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT127), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT127), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n964), .B(new_n972), .C1(new_n968), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n973), .ZN(G57));
endmodule


