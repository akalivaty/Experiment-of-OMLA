//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n193), .A3(new_n196), .A4(new_n191), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n200), .A2(new_n202), .A3(G128), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n200), .B2(new_n202), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT0), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G128), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n198), .A2(KEYINPUT67), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G128), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n199), .B(G146), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n200), .A2(new_n202), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n211), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n192), .A2(KEYINPUT64), .A3(G134), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n191), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT64), .B1(new_n192), .B2(G134), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n197), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n200), .A2(new_n202), .A3(G128), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n226), .B1(new_n210), .B2(new_n204), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n227), .A2(KEYINPUT0), .B1(G128), .B2(new_n205), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT67), .B1(new_n228), .B2(new_n198), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT30), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n197), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n223), .A2(KEYINPUT65), .A3(new_n197), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n219), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n228), .A2(new_n198), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G116), .B(G119), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT68), .A2(G953), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT68), .A2(G953), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G237), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(G210), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT27), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n225), .A2(new_n229), .A3(new_n243), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n244), .A2(new_n255), .A3(KEYINPUT31), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT31), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n242), .B1(new_n230), .B2(new_n238), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n237), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(new_n242), .A3(new_n224), .A4(new_n208), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n252), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n242), .B1(new_n235), .B2(new_n237), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT28), .B1(new_n254), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g079(.A1(new_n224), .A2(new_n242), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT28), .B1(new_n266), .B2(new_n237), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n256), .A2(new_n263), .B1(new_n253), .B2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(G472), .A2(G902), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n187), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(new_n253), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT31), .B1(new_n244), .B2(new_n255), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n258), .A2(new_n262), .A3(new_n257), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT69), .A3(new_n271), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n273), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(KEYINPUT32), .A3(new_n271), .ZN(new_n281));
  INV_X1    g095(.A(G472), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n253), .B1(new_n258), .B2(new_n254), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n265), .A2(new_n252), .A3(new_n268), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n243), .B1(new_n225), .B2(new_n229), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n261), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n267), .B1(new_n288), .B2(KEYINPUT28), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n253), .A2(new_n285), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g105(.A(KEYINPUT70), .B(new_n282), .C1(new_n286), .C2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n291), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(G472), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n280), .B(new_n281), .C1(new_n292), .C2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G475), .A2(G902), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G125), .ZN(new_n299));
  INV_X1    g113(.A(G125), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G140), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n301), .A3(KEYINPUT71), .ZN(new_n302));
  OR3_X1    g116(.A1(new_n300), .A2(KEYINPUT71), .A3(G140), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT16), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT16), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n304), .A2(new_n201), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n201), .B1(new_n304), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OR2_X1    g123(.A1(KEYINPUT68), .A2(G953), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT68), .A2(G953), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n310), .A2(G214), .A3(new_n248), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n199), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n247), .A2(G143), .A3(G214), .A4(new_n248), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT17), .A3(G131), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(G131), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n314), .A3(new_n196), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n309), .B(new_n316), .C1(new_n319), .C2(KEYINPUT17), .ZN(new_n320));
  XNOR2_X1  g134(.A(G113), .B(G122), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT96), .B(G104), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(KEYINPUT18), .A2(G131), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n315), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT95), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n313), .A2(new_n314), .A3(new_n324), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n299), .A2(new_n301), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n201), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n302), .A2(new_n303), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(new_n201), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n315), .A2(KEYINPUT95), .A3(new_n325), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n328), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n320), .A2(new_n323), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n330), .A2(KEYINPUT19), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n308), .B1(new_n340), .B2(new_n201), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n319), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n323), .B1(new_n336), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT97), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n337), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT95), .B1(new_n315), .B2(new_n325), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n329), .A2(new_n333), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n348), .A2(new_n335), .B1(new_n341), .B2(new_n319), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n349), .A2(KEYINPUT97), .A3(new_n323), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n297), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(KEYINPUT20), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n353), .B(new_n297), .C1(new_n345), .C2(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n320), .A2(new_n336), .ZN(new_n355));
  INV_X1    g169(.A(new_n323), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT98), .A3(new_n337), .ZN(new_n358));
  INV_X1    g172(.A(G902), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n360), .A3(new_n356), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n352), .A2(new_n354), .B1(new_n362), .B2(G475), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT9), .B(G234), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT78), .ZN(new_n365));
  INV_X1    g179(.A(G953), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(KEYINPUT78), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n365), .A2(G217), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G116), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(G122), .ZN(new_n371));
  INV_X1    g185(.A(G122), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G116), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT80), .A2(G107), .ZN(new_n374));
  AND2_X1   g188(.A1(KEYINPUT80), .A2(G107), .ZN(new_n375));
  OAI22_X1  g189(.A1(new_n371), .A2(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OR2_X1    g190(.A1(KEYINPUT80), .A2(G107), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(G116), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n370), .A2(G122), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT80), .A2(G107), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n376), .A2(KEYINPUT99), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT99), .B1(new_n376), .B2(new_n381), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n199), .A2(G128), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n217), .A2(G143), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT13), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n199), .B2(G128), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(G134), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n384), .B(new_n385), .C1(new_n387), .C2(new_n189), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n382), .A2(new_n383), .A3(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT14), .B1(new_n372), .B2(G116), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n370), .A3(G122), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n395), .A3(new_n378), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n396), .A2(G107), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(new_n189), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n384), .A2(new_n385), .A3(G134), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n381), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n369), .B1(new_n392), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n376), .A2(new_n381), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n376), .A2(KEYINPUT99), .A3(new_n381), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n389), .A4(new_n390), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n397), .A2(new_n400), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n368), .A3(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n402), .A2(new_n359), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT100), .ZN(new_n411));
  INV_X1    g225(.A(G478), .ZN(new_n412));
  NOR2_X1   g226(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(KEYINPUT101), .A2(KEYINPUT15), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT100), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n402), .A2(new_n409), .A3(new_n417), .A4(new_n359), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n410), .A2(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n363), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G952), .ZN(new_n424));
  AOI211_X1 g238(.A(G953), .B(new_n424), .C1(G234), .C2(G237), .ZN(new_n425));
  AOI211_X1 g239(.A(new_n359), .B(new_n247), .C1(G234), .C2(G237), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(G898), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G217), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n430), .B1(G234), .B2(new_n359), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n433), .B2(KEYINPUT75), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT22), .B(G137), .Z(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT74), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n247), .A2(G221), .A3(G234), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT73), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT23), .ZN(new_n441));
  INV_X1    g255(.A(G119), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(G128), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n443), .B(new_n444), .C1(G119), .C2(new_n217), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G110), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT24), .B(G110), .Z(new_n447));
  XNOR2_X1  g261(.A(G119), .B(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n304), .A2(new_n306), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G146), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n304), .A2(new_n201), .A3(new_n306), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT72), .B(G110), .Z(new_n455));
  OAI22_X1  g269(.A1(new_n445), .A2(new_n455), .B1(new_n448), .B2(new_n447), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n331), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n308), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n440), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n449), .B(new_n446), .C1(new_n307), .C2(new_n308), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n452), .A2(new_n331), .A3(new_n456), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT73), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n439), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n438), .B1(new_n460), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n434), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n433), .A2(KEYINPUT75), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n432), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI221_X1 g281(.A(new_n434), .B1(KEYINPUT75), .B2(new_n433), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OR3_X1    g283(.A1(new_n463), .A2(KEYINPUT76), .A3(new_n464), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n432), .A2(new_n359), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT77), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT76), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n296), .A2(new_n429), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT4), .ZN(new_n478));
  INV_X1    g292(.A(G101), .ZN(new_n479));
  INV_X1    g293(.A(G107), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT81), .B1(new_n480), .B2(G104), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT81), .ZN(new_n482));
  INV_X1    g296(.A(G104), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(G107), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(G104), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n481), .A2(new_n484), .B1(new_n485), .B2(KEYINPUT3), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n483), .A2(KEYINPUT3), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n377), .A3(new_n380), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n479), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n242), .B1(new_n478), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n481), .A2(new_n484), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n485), .A2(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT82), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(G101), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT83), .B(G101), .Z(new_n496));
  NAND4_X1  g310(.A1(new_n496), .A2(new_n488), .A3(new_n491), .A4(new_n492), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n493), .B2(G101), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(G104), .B1(new_n377), .B2(new_n380), .ZN(new_n501));
  INV_X1    g315(.A(new_n485), .ZN(new_n502));
  OAI21_X1  g316(.A(G101), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n240), .A2(KEYINPUT5), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n370), .A2(KEYINPUT5), .A3(G119), .ZN(new_n505));
  INV_X1    g319(.A(G113), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n241), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n240), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n497), .A2(new_n503), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G110), .B(G122), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n219), .A2(new_n300), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n206), .A2(new_n207), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(new_n300), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n366), .A2(G224), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n516), .A2(KEYINPUT92), .A3(KEYINPUT7), .A4(new_n520), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n513), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n497), .A2(new_n503), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n508), .A2(new_n510), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(new_n511), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n512), .B(KEYINPUT8), .Z(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT91), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n532));
  AOI211_X1 g346(.A(new_n532), .B(new_n529), .C1(new_n527), .C2(new_n511), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n359), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT93), .B(new_n359), .C1(new_n524), .C2(new_n534), .ZN(new_n538));
  INV_X1    g352(.A(new_n512), .ZN(new_n539));
  INV_X1    g353(.A(new_n500), .ZN(new_n540));
  INV_X1    g354(.A(new_n511), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(KEYINPUT6), .A3(new_n513), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n516), .B(new_n520), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n537), .A2(new_n538), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n537), .A2(new_n547), .A3(new_n549), .A4(new_n538), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(KEYINPUT94), .A3(new_n552), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n552), .A2(KEYINPUT94), .ZN(new_n554));
  OAI21_X1  g368(.A(G214), .B1(G237), .B2(G902), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT90), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G221), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT78), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n364), .B(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n561), .B2(new_n359), .ZN(new_n562));
  INV_X1    g376(.A(G469), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n211), .B(new_n218), .C1(new_n212), .C2(new_n200), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n497), .A3(new_n503), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n497), .A2(new_n503), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(new_n219), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT86), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n568), .A2(KEYINPUT85), .A3(KEYINPUT12), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(KEYINPUT86), .B2(new_n567), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT85), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n572), .A3(new_n198), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n571), .A2(new_n198), .B1(KEYINPUT12), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n247), .A2(G227), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT79), .ZN(new_n576));
  XNOR2_X1  g390(.A(G110), .B(G140), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT84), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n566), .A2(new_n579), .A3(KEYINPUT10), .A4(new_n219), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n219), .A2(KEYINPUT10), .A3(new_n497), .A4(new_n503), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT84), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n489), .A2(new_n478), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n584), .B(new_n228), .C1(new_n498), .C2(new_n499), .ZN(new_n585));
  INV_X1    g399(.A(new_n198), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n565), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n583), .A2(new_n585), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n574), .A2(new_n578), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT88), .ZN(new_n591));
  AOI211_X1 g405(.A(KEYINPUT82), .B(new_n479), .C1(new_n486), .C2(new_n488), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n592), .A2(new_n499), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n228), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n581), .B(new_n579), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n583), .A2(new_n585), .A3(KEYINPUT88), .A4(new_n588), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(new_n198), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n578), .B1(new_n600), .B2(new_n589), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT89), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n590), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n589), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n583), .A2(new_n585), .A3(new_n588), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n586), .B1(new_n605), .B2(new_n591), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n604), .B1(new_n606), .B2(new_n599), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n607), .A2(KEYINPUT89), .A3(new_n578), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n563), .B(new_n359), .C1(new_n603), .C2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n563), .A2(new_n359), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n578), .B1(new_n574), .B2(new_n589), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT87), .B1(new_n589), .B2(new_n578), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n612), .B1(new_n599), .B2(new_n606), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n589), .A2(KEYINPUT87), .A3(new_n578), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n610), .B1(new_n615), .B2(G469), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n562), .B1(new_n609), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n558), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n477), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n496), .ZN(G3));
  AND3_X1   g434(.A1(new_n357), .A2(KEYINPUT98), .A3(new_n337), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n361), .A2(new_n359), .ZN(new_n622));
  OAI21_X1  g436(.A(G475), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n354), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT97), .B1(new_n349), .B2(new_n323), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n336), .A2(new_n342), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n626), .A2(new_n344), .A3(new_n356), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n625), .A2(new_n337), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n353), .B1(new_n628), .B2(new_n297), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n623), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n368), .A2(KEYINPUT103), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n631), .B1(new_n392), .B2(new_n401), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n368), .A2(KEYINPUT103), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n407), .A2(new_n408), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(KEYINPUT33), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT102), .B(KEYINPUT33), .Z(new_n636));
  NAND3_X1  g450(.A1(new_n402), .A2(new_n409), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n412), .A2(G902), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n411), .A2(new_n412), .A3(new_n418), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n635), .A2(new_n637), .A3(KEYINPUT104), .A4(new_n638), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT105), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT105), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n641), .A2(new_n642), .A3(new_n646), .A4(new_n643), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n630), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT106), .ZN(new_n650));
  INV_X1    g464(.A(new_n555), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n651), .B1(new_n551), .B2(new_n552), .ZN(new_n652));
  INV_X1    g466(.A(new_n428), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n270), .B2(G902), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n273), .A2(new_n656), .A3(new_n278), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n475), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n617), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT34), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  NAND2_X1  g476(.A1(new_n363), .A2(new_n421), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n659), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT35), .B(G107), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n459), .A2(new_n462), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT36), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n439), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n459), .B(new_n462), .C1(KEYINPUT36), .C2(new_n438), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n671), .A2(new_n472), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n469), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n363), .A2(new_n675), .A3(new_n653), .A4(new_n422), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n657), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n558), .A2(new_n677), .A3(new_n617), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n426), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT107), .ZN(new_n683));
  INV_X1    g497(.A(new_n425), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(KEYINPUT107), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n663), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n673), .B1(new_n467), .B2(new_n468), .ZN(new_n689));
  AOI211_X1 g503(.A(new_n651), .B(new_n689), .C1(new_n551), .C2(new_n552), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n296), .A2(new_n617), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G128), .ZN(G30));
  XNOR2_X1  g506(.A(new_n686), .B(KEYINPUT39), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n617), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n694), .A2(KEYINPUT40), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n553), .A2(new_n554), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT38), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n258), .A2(new_n254), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n253), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n359), .B1(new_n288), .B2(new_n252), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n280), .A2(new_n281), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n352), .A2(new_n354), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n422), .B1(new_n704), .B2(new_n623), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n703), .A2(new_n555), .A3(new_n689), .A4(new_n705), .ZN(new_n706));
  NOR4_X1   g520(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT108), .B(G143), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G45));
  AND3_X1   g523(.A1(new_n296), .A2(new_n617), .A3(new_n690), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n630), .A2(new_n648), .A3(new_n686), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n630), .A2(new_n648), .A3(KEYINPUT109), .A4(new_n686), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  INV_X1    g532(.A(new_n609), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT89), .B1(new_n607), .B2(new_n578), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n600), .A2(new_n589), .ZN(new_n721));
  INV_X1    g535(.A(new_n578), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n602), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n720), .A2(new_n723), .A3(new_n590), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n563), .B1(new_n724), .B2(new_n359), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n562), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n476), .A4(new_n296), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n655), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT41), .B(G113), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NOR2_X1   g545(.A1(new_n728), .A2(new_n665), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n370), .ZN(G18));
  NAND3_X1  g547(.A1(new_n296), .A2(new_n429), .A3(new_n675), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n359), .B1(new_n603), .B2(new_n608), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(G469), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(new_n727), .A3(new_n609), .A4(new_n652), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n442), .ZN(G21));
  NAND2_X1  g553(.A1(new_n551), .A2(new_n552), .ZN(new_n740));
  AND4_X1   g554(.A1(new_n740), .A2(new_n705), .A3(new_n555), .A4(new_n653), .ZN(new_n741));
  OAI22_X1  g555(.A1(new_n275), .A2(new_n276), .B1(new_n252), .B2(new_n289), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n271), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n656), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n475), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n469), .A2(KEYINPUT110), .A3(new_n474), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n726), .A2(new_n741), .A3(new_n727), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G122), .ZN(G24));
  AND3_X1   g564(.A1(new_n675), .A2(new_n656), .A3(new_n743), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n713), .A2(new_n714), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n737), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n300), .ZN(G27));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n279), .B1(new_n270), .B2(new_n272), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n756), .B(new_n281), .C1(new_n295), .C2(new_n292), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n746), .A2(new_n747), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n713), .A2(new_n757), .A3(new_n758), .A4(new_n714), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n651), .B1(new_n553), .B2(new_n554), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n617), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n617), .A2(new_n760), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n280), .A2(new_n281), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n295), .A2(new_n292), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n476), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n713), .A2(new_n755), .A3(new_n714), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n763), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT111), .B1(new_n762), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n763), .A2(new_n766), .ZN(new_n770));
  INV_X1    g584(.A(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n757), .A2(new_n713), .A3(new_n714), .A4(new_n758), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT42), .B1(new_n763), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n196), .ZN(G33));
  INV_X1    g592(.A(new_n688), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n763), .A2(new_n766), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n189), .ZN(G36));
  NAND2_X1  g595(.A1(new_n657), .A2(new_n675), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g597(.A1(KEYINPUT112), .A2(KEYINPUT43), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n363), .A2(new_n648), .ZN(new_n786));
  MUX2_X1   g600(.A(new_n784), .B(new_n785), .S(new_n786), .Z(new_n787));
  NAND2_X1  g601(.A1(new_n783), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n760), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(G469), .B1(new_n615), .B2(KEYINPUT45), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(KEYINPUT45), .B2(new_n615), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(new_n794), .B2(new_n610), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n609), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n794), .A2(new_n792), .A3(new_n610), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n727), .B(new_n693), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n798), .B1(new_n789), .B2(new_n788), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n791), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(new_n296), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n716), .A2(new_n803), .A3(new_n475), .A4(new_n760), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n727), .B1(new_n796), .B2(new_n797), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(KEYINPUT47), .B(new_n727), .C1(new_n796), .C2(new_n797), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n298), .ZN(G42));
  AND2_X1   g624(.A1(new_n748), .A2(new_n425), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n787), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n719), .A2(new_n725), .A3(new_n562), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n698), .A2(new_n651), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n816), .B1(new_n814), .B2(new_n815), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n813), .A2(new_n425), .A3(new_n760), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(new_n787), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n817), .A2(new_n818), .B1(new_n751), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n726), .A2(new_n562), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n807), .A2(new_n808), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(new_n760), .A3(new_n812), .ZN(new_n824));
  INV_X1    g638(.A(new_n703), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n819), .A2(new_n476), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(KEYINPUT118), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n630), .A2(new_n648), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n821), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT51), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n757), .A2(new_n758), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n820), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n836));
  XNOR2_X1  g650(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n827), .A2(new_n650), .A3(new_n828), .ZN(new_n838));
  INV_X1    g652(.A(new_n737), .ZN(new_n839));
  AOI211_X1 g653(.A(new_n424), .B(G953), .C1(new_n812), .C2(new_n839), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n821), .A2(KEYINPUT51), .A3(new_n824), .A4(new_n830), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n833), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n687), .B(new_n673), .C1(new_n467), .C2(new_n468), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n652), .A2(new_n705), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n825), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n710), .A2(new_n716), .B1(new_n846), .B2(new_n617), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n617), .A2(new_n296), .A3(new_n688), .A4(new_n690), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n753), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT116), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n691), .B1(new_n737), .B2(new_n752), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n740), .A2(new_n705), .A3(new_n555), .A4(new_n844), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n617), .A3(new_n703), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n296), .A2(new_n617), .A3(new_n690), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n856), .B2(new_n715), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n852), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n851), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n728), .A2(new_n665), .B1(new_n737), .B2(new_n734), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n749), .B1(new_n728), .B2(new_n655), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT117), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n862), .B2(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n428), .B1(new_n663), .B2(new_n649), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n558), .A2(new_n617), .A3(new_n658), .A4(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n870), .B(new_n678), .C1(new_n618), .C2(new_n477), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT115), .B1(new_n423), .B2(new_n687), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n363), .A2(new_n873), .A3(new_n422), .A4(new_n686), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n296), .A2(new_n675), .A3(new_n872), .A4(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n763), .B1(new_n875), .B2(new_n752), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n871), .A2(new_n876), .A3(new_n780), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n762), .A2(new_n768), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n861), .A2(new_n868), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n877), .A2(new_n864), .A3(new_n769), .A4(new_n776), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT116), .B1(new_n847), .B2(new_n849), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n853), .A2(new_n857), .A3(new_n852), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT52), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n883), .B1(new_n886), .B2(new_n859), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n881), .B(new_n882), .C1(new_n887), .C2(KEYINPUT53), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n861), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n887), .B2(new_n878), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n891), .B2(new_n882), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n843), .A2(new_n892), .B1(G952), .B2(G953), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n726), .B(KEYINPUT49), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n758), .A2(new_n727), .A3(new_n557), .A4(new_n786), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n703), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n698), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n893), .A2(new_n897), .ZN(G75));
  OAI21_X1  g712(.A(new_n881), .B1(new_n887), .B2(KEYINPUT53), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(G210), .A3(G902), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n543), .A2(new_n545), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n546), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT120), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n900), .B2(new_n901), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n247), .A2(G952), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT121), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n610), .B(KEYINPUT57), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n850), .A2(new_n851), .A3(new_n858), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n851), .B1(new_n850), .B2(new_n858), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n878), .B1(new_n915), .B2(new_n883), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n882), .B1(new_n916), .B2(new_n881), .ZN(new_n917));
  INV_X1    g731(.A(new_n888), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n724), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n899), .A2(G902), .A3(new_n794), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n920), .B2(new_n921), .ZN(G54));
  NAND2_X1  g736(.A1(new_n899), .A2(G902), .ZN(new_n923));
  NAND2_X1  g737(.A1(KEYINPUT58), .A2(G475), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(new_n628), .ZN(new_n926));
  INV_X1    g740(.A(new_n628), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n923), .A2(new_n927), .A3(new_n924), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n908), .A3(new_n928), .ZN(G60));
  AND2_X1   g743(.A1(new_n635), .A2(new_n637), .ZN(new_n930));
  XNOR2_X1  g744(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n412), .A2(new_n359), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n930), .B1(new_n892), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n930), .A2(new_n933), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n899), .A2(KEYINPUT54), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n888), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n934), .A2(new_n910), .A3(new_n937), .ZN(G63));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n671), .A2(new_n672), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n430), .A2(new_n359), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n899), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n909), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n470), .A2(new_n473), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n899), .B2(new_n944), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n939), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n950));
  INV_X1    g764(.A(new_n944), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n916), .B2(new_n881), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(new_n947), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(KEYINPUT124), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n909), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n955), .B2(new_n956), .ZN(G66));
  OR3_X1    g771(.A1(new_n862), .A2(new_n863), .A3(new_n871), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n247), .ZN(new_n959));
  INV_X1    g773(.A(G224), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n427), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n902), .B1(G898), .B2(new_n247), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT125), .Z(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  AOI21_X1  g779(.A(new_n247), .B1(G227), .B2(G900), .ZN(new_n966));
  INV_X1    g780(.A(new_n809), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n834), .A2(new_n652), .A3(new_n705), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n798), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n849), .A2(new_n717), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n780), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n777), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n801), .A2(new_n967), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n247), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n239), .B(new_n340), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(G900), .B2(new_n974), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n663), .A2(new_n649), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n760), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n694), .A2(new_n981), .A3(new_n766), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n809), .A2(new_n982), .ZN(new_n983));
  OR3_X1    g797(.A1(new_n707), .A2(new_n970), .A3(KEYINPUT62), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT62), .B1(new_n707), .B2(new_n970), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n983), .A2(new_n801), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n976), .B1(new_n986), .B2(new_n247), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n966), .B1(new_n979), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n975), .B2(new_n978), .ZN(new_n989));
  INV_X1    g803(.A(new_n966), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n988), .A2(new_n991), .ZN(G72));
  XNOR2_X1  g806(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n282), .A2(new_n359), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n993), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n986), .B2(new_n958), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n908), .B1(new_n996), .B2(new_n700), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n283), .B1(new_n258), .B2(new_n262), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n995), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n997), .B1(new_n891), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n699), .A2(new_n253), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n995), .B1(new_n973), .B2(new_n958), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(KEYINPUT127), .B(new_n995), .C1(new_n973), .C2(new_n958), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1000), .A2(new_n1006), .ZN(G57));
endmodule


