

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U556 ( .A1(n549), .A2(n530), .ZN(n548) );
  AND2_X2 U557 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U558 ( .A(n839), .B(KEYINPUT32), .ZN(n540) );
  NOR2_X1 U559 ( .A1(n827), .A2(n826), .ZN(n829) );
  NOR2_X1 U560 ( .A1(n807), .A2(n987), .ZN(n796) );
  NOR2_X1 U561 ( .A1(n533), .A2(n531), .ZN(n804) );
  NOR2_X1 U562 ( .A1(n793), .A2(n792), .ZN(n807) );
  NOR2_X1 U563 ( .A1(G1966), .A2(n865), .ZN(n842) );
  NAND2_X1 U564 ( .A1(G8), .A2(n818), .ZN(n865) );
  AND2_X1 U565 ( .A1(n866), .A2(n536), .ZN(n819) );
  AND2_X1 U566 ( .A1(n576), .A2(n575), .ZN(G164) );
  AND2_X2 U567 ( .A1(n555), .A2(G2105), .ZN(n628) );
  NOR2_X1 U568 ( .A1(n854), .A2(n853), .ZN(n855) );
  INV_X1 U569 ( .A(n1002), .ZN(n853) );
  INV_X1 U570 ( .A(n991), .ZN(n539) );
  NAND2_X1 U571 ( .A1(n548), .A2(n526), .ZN(n544) );
  INV_X1 U572 ( .A(KEYINPUT19), .ZN(n703) );
  NAND2_X1 U573 ( .A1(n535), .A2(n534), .ZN(n533) );
  NAND2_X1 U574 ( .A1(n818), .A2(G1341), .ZN(n535) );
  NAND2_X1 U575 ( .A1(n528), .A2(n539), .ZN(n538) );
  NAND2_X1 U576 ( .A1(n550), .A2(KEYINPUT98), .ZN(n549) );
  NOR2_X1 U577 ( .A1(G164), .A2(G1384), .ZN(n866) );
  INV_X1 U578 ( .A(G2105), .ZN(n543) );
  NAND2_X1 U579 ( .A1(n527), .A2(n523), .ZN(n546) );
  XNOR2_X1 U580 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U581 ( .A(n704), .B(n703), .ZN(n705) );
  NOR2_X1 U582 ( .A1(G651), .A2(n660), .ZN(n735) );
  AND2_X1 U583 ( .A1(n846), .A2(n528), .ZN(n521) );
  NOR2_X1 U584 ( .A1(n872), .A2(n529), .ZN(n522) );
  AND2_X1 U585 ( .A1(n522), .A2(KEYINPUT98), .ZN(n523) );
  AND2_X1 U586 ( .A1(n544), .A2(n522), .ZN(n524) );
  XOR2_X1 U587 ( .A(n849), .B(KEYINPUT64), .Z(n525) );
  INV_X1 U588 ( .A(n819), .ZN(n818) );
  NAND2_X1 U589 ( .A1(n861), .A2(n551), .ZN(n526) );
  AND2_X1 U590 ( .A1(n856), .A2(n855), .ZN(n527) );
  NOR2_X2 U591 ( .A1(G2105), .A2(n555), .ZN(n570) );
  NOR2_X1 U592 ( .A1(n848), .A2(n865), .ZN(n528) );
  AND2_X1 U593 ( .A1(n887), .A2(n936), .ZN(n529) );
  OR2_X1 U594 ( .A1(n865), .A2(n864), .ZN(n530) );
  INV_X1 U595 ( .A(KEYINPUT98), .ZN(n551) );
  XNOR2_X1 U596 ( .A(n532), .B(KEYINPUT26), .ZN(n531) );
  NOR2_X1 U597 ( .A1(n818), .A2(n797), .ZN(n532) );
  INV_X1 U598 ( .A(n985), .ZN(n534) );
  INV_X1 U599 ( .A(n867), .ZN(n536) );
  NAND2_X1 U600 ( .A1(n540), .A2(n521), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n537), .A2(n538), .ZN(n849) );
  NAND2_X1 U602 ( .A1(n540), .A2(n846), .ZN(n859) );
  NAND2_X1 U603 ( .A1(n571), .A2(n541), .ZN(n572) );
  NAND2_X1 U604 ( .A1(n633), .A2(G138), .ZN(n541) );
  XNOR2_X2 U605 ( .A(n542), .B(KEYINPUT17), .ZN(n633) );
  NAND2_X1 U606 ( .A1(n543), .A2(n555), .ZN(n542) );
  NAND2_X1 U607 ( .A1(n545), .A2(n524), .ZN(n547) );
  NAND2_X1 U608 ( .A1(n527), .A2(n548), .ZN(n545) );
  INV_X1 U609 ( .A(n861), .ZN(n550) );
  NAND2_X1 U610 ( .A1(n547), .A2(n546), .ZN(n873) );
  NOR2_X2 U611 ( .A1(n569), .A2(n568), .ZN(G160) );
  AND2_X1 U612 ( .A1(n629), .A2(G114), .ZN(n552) );
  XNOR2_X1 U613 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n823) );
  XNOR2_X1 U614 ( .A(n824), .B(n823), .ZN(n825) );
  INV_X1 U615 ( .A(KEYINPUT29), .ZN(n812) );
  INV_X1 U616 ( .A(KEYINPUT31), .ZN(n828) );
  NOR2_X1 U617 ( .A1(G395), .A2(G397), .ZN(n776) );
  XNOR2_X1 U618 ( .A(G286), .B(n534), .ZN(n738) );
  INV_X1 U619 ( .A(G2104), .ZN(n555) );
  NAND2_X1 U620 ( .A1(G124), .A2(n628), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n553), .B(KEYINPUT44), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(KEYINPUT104), .ZN(n557) );
  NAND2_X1 U623 ( .A1(G100), .A2(n570), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U625 ( .A1(G136), .A2(n633), .ZN(n559) );
  AND2_X1 U626 ( .A1(G2105), .A2(G2104), .ZN(n629) );
  NAND2_X1 U627 ( .A1(G112), .A2(n629), .ZN(n558) );
  NAND2_X1 U628 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U629 ( .A1(n561), .A2(n560), .ZN(G162) );
  NAND2_X1 U630 ( .A1(G101), .A2(n570), .ZN(n562) );
  XOR2_X1 U631 ( .A(KEYINPUT23), .B(n562), .Z(n565) );
  NAND2_X1 U632 ( .A1(G125), .A2(n628), .ZN(n563) );
  XOR2_X1 U633 ( .A(KEYINPUT65), .B(n563), .Z(n564) );
  NAND2_X1 U634 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G137), .A2(n633), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G113), .A2(n629), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U638 ( .A1(G102), .A2(n570), .ZN(n571) );
  XOR2_X1 U639 ( .A(n572), .B(KEYINPUT82), .Z(n576) );
  NAND2_X1 U640 ( .A1(G126), .A2(n628), .ZN(n573) );
  XNOR2_X1 U641 ( .A(KEYINPUT81), .B(n573), .ZN(n574) );
  NOR2_X1 U642 ( .A1(n552), .A2(n574), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G105), .A2(n570), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n577), .B(KEYINPUT38), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G141), .A2(n633), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G117), .A2(n629), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U648 ( .A1(G129), .A2(n628), .ZN(n580) );
  XNOR2_X1 U649 ( .A(KEYINPUT87), .B(n580), .ZN(n581) );
  NOR2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n875) );
  NAND2_X1 U652 ( .A1(G123), .A2(n628), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n585), .B(KEYINPUT18), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G99), .A2(n570), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT73), .B(n586), .Z(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G135), .A2(n633), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G111), .A2(n629), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U660 ( .A1(n592), .A2(n591), .ZN(n937) );
  XOR2_X1 U661 ( .A(G162), .B(n937), .Z(n593) );
  XNOR2_X1 U662 ( .A(n875), .B(n593), .ZN(n606) );
  XOR2_X1 U663 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n595) );
  XNOR2_X1 U664 ( .A(KEYINPUT48), .B(KEYINPUT111), .ZN(n594) );
  XNOR2_X1 U665 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U666 ( .A(KEYINPUT107), .B(n596), .ZN(n604) );
  NAND2_X1 U667 ( .A1(G95), .A2(n570), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G119), .A2(n628), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U670 ( .A1(G131), .A2(n633), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G107), .A2(n629), .ZN(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  OR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n876) );
  XNOR2_X1 U674 ( .A(n876), .B(KEYINPUT106), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n604), .B(n603), .ZN(n605) );
  XOR2_X1 U676 ( .A(n606), .B(n605), .Z(n617) );
  XNOR2_X1 U677 ( .A(KEYINPUT47), .B(KEYINPUT109), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G127), .A2(n628), .ZN(n608) );
  NAND2_X1 U679 ( .A1(G115), .A2(n629), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n610), .B(n609), .ZN(n615) );
  NAND2_X1 U682 ( .A1(n570), .A2(G103), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n611), .B(KEYINPUT108), .ZN(n613) );
  NAND2_X1 U684 ( .A1(G139), .A2(n633), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n942) );
  XNOR2_X1 U687 ( .A(G160), .B(n942), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n617), .B(n616), .ZN(n627) );
  NAND2_X1 U689 ( .A1(G130), .A2(n628), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G118), .A2(n629), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n625) );
  NAND2_X1 U692 ( .A1(n570), .A2(G106), .ZN(n620) );
  XOR2_X1 U693 ( .A(KEYINPUT105), .B(n620), .Z(n622) );
  NAND2_X1 U694 ( .A1(n633), .A2(G142), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U696 ( .A(KEYINPUT45), .B(n623), .Z(n624) );
  NOR2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U698 ( .A(n627), .B(n626), .Z(n643) );
  XNOR2_X1 U699 ( .A(KEYINPUT86), .B(KEYINPUT36), .ZN(n641) );
  NAND2_X1 U700 ( .A1(G128), .A2(n628), .ZN(n631) );
  NAND2_X1 U701 ( .A1(G116), .A2(n629), .ZN(n630) );
  NAND2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U703 ( .A(n632), .B(KEYINPUT35), .ZN(n639) );
  XNOR2_X1 U704 ( .A(KEYINPUT85), .B(KEYINPUT34), .ZN(n637) );
  NAND2_X1 U705 ( .A1(G104), .A2(n570), .ZN(n635) );
  NAND2_X1 U706 ( .A1(G140), .A2(n633), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n638) );
  NAND2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U710 ( .A(n641), .B(n640), .Z(n884) );
  XNOR2_X1 U711 ( .A(G164), .B(n884), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n643), .B(n642), .ZN(n644) );
  NOR2_X1 U713 ( .A1(G37), .A2(n644), .ZN(G395) );
  INV_X1 U714 ( .A(G651), .ZN(n649) );
  NOR2_X1 U715 ( .A1(G543), .A2(n649), .ZN(n645) );
  XOR2_X1 U716 ( .A(KEYINPUT1), .B(n645), .Z(n724) );
  NAND2_X1 U717 ( .A1(G61), .A2(n724), .ZN(n647) );
  NOR2_X1 U718 ( .A1(G651), .A2(G543), .ZN(n726) );
  NAND2_X1 U719 ( .A1(G86), .A2(n726), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n653) );
  XOR2_X1 U721 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  XNOR2_X1 U722 ( .A(KEYINPUT66), .B(n648), .ZN(n660) );
  NOR2_X2 U723 ( .A1(n649), .A2(n660), .ZN(n728) );
  NAND2_X1 U724 ( .A1(G73), .A2(n728), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(KEYINPUT2), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n651), .B(KEYINPUT77), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n735), .A2(G48), .ZN(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G49), .A2(n735), .ZN(n657) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U733 ( .A(KEYINPUT76), .B(n658), .ZN(n659) );
  NOR2_X1 U734 ( .A1(n724), .A2(n659), .ZN(n662) );
  NAND2_X1 U735 ( .A1(G87), .A2(n660), .ZN(n661) );
  NAND2_X1 U736 ( .A1(n662), .A2(n661), .ZN(G288) );
  NAND2_X1 U737 ( .A1(n724), .A2(G62), .ZN(n663) );
  XNOR2_X1 U738 ( .A(n663), .B(KEYINPUT78), .ZN(n665) );
  NAND2_X1 U739 ( .A1(G88), .A2(n726), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n665), .A2(n664), .ZN(n669) );
  NAND2_X1 U741 ( .A1(G75), .A2(n728), .ZN(n667) );
  NAND2_X1 U742 ( .A1(G50), .A2(n735), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U744 ( .A1(n669), .A2(n668), .ZN(G166) );
  INV_X1 U745 ( .A(G166), .ZN(G303) );
  AND2_X1 U746 ( .A1(n724), .A2(G60), .ZN(n673) );
  NAND2_X1 U747 ( .A1(G85), .A2(n726), .ZN(n671) );
  NAND2_X1 U748 ( .A1(G72), .A2(n728), .ZN(n670) );
  NAND2_X1 U749 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U750 ( .A1(n673), .A2(n672), .ZN(n675) );
  NAND2_X1 U751 ( .A1(n735), .A2(G47), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n675), .A2(n674), .ZN(G290) );
  NAND2_X1 U753 ( .A1(G64), .A2(n724), .ZN(n677) );
  NAND2_X1 U754 ( .A1(G52), .A2(n735), .ZN(n676) );
  NAND2_X1 U755 ( .A1(n677), .A2(n676), .ZN(n684) );
  XNOR2_X1 U756 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n728), .A2(G77), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n726), .A2(G90), .ZN(n678) );
  XOR2_X1 U759 ( .A(KEYINPUT67), .B(n678), .Z(n679) );
  NAND2_X1 U760 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U761 ( .A(n682), .B(n681), .Z(n683) );
  NOR2_X1 U762 ( .A1(n684), .A2(n683), .ZN(G171) );
  INV_X1 U763 ( .A(G171), .ZN(G301) );
  NAND2_X1 U764 ( .A1(n726), .A2(G89), .ZN(n685) );
  XNOR2_X1 U765 ( .A(n685), .B(KEYINPUT4), .ZN(n687) );
  NAND2_X1 U766 ( .A1(G76), .A2(n728), .ZN(n686) );
  NAND2_X1 U767 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U768 ( .A(n688), .B(KEYINPUT5), .ZN(n693) );
  NAND2_X1 U769 ( .A1(G63), .A2(n724), .ZN(n690) );
  NAND2_X1 U770 ( .A1(G51), .A2(n735), .ZN(n689) );
  NAND2_X1 U771 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U772 ( .A(KEYINPUT6), .B(n691), .Z(n692) );
  NAND2_X1 U773 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U774 ( .A(n694), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U775 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U776 ( .A1(G67), .A2(n724), .ZN(n696) );
  NAND2_X1 U777 ( .A1(G93), .A2(n726), .ZN(n695) );
  NAND2_X1 U778 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U779 ( .A1(G80), .A2(n728), .ZN(n697) );
  XNOR2_X1 U780 ( .A(KEYINPUT75), .B(n697), .ZN(n698) );
  NOR2_X1 U781 ( .A1(n699), .A2(n698), .ZN(n701) );
  NAND2_X1 U782 ( .A1(n735), .A2(G55), .ZN(n700) );
  NAND2_X1 U783 ( .A1(n701), .A2(n700), .ZN(n915) );
  XOR2_X1 U784 ( .A(G305), .B(G288), .Z(n702) );
  XNOR2_X1 U785 ( .A(n915), .B(n702), .ZN(n706) );
  XOR2_X1 U786 ( .A(G303), .B(KEYINPUT79), .Z(n704) );
  XNOR2_X1 U787 ( .A(n707), .B(G290), .ZN(n714) );
  NAND2_X1 U788 ( .A1(G65), .A2(n724), .ZN(n709) );
  NAND2_X1 U789 ( .A1(G53), .A2(n735), .ZN(n708) );
  NAND2_X1 U790 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U791 ( .A1(G91), .A2(n726), .ZN(n711) );
  NAND2_X1 U792 ( .A1(G78), .A2(n728), .ZN(n710) );
  NAND2_X1 U793 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U794 ( .A1(n713), .A2(n712), .ZN(n987) );
  XOR2_X1 U795 ( .A(n714), .B(n987), .Z(n912) );
  XOR2_X1 U796 ( .A(KEYINPUT112), .B(n912), .Z(n723) );
  NAND2_X1 U797 ( .A1(G66), .A2(n724), .ZN(n716) );
  NAND2_X1 U798 ( .A1(G92), .A2(n726), .ZN(n715) );
  NAND2_X1 U799 ( .A1(n716), .A2(n715), .ZN(n720) );
  NAND2_X1 U800 ( .A1(G79), .A2(n728), .ZN(n718) );
  NAND2_X1 U801 ( .A1(G54), .A2(n735), .ZN(n717) );
  NAND2_X1 U802 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U803 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U804 ( .A(KEYINPUT15), .B(n721), .Z(n982) );
  XOR2_X1 U805 ( .A(G301), .B(n982), .Z(n722) );
  XNOR2_X1 U806 ( .A(n723), .B(n722), .ZN(n739) );
  NAND2_X1 U807 ( .A1(n724), .A2(G56), .ZN(n725) );
  XNOR2_X1 U808 ( .A(KEYINPUT14), .B(n725), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n726), .A2(G81), .ZN(n727) );
  XNOR2_X1 U810 ( .A(n727), .B(KEYINPUT12), .ZN(n730) );
  NAND2_X1 U811 ( .A1(G68), .A2(n728), .ZN(n729) );
  NAND2_X1 U812 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U813 ( .A(KEYINPUT13), .B(n731), .ZN(n732) );
  NAND2_X1 U814 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U815 ( .A(n734), .B(KEYINPUT69), .ZN(n737) );
  NAND2_X1 U816 ( .A1(n735), .A2(G43), .ZN(n736) );
  NAND2_X1 U817 ( .A1(n737), .A2(n736), .ZN(n985) );
  XNOR2_X1 U818 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U819 ( .A1(G37), .A2(n740), .ZN(G397) );
  XOR2_X1 U820 ( .A(G2443), .B(G2446), .Z(n742) );
  XNOR2_X1 U821 ( .A(G2427), .B(G2451), .ZN(n741) );
  XNOR2_X1 U822 ( .A(n742), .B(n741), .ZN(n748) );
  XOR2_X1 U823 ( .A(G2430), .B(G2454), .Z(n744) );
  XNOR2_X1 U824 ( .A(G1341), .B(G1348), .ZN(n743) );
  XNOR2_X1 U825 ( .A(n744), .B(n743), .ZN(n746) );
  XOR2_X1 U826 ( .A(G2435), .B(G2438), .Z(n745) );
  XNOR2_X1 U827 ( .A(n746), .B(n745), .ZN(n747) );
  XOR2_X1 U828 ( .A(n748), .B(n747), .Z(n749) );
  AND2_X1 U829 ( .A1(G14), .A2(n749), .ZN(G401) );
  XNOR2_X1 U830 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U831 ( .A(G82), .ZN(G220) );
  INV_X1 U832 ( .A(G132), .ZN(G219) );
  INV_X1 U833 ( .A(G57), .ZN(G237) );
  NOR2_X1 U834 ( .A1(G220), .A2(G219), .ZN(n750) );
  XOR2_X1 U835 ( .A(KEYINPUT22), .B(n750), .Z(n751) );
  NOR2_X1 U836 ( .A1(G218), .A2(n751), .ZN(n752) );
  NAND2_X1 U837 ( .A1(G96), .A2(n752), .ZN(n1043) );
  NAND2_X1 U838 ( .A1(n1043), .A2(G2106), .ZN(n756) );
  NAND2_X1 U839 ( .A1(G69), .A2(G120), .ZN(n753) );
  NOR2_X1 U840 ( .A1(G237), .A2(n753), .ZN(n754) );
  NAND2_X1 U841 ( .A1(G108), .A2(n754), .ZN(n1044) );
  NAND2_X1 U842 ( .A1(n1044), .A2(G567), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n925) );
  INV_X1 U844 ( .A(n925), .ZN(G319) );
  XOR2_X1 U845 ( .A(KEYINPUT102), .B(G2678), .Z(n758) );
  XNOR2_X1 U846 ( .A(G2090), .B(G2072), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n758), .B(n757), .ZN(n762) );
  XOR2_X1 U848 ( .A(KEYINPUT43), .B(KEYINPUT103), .Z(n760) );
  XNOR2_X1 U849 ( .A(G2067), .B(KEYINPUT42), .ZN(n759) );
  XNOR2_X1 U850 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U851 ( .A(n762), .B(n761), .Z(n764) );
  INV_X1 U852 ( .A(G2100), .ZN(n907) );
  XOR2_X1 U853 ( .A(G2096), .B(n907), .Z(n763) );
  XNOR2_X1 U854 ( .A(n764), .B(n763), .ZN(n766) );
  XOR2_X1 U855 ( .A(G2078), .B(G2084), .Z(n765) );
  XNOR2_X1 U856 ( .A(n766), .B(n765), .ZN(G227) );
  INV_X1 U857 ( .A(G1971), .ZN(n1023) );
  XNOR2_X1 U858 ( .A(n1023), .B(G1956), .ZN(n768) );
  XNOR2_X1 U859 ( .A(G1986), .B(G1961), .ZN(n767) );
  XNOR2_X1 U860 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U861 ( .A(n769), .B(G2474), .Z(n771) );
  XNOR2_X1 U862 ( .A(G1966), .B(G1976), .ZN(n770) );
  XNOR2_X1 U863 ( .A(n771), .B(n770), .ZN(n775) );
  XOR2_X1 U864 ( .A(KEYINPUT41), .B(G1981), .Z(n773) );
  INV_X1 U865 ( .A(G1996), .ZN(n797) );
  XOR2_X1 U866 ( .A(n797), .B(G1991), .Z(n772) );
  XNOR2_X1 U867 ( .A(n773), .B(n772), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n775), .B(n774), .ZN(G229) );
  XNOR2_X1 U869 ( .A(KEYINPUT114), .B(n776), .ZN(n782) );
  NOR2_X1 U870 ( .A1(G227), .A2(G229), .ZN(n777) );
  XOR2_X1 U871 ( .A(KEYINPUT49), .B(n777), .Z(n778) );
  NAND2_X1 U872 ( .A1(G319), .A2(n778), .ZN(n779) );
  NOR2_X1 U873 ( .A1(G401), .A2(n779), .ZN(n780) );
  XOR2_X1 U874 ( .A(KEYINPUT113), .B(n780), .Z(n781) );
  NAND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(G225) );
  XNOR2_X1 U876 ( .A(G225), .B(KEYINPUT115), .ZN(G308) );
  XOR2_X1 U877 ( .A(G2078), .B(KEYINPUT25), .Z(n783) );
  XNOR2_X1 U878 ( .A(KEYINPUT92), .B(n783), .ZN(n961) );
  NAND2_X1 U879 ( .A1(G40), .A2(G160), .ZN(n785) );
  INV_X1 U880 ( .A(KEYINPUT83), .ZN(n784) );
  XNOR2_X1 U881 ( .A(n785), .B(n784), .ZN(n867) );
  INV_X1 U882 ( .A(KEYINPUT91), .ZN(n786) );
  XNOR2_X1 U883 ( .A(n819), .B(n786), .ZN(n789) );
  INV_X1 U884 ( .A(n789), .ZN(n799) );
  NOR2_X1 U885 ( .A1(n961), .A2(n799), .ZN(n788) );
  INV_X1 U886 ( .A(n818), .ZN(n798) );
  NOR2_X1 U887 ( .A1(n798), .A2(G1961), .ZN(n787) );
  NOR2_X1 U888 ( .A1(n788), .A2(n787), .ZN(n816) );
  OR2_X1 U889 ( .A1(n816), .A2(G301), .ZN(n815) );
  XOR2_X1 U890 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n791) );
  NAND2_X1 U891 ( .A1(G2072), .A2(n789), .ZN(n790) );
  XNOR2_X1 U892 ( .A(n791), .B(n790), .ZN(n793) );
  AND2_X1 U893 ( .A1(n799), .A2(G1956), .ZN(n792) );
  XNOR2_X1 U894 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n794) );
  XNOR2_X1 U895 ( .A(n794), .B(KEYINPUT28), .ZN(n795) );
  XNOR2_X1 U896 ( .A(n796), .B(n795), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n982), .A2(n804), .ZN(n803) );
  NAND2_X1 U898 ( .A1(G2067), .A2(n789), .ZN(n801) );
  NAND2_X1 U899 ( .A1(G1348), .A2(n818), .ZN(n800) );
  NAND2_X1 U900 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U901 ( .A1(n803), .A2(n802), .ZN(n806) );
  OR2_X1 U902 ( .A1(n982), .A2(n804), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n807), .A2(n987), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n813), .B(n812), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n831) );
  NAND2_X1 U909 ( .A1(n816), .A2(G301), .ZN(n817) );
  XNOR2_X1 U910 ( .A(n817), .B(KEYINPUT97), .ZN(n827) );
  INV_X1 U911 ( .A(G2084), .ZN(n820) );
  AND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U913 ( .A(n821), .B(KEYINPUT90), .ZN(n840) );
  NOR2_X1 U914 ( .A1(n842), .A2(n840), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n822), .A2(G8), .ZN(n824) );
  NOR2_X1 U916 ( .A1(n825), .A2(G168), .ZN(n826) );
  XNOR2_X1 U917 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U918 ( .A1(n831), .A2(n830), .ZN(n841) );
  NAND2_X1 U919 ( .A1(n841), .A2(G286), .ZN(n838) );
  INV_X1 U920 ( .A(G8), .ZN(n836) );
  NOR2_X1 U921 ( .A1(G1971), .A2(n865), .ZN(n833) );
  NOR2_X1 U922 ( .A1(G2090), .A2(n818), .ZN(n832) );
  NOR2_X1 U923 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U924 ( .A1(n834), .A2(G303), .ZN(n835) );
  OR2_X1 U925 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U926 ( .A1(n840), .A2(G8), .ZN(n845) );
  INV_X1 U927 ( .A(n841), .ZN(n843) );
  NOR2_X1 U928 ( .A1(n843), .A2(n842), .ZN(n844) );
  NAND2_X1 U929 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U930 ( .A1(G1976), .A2(G288), .ZN(n851) );
  NOR2_X1 U931 ( .A1(G1971), .A2(G303), .ZN(n847) );
  NOR2_X1 U932 ( .A1(n851), .A2(n847), .ZN(n991) );
  NAND2_X1 U933 ( .A1(G1976), .A2(G288), .ZN(n995) );
  INV_X1 U934 ( .A(n995), .ZN(n848) );
  INV_X1 U935 ( .A(KEYINPUT33), .ZN(n850) );
  NAND2_X1 U936 ( .A1(n525), .A2(n850), .ZN(n856) );
  NAND2_X1 U937 ( .A1(n851), .A2(KEYINPUT33), .ZN(n852) );
  NOR2_X1 U938 ( .A1(n852), .A2(n865), .ZN(n854) );
  XOR2_X1 U939 ( .A(G1981), .B(G305), .Z(n1002) );
  NOR2_X1 U940 ( .A1(G2090), .A2(G303), .ZN(n857) );
  NAND2_X1 U941 ( .A1(G8), .A2(n857), .ZN(n858) );
  NAND2_X1 U942 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U943 ( .A1(n860), .A2(n865), .ZN(n861) );
  NOR2_X1 U944 ( .A1(G1981), .A2(G305), .ZN(n862) );
  XNOR2_X1 U945 ( .A(n862), .B(KEYINPUT89), .ZN(n863) );
  XNOR2_X1 U946 ( .A(n863), .B(KEYINPUT24), .ZN(n864) );
  NOR2_X1 U947 ( .A1(n867), .A2(n866), .ZN(n887) );
  XNOR2_X1 U948 ( .A(G1986), .B(G290), .ZN(n993) );
  NAND2_X1 U949 ( .A1(n887), .A2(n993), .ZN(n868) );
  XOR2_X1 U950 ( .A(KEYINPUT84), .B(n868), .Z(n872) );
  NAND2_X1 U951 ( .A1(n875), .A2(G1996), .ZN(n870) );
  NAND2_X1 U952 ( .A1(G1991), .A2(n876), .ZN(n869) );
  NAND2_X1 U953 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U954 ( .A(n871), .B(KEYINPUT88), .ZN(n936) );
  XNOR2_X1 U955 ( .A(G2067), .B(KEYINPUT37), .ZN(n883) );
  NOR2_X1 U956 ( .A1(n883), .A2(n884), .ZN(n932) );
  NAND2_X1 U957 ( .A1(n887), .A2(n932), .ZN(n881) );
  AND2_X1 U958 ( .A1(n873), .A2(n881), .ZN(n874) );
  XNOR2_X1 U959 ( .A(n874), .B(KEYINPUT99), .ZN(n889) );
  NOR2_X1 U960 ( .A1(G1996), .A2(n875), .ZN(n947) );
  NOR2_X1 U961 ( .A1(G1991), .A2(n876), .ZN(n938) );
  NOR2_X1 U962 ( .A1(G1986), .A2(G290), .ZN(n877) );
  NOR2_X1 U963 ( .A1(n938), .A2(n877), .ZN(n878) );
  NOR2_X1 U964 ( .A1(n529), .A2(n878), .ZN(n879) );
  NOR2_X1 U965 ( .A1(n947), .A2(n879), .ZN(n880) );
  XNOR2_X1 U966 ( .A(n880), .B(KEYINPUT39), .ZN(n882) );
  NAND2_X1 U967 ( .A1(n882), .A2(n881), .ZN(n885) );
  NAND2_X1 U968 ( .A1(n884), .A2(n883), .ZN(n952) );
  NAND2_X1 U969 ( .A1(n885), .A2(n952), .ZN(n886) );
  NAND2_X1 U970 ( .A1(n887), .A2(n886), .ZN(n888) );
  NAND2_X1 U971 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U972 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n890) );
  XNOR2_X1 U973 ( .A(n891), .B(n890), .ZN(G329) );
  AND2_X1 U974 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U975 ( .A1(G7), .A2(G661), .ZN(n892) );
  XOR2_X1 U976 ( .A(n892), .B(KEYINPUT10), .Z(n926) );
  NAND2_X1 U977 ( .A1(n926), .A2(G567), .ZN(n893) );
  XOR2_X1 U978 ( .A(KEYINPUT11), .B(n893), .Z(G234) );
  INV_X1 U979 ( .A(G860), .ZN(n899) );
  OR2_X1 U980 ( .A1(n985), .A2(n899), .ZN(G153) );
  OR2_X1 U981 ( .A1(n982), .A2(G868), .ZN(n894) );
  XNOR2_X1 U982 ( .A(n894), .B(KEYINPUT70), .ZN(n896) );
  NAND2_X1 U983 ( .A1(G868), .A2(G301), .ZN(n895) );
  NAND2_X1 U984 ( .A1(n896), .A2(n895), .ZN(G284) );
  INV_X1 U985 ( .A(n987), .ZN(G299) );
  INV_X1 U986 ( .A(G868), .ZN(n916) );
  NOR2_X1 U987 ( .A1(G286), .A2(n916), .ZN(n898) );
  NOR2_X1 U988 ( .A1(G868), .A2(G299), .ZN(n897) );
  NOR2_X1 U989 ( .A1(n898), .A2(n897), .ZN(G297) );
  NAND2_X1 U990 ( .A1(n899), .A2(G559), .ZN(n900) );
  NAND2_X1 U991 ( .A1(n900), .A2(n982), .ZN(n901) );
  XNOR2_X1 U992 ( .A(n901), .B(KEYINPUT16), .ZN(n902) );
  XOR2_X1 U993 ( .A(KEYINPUT71), .B(n902), .Z(G148) );
  NOR2_X1 U994 ( .A1(G868), .A2(n985), .ZN(n903) );
  XNOR2_X1 U995 ( .A(KEYINPUT72), .B(n903), .ZN(n906) );
  NAND2_X1 U996 ( .A1(G868), .A2(n982), .ZN(n904) );
  NOR2_X1 U997 ( .A1(G559), .A2(n904), .ZN(n905) );
  NOR2_X1 U998 ( .A1(n906), .A2(n905), .ZN(G282) );
  XNOR2_X1 U999 ( .A(n937), .B(G2096), .ZN(n908) );
  NAND2_X1 U1000 ( .A1(n908), .A2(n907), .ZN(G156) );
  NAND2_X1 U1001 ( .A1(G559), .A2(n982), .ZN(n909) );
  XNOR2_X1 U1002 ( .A(n985), .B(n909), .ZN(n913) );
  NOR2_X1 U1003 ( .A1(n913), .A2(G860), .ZN(n911) );
  XOR2_X1 U1004 ( .A(n915), .B(KEYINPUT74), .Z(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(G145) );
  XOR2_X1 U1006 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1007 ( .A1(n914), .A2(G868), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1009 ( .A1(n918), .A2(n917), .ZN(G295) );
  NAND2_X1 U1010 ( .A1(G2078), .A2(G2084), .ZN(n919) );
  XOR2_X1 U1011 ( .A(KEYINPUT20), .B(n919), .Z(n920) );
  NAND2_X1 U1012 ( .A1(G2090), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1013 ( .A(KEYINPUT80), .B(KEYINPUT21), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(n922), .B(n921), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(G2072), .A2(n923), .ZN(G158) );
  NAND2_X1 U1016 ( .A1(G483), .A2(G661), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(n925), .A2(n924), .ZN(n931) );
  NAND2_X1 U1018 ( .A1(n931), .A2(G36), .ZN(G176) );
  NAND2_X1 U1019 ( .A1(G2106), .A2(n926), .ZN(G217) );
  INV_X1 U1020 ( .A(n926), .ZN(G223) );
  NAND2_X1 U1021 ( .A1(G15), .A2(G2), .ZN(n928) );
  INV_X1 U1022 ( .A(G661), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1024 ( .A(n929), .B(KEYINPUT101), .ZN(G259) );
  NAND2_X1 U1025 ( .A1(G3), .A2(G1), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(G188) );
  XNOR2_X1 U1028 ( .A(G2084), .B(G160), .ZN(n934) );
  INV_X1 U1029 ( .A(n932), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n940) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT116), .B(n941), .ZN(n955) );
  XOR2_X1 U1035 ( .A(G2072), .B(n942), .Z(n944) );
  XOR2_X1 U1036 ( .A(G164), .B(G2078), .Z(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1038 ( .A(KEYINPUT50), .B(n945), .Z(n951) );
  XOR2_X1 U1039 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1041 ( .A(KEYINPUT117), .B(n948), .Z(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT51), .B(n949), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n953) );
  NAND2_X1 U1044 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1045 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n956), .ZN(n958) );
  INV_X1 U1047 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1049 ( .A1(n959), .A2(G29), .ZN(n1041) );
  XNOR2_X1 U1050 ( .A(G2090), .B(G35), .ZN(n974) );
  XOR2_X1 U1051 ( .A(G2072), .B(G33), .Z(n960) );
  NAND2_X1 U1052 ( .A1(n960), .A2(G28), .ZN(n971) );
  XOR2_X1 U1053 ( .A(n961), .B(G27), .Z(n964) );
  XOR2_X1 U1054 ( .A(G32), .B(G1996), .Z(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT118), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(KEYINPUT119), .B(n965), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(G2067), .B(G26), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G1991), .B(G25), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1062 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n972), .ZN(n973) );
  NOR2_X1 U1064 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n975) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n975), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1068 ( .A(KEYINPUT55), .B(n978), .Z(n980) );
  INV_X1 U1069 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n981), .ZN(n1039) );
  INV_X1 U1072 ( .A(G16), .ZN(n1035) );
  XOR2_X1 U1073 ( .A(n1035), .B(KEYINPUT56), .Z(n1008) );
  XNOR2_X1 U1074 ( .A(n982), .B(G1348), .ZN(n984) );
  XOR2_X1 U1075 ( .A(G301), .B(G1961), .Z(n983) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n1000) );
  XNOR2_X1 U1077 ( .A(n985), .B(G1341), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n986), .B(KEYINPUT121), .ZN(n998) );
  XOR2_X1 U1079 ( .A(G1956), .B(n987), .Z(n989) );
  NOR2_X1 U1080 ( .A1(n1023), .A2(G166), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1085 ( .A(KEYINPUT120), .B(n996), .Z(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(n1001), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G1966), .B(G168), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT57), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1037) );
  XNOR2_X1 U1094 ( .A(KEYINPUT123), .B(G1961), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(n1009), .B(G5), .ZN(n1022) );
  XNOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(n1010), .B(G4), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G1341), .B(G19), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1102 ( .A(KEYINPUT124), .B(G1956), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(G20), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1105 ( .A(KEYINPUT60), .B(n1018), .Z(n1020) );
  XNOR2_X1 U1106 ( .A(G1966), .B(G21), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1032) );
  XNOR2_X1 U1109 ( .A(n1023), .B(G22), .ZN(n1024) );
  XNOR2_X1 U1110 ( .A(KEYINPUT125), .B(n1024), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(G23), .B(G1976), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1113 ( .A(KEYINPUT126), .B(n1027), .Z(n1029) );
  XNOR2_X1 U1114 ( .A(G1986), .B(G24), .ZN(n1028) );
  NOR2_X1 U1115 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1116 ( .A(KEYINPUT58), .B(n1030), .Z(n1031) );
  NOR2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1118 ( .A(KEYINPUT61), .B(n1033), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1120 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1121 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1122 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XOR2_X1 U1123 ( .A(KEYINPUT62), .B(n1042), .Z(G311) );
  XNOR2_X1 U1124 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1125 ( .A(G120), .ZN(G236) );
  INV_X1 U1126 ( .A(G96), .ZN(G221) );
  INV_X1 U1127 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1128 ( .A1(n1044), .A2(n1043), .ZN(G325) );
  INV_X1 U1129 ( .A(G325), .ZN(G261) );
  INV_X1 U1130 ( .A(G108), .ZN(G238) );
endmodule

