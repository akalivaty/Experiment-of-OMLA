

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768;

  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n547) );
  AND2_X1 U372 ( .A1(n377), .A2(n353), .ZN(n374) );
  NOR2_X1 U373 ( .A1(n730), .A2(G902), .ZN(n559) );
  OR2_X2 U374 ( .A1(n436), .A2(n432), .ZN(n700) );
  INV_X1 U375 ( .A(G953), .ZN(n760) );
  XNOR2_X1 U376 ( .A(n407), .B(KEYINPUT42), .ZN(n467) );
  XNOR2_X1 U377 ( .A(n402), .B(KEYINPUT35), .ZN(n765) );
  XOR2_X1 U378 ( .A(n575), .B(n574), .Z(n349) );
  XNOR2_X1 U379 ( .A(n618), .B(KEYINPUT38), .ZN(n710) );
  XNOR2_X2 U380 ( .A(n700), .B(n357), .ZN(n626) );
  XNOR2_X2 U381 ( .A(G116), .B(G119), .ZN(n505) );
  XNOR2_X2 U382 ( .A(n637), .B(KEYINPUT112), .ZN(n714) );
  XNOR2_X2 U383 ( .A(n409), .B(n502), .ZN(n553) );
  NOR2_X2 U384 ( .A1(n694), .A2(n693), .ZN(n594) );
  NOR2_X1 U385 ( .A1(n590), .A2(n589), .ZN(n679) );
  XNOR2_X1 U386 ( .A(n487), .B(n485), .ZN(n723) );
  NOR2_X1 U387 ( .A1(n638), .A2(n478), .ZN(n477) );
  OR2_X1 U388 ( .A1(n464), .A2(n404), .ZN(n638) );
  XNOR2_X1 U389 ( .A(n629), .B(n465), .ZN(n613) );
  AND2_X1 U390 ( .A1(n450), .A2(n448), .ZN(n447) );
  BUF_X1 U391 ( .A(n686), .Z(n758) );
  XNOR2_X1 U392 ( .A(n650), .B(KEYINPUT82), .ZN(n686) );
  NAND2_X1 U393 ( .A1(n351), .A2(n401), .ZN(n764) );
  NAND2_X1 U394 ( .A1(n588), .A2(n696), .ZN(n662) );
  XNOR2_X1 U395 ( .A(n587), .B(KEYINPUT85), .ZN(n588) );
  AND2_X1 U396 ( .A1(n426), .A2(n630), .ZN(n500) );
  XNOR2_X1 U397 ( .A(n494), .B(n493), .ZN(n767) );
  NAND2_X1 U398 ( .A1(n408), .A2(n477), .ZN(n407) );
  XNOR2_X1 U399 ( .A(n460), .B(n468), .ZN(n675) );
  AND2_X1 U400 ( .A1(n479), .A2(n482), .ZN(n408) );
  NOR2_X1 U401 ( .A1(n638), .A2(n613), .ZN(n460) );
  NOR2_X1 U402 ( .A1(n595), .A2(n498), .ZN(n497) );
  INV_X1 U403 ( .A(n609), .ZN(n696) );
  XNOR2_X1 U404 ( .A(n576), .B(n349), .ZN(n609) );
  XNOR2_X1 U405 ( .A(n496), .B(n741), .ZN(n659) );
  XNOR2_X1 U406 ( .A(n505), .B(n504), .ZN(n506) );
  NOR2_X2 U407 ( .A1(n375), .A2(n374), .ZN(n650) );
  NAND2_X1 U408 ( .A1(n645), .A2(n709), .ZN(n629) );
  XNOR2_X1 U409 ( .A(G134), .B(G131), .ZN(n502) );
  AND2_X1 U410 ( .A1(n675), .A2(n419), .ZN(n616) );
  XOR2_X1 U411 ( .A(G902), .B(KEYINPUT15), .Z(n653) );
  AND2_X1 U412 ( .A1(n597), .A2(n662), .ZN(n393) );
  NOR2_X1 U413 ( .A1(n758), .A2(KEYINPUT2), .ZN(n687) );
  INV_X1 U414 ( .A(KEYINPUT0), .ZN(n499) );
  NAND2_X1 U415 ( .A1(n438), .A2(n437), .ZN(n436) );
  NAND2_X1 U416 ( .A1(n435), .A2(n434), .ZN(n433) );
  XNOR2_X1 U417 ( .A(n540), .B(n539), .ZN(n590) );
  XNOR2_X1 U418 ( .A(n639), .B(KEYINPUT46), .ZN(n424) );
  NOR2_X1 U419 ( .A1(n500), .A2(n633), .ZN(n634) );
  AND2_X1 U420 ( .A1(n443), .A2(n475), .ZN(n442) );
  NAND2_X1 U421 ( .A1(n764), .A2(n671), .ZN(n400) );
  NAND2_X1 U422 ( .A1(n710), .A2(n709), .ZN(n637) );
  NOR2_X1 U423 ( .A1(n663), .A2(n628), .ZN(n641) );
  XNOR2_X1 U424 ( .A(n486), .B(KEYINPUT87), .ZN(n485) );
  INV_X1 U425 ( .A(KEYINPUT33), .ZN(n486) );
  AND2_X1 U426 ( .A1(n709), .A2(n386), .ZN(n383) );
  AND2_X1 U427 ( .A1(n385), .A2(n381), .ZN(n380) );
  OR2_X1 U428 ( .A1(n709), .A2(n386), .ZN(n381) );
  INV_X1 U429 ( .A(n607), .ZN(n385) );
  INV_X1 U430 ( .A(KEYINPUT30), .ZN(n386) );
  OR2_X1 U431 ( .A1(G902), .A2(G237), .ZN(n521) );
  INV_X1 U432 ( .A(n653), .ZN(n517) );
  XNOR2_X1 U433 ( .A(n573), .B(n572), .ZN(n575) );
  XNOR2_X1 U434 ( .A(n363), .B(n545), .ZN(n548) );
  XNOR2_X1 U435 ( .A(n546), .B(n356), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n553), .B(n552), .ZN(n755) );
  XNOR2_X1 U437 ( .A(n565), .B(KEYINPUT93), .ZN(n552) );
  AND2_X1 U438 ( .A1(n654), .A2(n653), .ZN(n472) );
  XNOR2_X1 U439 ( .A(n397), .B(n516), .ZN(n496) );
  XNOR2_X1 U440 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U441 ( .A(n409), .B(n398), .ZN(n397) );
  XNOR2_X1 U442 ( .A(n604), .B(n390), .ZN(n389) );
  INV_X1 U443 ( .A(KEYINPUT39), .ZN(n390) );
  NOR2_X1 U444 ( .A1(n617), .A2(n636), .ZN(n604) );
  INV_X1 U445 ( .A(n710), .ZN(n636) );
  INV_X1 U446 ( .A(KEYINPUT19), .ZN(n465) );
  INV_X1 U447 ( .A(KEYINPUT28), .ZN(n611) );
  NOR2_X1 U448 ( .A1(n625), .A2(n610), .ZN(n612) );
  XNOR2_X1 U449 ( .A(n595), .B(n583), .ZN(n591) );
  XNOR2_X1 U450 ( .A(n553), .B(n490), .ZN(n655) );
  XNOR2_X1 U451 ( .A(n492), .B(n508), .ZN(n491) );
  XOR2_X1 U452 ( .A(KEYINPUT5), .B(G137), .Z(n508) );
  XNOR2_X1 U453 ( .A(n461), .B(n536), .ZN(n736) );
  XNOR2_X1 U454 ( .A(n535), .B(n355), .ZN(n461) );
  XNOR2_X1 U455 ( .A(G116), .B(G122), .ZN(n530) );
  BUF_X1 U456 ( .A(n734), .Z(n737) );
  XNOR2_X1 U457 ( .A(n755), .B(n484), .ZN(n730) );
  XNOR2_X1 U458 ( .A(n557), .B(n558), .ZN(n484) );
  XNOR2_X1 U459 ( .A(n556), .B(G140), .ZN(n557) );
  XNOR2_X1 U460 ( .A(n415), .B(n555), .ZN(n556) );
  NAND2_X1 U461 ( .A1(n734), .A2(G210), .ZN(n471) );
  NOR2_X1 U462 ( .A1(n727), .A2(KEYINPUT123), .ZN(n449) );
  INV_X1 U463 ( .A(KEYINPUT48), .ZN(n378) );
  NAND2_X1 U464 ( .A1(n424), .A2(n378), .ZN(n370) );
  NAND2_X1 U465 ( .A1(n766), .A2(n367), .ZN(n443) );
  NAND2_X1 U466 ( .A1(G234), .A2(G237), .ZN(n522) );
  XNOR2_X1 U467 ( .A(n594), .B(KEYINPUT108), .ZN(n488) );
  XOR2_X1 U468 ( .A(G125), .B(G146), .Z(n541) );
  XOR2_X1 U469 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n538) );
  XNOR2_X1 U470 ( .A(G107), .B(KEYINPUT101), .ZN(n528) );
  XNOR2_X1 U471 ( .A(G113), .B(G122), .ZN(n542) );
  XOR2_X1 U472 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n544) );
  XNOR2_X1 U473 ( .A(G104), .B(G143), .ZN(n543) );
  INV_X1 U474 ( .A(KEYINPUT4), .ZN(n501) );
  XNOR2_X1 U475 ( .A(n399), .B(n405), .ZN(n398) );
  NAND2_X1 U476 ( .A1(n760), .A2(G224), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n474), .B(KEYINPUT90), .ZN(n399) );
  XNOR2_X1 U478 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n474) );
  INV_X1 U479 ( .A(KEYINPUT80), .ZN(n425) );
  AND2_X1 U480 ( .A1(n650), .A2(KEYINPUT2), .ZN(n648) );
  INV_X1 U481 ( .A(KEYINPUT41), .ZN(n483) );
  NAND2_X1 U482 ( .A1(n712), .A2(n483), .ZN(n481) );
  INV_X1 U483 ( .A(G902), .ZN(n434) );
  INV_X1 U484 ( .A(G472), .ZN(n435) );
  NAND2_X1 U485 ( .A1(n655), .A2(G472), .ZN(n438) );
  NAND2_X1 U486 ( .A1(G902), .A2(G472), .ZN(n437) );
  XNOR2_X1 U487 ( .A(n459), .B(n458), .ZN(n492) );
  INV_X1 U488 ( .A(G146), .ZN(n458) );
  XOR2_X1 U489 ( .A(G137), .B(KEYINPUT67), .Z(n565) );
  XNOR2_X1 U490 ( .A(G119), .B(G110), .ZN(n560) );
  XNOR2_X1 U491 ( .A(n541), .B(n418), .ZN(n754) );
  XNOR2_X1 U492 ( .A(G140), .B(KEYINPUT10), .ZN(n418) );
  XNOR2_X1 U493 ( .A(n462), .B(n529), .ZN(n531) );
  XOR2_X1 U494 ( .A(KEYINPUT9), .B(KEYINPUT102), .Z(n529) );
  XNOR2_X1 U495 ( .A(n528), .B(n463), .ZN(n462) );
  INV_X1 U496 ( .A(KEYINPUT7), .ZN(n463) );
  XNOR2_X1 U497 ( .A(n554), .B(n416), .ZN(n415) );
  INV_X1 U498 ( .A(KEYINPUT94), .ZN(n416) );
  XOR2_X1 U499 ( .A(G104), .B(G107), .Z(n512) );
  AND2_X1 U500 ( .A1(n727), .A2(KEYINPUT123), .ZN(n451) );
  INV_X1 U501 ( .A(n481), .ZN(n478) );
  NOR2_X1 U502 ( .A1(n384), .A2(n379), .ZN(n602) );
  NAND2_X1 U503 ( .A1(n382), .A2(n380), .ZN(n379) );
  XNOR2_X1 U504 ( .A(n518), .B(KEYINPUT77), .ZN(n519) );
  NOR2_X1 U505 ( .A1(G902), .A2(n739), .ZN(n576) );
  NAND2_X1 U506 ( .A1(n480), .A2(n697), .ZN(n498) );
  INV_X1 U507 ( .A(n700), .ZN(n610) );
  INV_X1 U508 ( .A(KEYINPUT123), .ZN(n445) );
  XNOR2_X1 U509 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U510 ( .A(n428), .B(n427), .ZN(n426) );
  INV_X1 U511 ( .A(KEYINPUT36), .ZN(n427) );
  XNOR2_X1 U512 ( .A(n364), .B(n584), .ZN(n403) );
  XNOR2_X1 U513 ( .A(n396), .B(n395), .ZN(n680) );
  XNOR2_X1 U514 ( .A(KEYINPUT31), .B(KEYINPUT98), .ZN(n395) );
  INV_X1 U515 ( .A(KEYINPUT75), .ZN(n468) );
  XOR2_X1 U516 ( .A(n655), .B(KEYINPUT62), .Z(n656) );
  XNOR2_X1 U517 ( .A(n738), .B(n739), .ZN(n417) );
  XNOR2_X1 U518 ( .A(n735), .B(n736), .ZN(n421) );
  INV_X1 U519 ( .A(KEYINPUT60), .ZN(n422) );
  XNOR2_X1 U520 ( .A(n728), .B(n466), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n730), .B(n729), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n456), .A2(n455), .ZN(n454) );
  XNOR2_X1 U523 ( .A(n471), .B(n359), .ZN(n456) );
  INV_X1 U524 ( .A(KEYINPUT53), .ZN(n469) );
  NAND2_X1 U525 ( .A1(n446), .A2(n445), .ZN(n444) );
  AND2_X1 U526 ( .A1(n480), .A2(KEYINPUT41), .ZN(n350) );
  AND2_X1 U527 ( .A1(n413), .A2(n412), .ZN(n351) );
  AND2_X1 U528 ( .A1(n605), .A2(n663), .ZN(n352) );
  AND2_X1 U529 ( .A1(n647), .A2(KEYINPUT83), .ZN(n353) );
  AND2_X1 U530 ( .A1(n370), .A2(n371), .ZN(n354) );
  AND2_X1 U531 ( .A1(G217), .A2(n566), .ZN(n355) );
  AND2_X1 U532 ( .A1(n547), .A2(G214), .ZN(n356) );
  XNOR2_X1 U533 ( .A(KEYINPUT6), .B(KEYINPUT106), .ZN(n357) );
  INV_X1 U534 ( .A(n663), .ZN(n387) );
  NAND2_X1 U535 ( .A1(n590), .A2(n585), .ZN(n712) );
  XNOR2_X1 U536 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n358) );
  XNOR2_X1 U537 ( .A(n661), .B(n660), .ZN(n359) );
  XOR2_X1 U538 ( .A(n732), .B(n731), .Z(n360) );
  INV_X1 U539 ( .A(n740), .ZN(n455) );
  XOR2_X1 U540 ( .A(KEYINPUT84), .B(KEYINPUT56), .Z(n361) );
  NAND2_X1 U541 ( .A1(n467), .A2(n414), .ZN(n639) );
  NAND2_X1 U542 ( .A1(n373), .A2(n372), .ZN(n369) );
  NAND2_X1 U543 ( .A1(n376), .A2(n442), .ZN(n375) );
  XNOR2_X1 U544 ( .A(n362), .B(n549), .ZN(n551) );
  NOR2_X1 U545 ( .A1(n732), .A2(G902), .ZN(n362) );
  NAND2_X1 U546 ( .A1(n591), .A2(n723), .ZN(n364) );
  XNOR2_X2 U547 ( .A(n527), .B(n499), .ZN(n595) );
  NAND2_X1 U548 ( .A1(n369), .A2(n354), .ZN(n377) );
  NAND2_X1 U549 ( .A1(n369), .A2(n365), .ZN(n376) );
  NOR2_X1 U550 ( .A1(n368), .A2(n366), .ZN(n365) );
  NAND2_X1 U551 ( .A1(n371), .A2(n367), .ZN(n366) );
  INV_X1 U552 ( .A(KEYINPUT83), .ZN(n367) );
  INV_X1 U553 ( .A(n370), .ZN(n368) );
  NAND2_X1 U554 ( .A1(n640), .A2(n378), .ZN(n371) );
  INV_X1 U555 ( .A(n640), .ZN(n372) );
  NOR2_X1 U556 ( .A1(n424), .A2(n378), .ZN(n373) );
  NAND2_X1 U557 ( .A1(n700), .A2(n383), .ZN(n382) );
  NOR2_X1 U558 ( .A1(n700), .A2(n386), .ZN(n384) );
  NAND2_X1 U559 ( .A1(n389), .A2(n387), .ZN(n494) );
  AND2_X1 U560 ( .A1(n389), .A2(n388), .ZN(n685) );
  INV_X1 U561 ( .A(n605), .ZN(n388) );
  XNOR2_X2 U562 ( .A(n391), .B(KEYINPUT45), .ZN(n744) );
  NAND2_X1 U563 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U564 ( .A(n394), .B(KEYINPUT44), .ZN(n392) );
  NOR2_X2 U565 ( .A1(n400), .A2(n765), .ZN(n394) );
  OR2_X1 U566 ( .A1(n595), .A2(n703), .ZN(n396) );
  XNOR2_X2 U567 ( .A(n532), .B(n501), .ZN(n409) );
  XNOR2_X2 U568 ( .A(n406), .B(G143), .ZN(n532) );
  NAND2_X1 U569 ( .A1(n411), .A2(n410), .ZN(n401) );
  NAND2_X1 U570 ( .A1(n403), .A2(n620), .ZN(n402) );
  NOR2_X1 U571 ( .A1(n693), .A2(n404), .ZN(n603) );
  XNOR2_X2 U572 ( .A(n404), .B(KEYINPUT1), .ZN(n694) );
  XNOR2_X2 U573 ( .A(n559), .B(G469), .ZN(n404) );
  XNOR2_X2 U574 ( .A(G128), .B(KEYINPUT76), .ZN(n406) );
  INV_X1 U575 ( .A(n467), .ZN(n768) );
  NOR2_X1 U576 ( .A1(n578), .A2(n358), .ZN(n410) );
  INV_X1 U577 ( .A(n586), .ZN(n411) );
  NAND2_X1 U578 ( .A1(n578), .A2(n358), .ZN(n412) );
  NAND2_X1 U579 ( .A1(n586), .A2(n358), .ZN(n413) );
  INV_X1 U580 ( .A(n767), .ZN(n414) );
  NAND2_X1 U581 ( .A1(n457), .A2(n350), .ZN(n479) );
  NAND2_X1 U582 ( .A1(n488), .A2(n582), .ZN(n487) );
  NAND2_X1 U583 ( .A1(n579), .A2(n626), .ZN(n586) );
  NOR2_X1 U584 ( .A1(n417), .A2(n740), .ZN(G66) );
  NOR2_X1 U585 ( .A1(n352), .A2(n614), .ZN(n419) );
  AND2_X2 U586 ( .A1(n473), .A2(n472), .ZN(n734) );
  NAND2_X1 U587 ( .A1(n734), .A2(G472), .ZN(n657) );
  NOR2_X1 U588 ( .A1(n420), .A2(n740), .ZN(G54) );
  NOR2_X1 U589 ( .A1(n421), .A2(n740), .ZN(G63) );
  NAND2_X1 U590 ( .A1(n744), .A2(n648), .ZN(n649) );
  XNOR2_X1 U591 ( .A(n454), .B(n361), .ZN(G51) );
  XNOR2_X1 U592 ( .A(n423), .B(n422), .ZN(G60) );
  NAND2_X1 U593 ( .A1(n453), .A2(n455), .ZN(n423) );
  NAND2_X1 U594 ( .A1(n602), .A2(n603), .ZN(n617) );
  NAND2_X1 U595 ( .A1(n690), .A2(n689), .ZN(n452) );
  XNOR2_X1 U596 ( .A(n688), .B(n425), .ZN(n440) );
  NAND2_X1 U597 ( .A1(n430), .A2(n429), .ZN(n428) );
  INV_X1 U598 ( .A(n629), .ZN(n429) );
  XNOR2_X1 U599 ( .A(n641), .B(n431), .ZN(n430) );
  INV_X1 U600 ( .A(KEYINPUT113), .ZN(n431) );
  NOR2_X1 U601 ( .A1(n655), .A2(n433), .ZN(n432) );
  AND2_X1 U602 ( .A1(n473), .A2(n440), .ZN(n689) );
  XNOR2_X2 U603 ( .A(n649), .B(n439), .ZN(n473) );
  INV_X1 U604 ( .A(KEYINPUT71), .ZN(n439) );
  XNOR2_X1 U605 ( .A(n491), .B(n441), .ZN(n490) );
  XNOR2_X2 U606 ( .A(n441), .B(KEYINPUT16), .ZN(n495) );
  XNOR2_X2 U607 ( .A(n506), .B(n507), .ZN(n441) );
  NAND2_X1 U608 ( .A1(n447), .A2(n444), .ZN(n470) );
  INV_X1 U609 ( .A(n452), .ZN(n446) );
  NOR2_X1 U610 ( .A1(n449), .A2(G953), .ZN(n448) );
  NAND2_X1 U611 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U612 ( .A(n733), .B(n360), .ZN(n453) );
  XNOR2_X1 U613 ( .A(n497), .B(KEYINPUT22), .ZN(n579) );
  XNOR2_X1 U614 ( .A(n687), .B(KEYINPUT81), .ZN(n690) );
  INV_X1 U615 ( .A(n714), .ZN(n457) );
  NAND2_X1 U616 ( .A1(n547), .A2(G210), .ZN(n459) );
  XOR2_X2 U617 ( .A(n558), .B(G122), .Z(n513) );
  XNOR2_X1 U618 ( .A(n612), .B(n611), .ZN(n464) );
  NOR2_X1 U619 ( .A1(n626), .A2(n625), .ZN(n627) );
  NAND2_X1 U620 ( .A1(n734), .A2(G475), .ZN(n733) );
  XNOR2_X2 U621 ( .A(n495), .B(n513), .ZN(n741) );
  XNOR2_X2 U622 ( .A(n503), .B(G101), .ZN(n507) );
  NAND2_X1 U623 ( .A1(n658), .A2(n455), .ZN(n489) );
  XNOR2_X1 U624 ( .A(n489), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X2 U625 ( .A(G113), .B(KEYINPUT88), .ZN(n503) );
  NAND2_X1 U626 ( .A1(n609), .A2(n608), .ZN(n625) );
  XNOR2_X1 U627 ( .A(n470), .B(n469), .ZN(G75) );
  INV_X1 U628 ( .A(n685), .ZN(n475) );
  NAND2_X1 U629 ( .A1(n476), .A2(n482), .ZN(n691) );
  AND2_X1 U630 ( .A1(n479), .A2(n481), .ZN(n476) );
  INV_X1 U631 ( .A(n712), .ZN(n480) );
  NAND2_X1 U632 ( .A1(n714), .A2(n483), .ZN(n482) );
  XNOR2_X2 U633 ( .A(n520), .B(n519), .ZN(n618) );
  XNOR2_X2 U634 ( .A(n512), .B(n511), .ZN(n558) );
  INV_X1 U635 ( .A(n618), .ZN(n645) );
  NOR2_X2 U636 ( .A1(n613), .A2(n526), .ZN(n527) );
  INV_X1 U637 ( .A(KEYINPUT69), .ZN(n615) );
  INV_X1 U638 ( .A(KEYINPUT89), .ZN(n514) );
  INV_X1 U639 ( .A(KEYINPUT103), .ZN(n533) );
  XNOR2_X1 U640 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U641 ( .A(KEYINPUT104), .B(G478), .ZN(n539) );
  INV_X1 U642 ( .A(n694), .ZN(n630) );
  NOR2_X1 U643 ( .A1(G952), .A2(n760), .ZN(n740) );
  INV_X1 U644 ( .A(KEYINPUT3), .ZN(n504) );
  NAND2_X1 U645 ( .A1(G234), .A2(n517), .ZN(n509) );
  XNOR2_X1 U646 ( .A(KEYINPUT20), .B(n509), .ZN(n571) );
  NAND2_X1 U647 ( .A1(n571), .A2(G221), .ZN(n510) );
  XOR2_X1 U648 ( .A(KEYINPUT21), .B(n510), .Z(n697) );
  XNOR2_X1 U649 ( .A(KEYINPUT70), .B(G110), .ZN(n511) );
  XNOR2_X1 U650 ( .A(n541), .B(KEYINPUT74), .ZN(n515) );
  NAND2_X1 U651 ( .A1(n659), .A2(n517), .ZN(n520) );
  AND2_X1 U652 ( .A1(G210), .A2(n521), .ZN(n518) );
  NAND2_X1 U653 ( .A1(G214), .A2(n521), .ZN(n709) );
  XNOR2_X1 U654 ( .A(n522), .B(KEYINPUT14), .ZN(n523) );
  NAND2_X1 U655 ( .A1(n523), .A2(G952), .ZN(n722) );
  NOR2_X1 U656 ( .A1(G953), .A2(n722), .ZN(n601) );
  NAND2_X1 U657 ( .A1(G902), .A2(n523), .ZN(n598) );
  INV_X1 U658 ( .A(G898), .ZN(n749) );
  NAND2_X1 U659 ( .A1(G953), .A2(n749), .ZN(n742) );
  NOR2_X1 U660 ( .A1(n598), .A2(n742), .ZN(n524) );
  NOR2_X1 U661 ( .A1(n601), .A2(n524), .ZN(n525) );
  XOR2_X1 U662 ( .A(KEYINPUT91), .B(n525), .Z(n526) );
  XNOR2_X1 U663 ( .A(n531), .B(n530), .ZN(n536) );
  XNOR2_X1 U664 ( .A(n532), .B(G134), .ZN(n534) );
  NAND2_X1 U665 ( .A1(G234), .A2(n760), .ZN(n537) );
  XNOR2_X1 U666 ( .A(n538), .B(n537), .ZN(n566) );
  NOR2_X1 U667 ( .A1(G902), .A2(n736), .ZN(n540) );
  XNOR2_X1 U668 ( .A(n542), .B(G131), .ZN(n546) );
  XNOR2_X1 U669 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U670 ( .A(n754), .B(n548), .ZN(n732) );
  XNOR2_X1 U671 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n549) );
  XOR2_X1 U672 ( .A(KEYINPUT13), .B(G475), .Z(n550) );
  XNOR2_X1 U673 ( .A(n551), .B(n550), .ZN(n589) );
  INV_X1 U674 ( .A(n589), .ZN(n585) );
  XOR2_X1 U675 ( .A(G101), .B(G146), .Z(n555) );
  NAND2_X1 U676 ( .A1(G227), .A2(n760), .ZN(n554) );
  XOR2_X1 U677 ( .A(KEYINPUT24), .B(G128), .Z(n561) );
  XNOR2_X1 U678 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U679 ( .A(KEYINPUT73), .B(KEYINPUT95), .Z(n562) );
  XNOR2_X1 U680 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U681 ( .A(n754), .B(n564), .ZN(n570) );
  XOR2_X1 U682 ( .A(n565), .B(KEYINPUT23), .Z(n568) );
  NAND2_X1 U683 ( .A1(G221), .A2(n566), .ZN(n567) );
  XNOR2_X1 U684 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U685 ( .A(n570), .B(n569), .ZN(n739) );
  XOR2_X1 U686 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n573) );
  NAND2_X1 U687 ( .A1(n571), .A2(G217), .ZN(n572) );
  XNOR2_X1 U688 ( .A(KEYINPUT72), .B(KEYINPUT97), .ZN(n574) );
  NOR2_X1 U689 ( .A1(n694), .A2(n696), .ZN(n577) );
  XNOR2_X1 U690 ( .A(n577), .B(KEYINPUT107), .ZN(n578) );
  NAND2_X1 U691 ( .A1(n694), .A2(n579), .ZN(n580) );
  NOR2_X1 U692 ( .A1(n700), .A2(n580), .ZN(n581) );
  NAND2_X1 U693 ( .A1(n609), .A2(n581), .ZN(n671) );
  NAND2_X1 U694 ( .A1(n696), .A2(n697), .ZN(n693) );
  INV_X1 U695 ( .A(n626), .ZN(n582) );
  INV_X1 U696 ( .A(KEYINPUT92), .ZN(n583) );
  XOR2_X1 U697 ( .A(KEYINPUT68), .B(KEYINPUT34), .Z(n584) );
  NOR2_X1 U698 ( .A1(n590), .A2(n585), .ZN(n620) );
  OR2_X1 U699 ( .A1(n630), .A2(n586), .ZN(n587) );
  XNOR2_X1 U700 ( .A(KEYINPUT105), .B(n679), .ZN(n605) );
  NAND2_X1 U701 ( .A1(n590), .A2(n589), .ZN(n663) );
  INV_X1 U702 ( .A(n603), .ZN(n593) );
  NAND2_X1 U703 ( .A1(n591), .A2(n610), .ZN(n592) );
  NOR2_X1 U704 ( .A1(n593), .A2(n592), .ZN(n668) );
  NAND2_X1 U705 ( .A1(n700), .A2(n594), .ZN(n703) );
  NOR2_X1 U706 ( .A1(n668), .A2(n680), .ZN(n596) );
  OR2_X1 U707 ( .A1(n352), .A2(n596), .ZN(n597) );
  OR2_X1 U708 ( .A1(n760), .A2(n598), .ZN(n599) );
  NOR2_X1 U709 ( .A1(G900), .A2(n599), .ZN(n600) );
  NOR2_X1 U710 ( .A1(n601), .A2(n600), .ZN(n607) );
  INV_X1 U711 ( .A(n697), .ZN(n606) );
  NOR2_X1 U712 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U713 ( .A(KEYINPUT65), .B(KEYINPUT47), .Z(n614) );
  XNOR2_X1 U714 ( .A(n616), .B(n615), .ZN(n624) );
  NAND2_X1 U715 ( .A1(KEYINPUT47), .A2(n352), .ZN(n621) );
  NOR2_X1 U716 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U717 ( .A1(n620), .A2(n619), .ZN(n674) );
  NAND2_X1 U718 ( .A1(n621), .A2(n674), .ZN(n622) );
  XNOR2_X1 U719 ( .A(KEYINPUT78), .B(n622), .ZN(n623) );
  NOR2_X1 U720 ( .A1(n624), .A2(n623), .ZN(n635) );
  XNOR2_X1 U721 ( .A(n627), .B(KEYINPUT109), .ZN(n628) );
  INV_X1 U722 ( .A(n675), .ZN(n631) );
  NAND2_X1 U723 ( .A1(KEYINPUT47), .A2(n631), .ZN(n632) );
  XNOR2_X1 U724 ( .A(KEYINPUT79), .B(n632), .ZN(n633) );
  NAND2_X1 U725 ( .A1(n635), .A2(n634), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n709), .ZN(n642) );
  NOR2_X1 U727 ( .A1(n630), .A2(n642), .ZN(n643) );
  XNOR2_X1 U728 ( .A(n643), .B(KEYINPUT43), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U730 ( .A(KEYINPUT110), .B(n646), .ZN(n766) );
  INV_X1 U731 ( .A(n766), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n686), .A2(n744), .ZN(n652) );
  INV_X1 U733 ( .A(KEYINPUT2), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U736 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n661) );
  XNOR2_X1 U737 ( .A(n659), .B(KEYINPUT86), .ZN(n660) );
  XNOR2_X1 U738 ( .A(G101), .B(n662), .ZN(G3) );
  NAND2_X1 U739 ( .A1(n387), .A2(n668), .ZN(n664) );
  XNOR2_X1 U740 ( .A(G104), .B(n664), .ZN(G6) );
  XOR2_X1 U741 ( .A(KEYINPUT27), .B(KEYINPUT115), .Z(n666) );
  XNOR2_X1 U742 ( .A(G107), .B(KEYINPUT114), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U744 ( .A(KEYINPUT26), .B(n667), .Z(n670) );
  NAND2_X1 U745 ( .A1(n668), .A2(n679), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n670), .B(n669), .ZN(G9) );
  XNOR2_X1 U747 ( .A(G110), .B(n671), .ZN(G12) );
  XOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U749 ( .A1(n675), .A2(n679), .ZN(n672) );
  XNOR2_X1 U750 ( .A(n673), .B(n672), .ZN(G30) );
  XNOR2_X1 U751 ( .A(G143), .B(n674), .ZN(G45) );
  NAND2_X1 U752 ( .A1(n675), .A2(n387), .ZN(n676) );
  XNOR2_X1 U753 ( .A(n676), .B(G146), .ZN(G48) );
  NAND2_X1 U754 ( .A1(n680), .A2(n387), .ZN(n677) );
  XNOR2_X1 U755 ( .A(n677), .B(KEYINPUT116), .ZN(n678) );
  XNOR2_X1 U756 ( .A(G113), .B(n678), .ZN(G15) );
  NAND2_X1 U757 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n681), .B(G116), .ZN(G18) );
  XOR2_X1 U759 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n683) );
  XNOR2_X1 U760 ( .A(G125), .B(KEYINPUT37), .ZN(n682) );
  XNOR2_X1 U761 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U762 ( .A(n500), .B(n684), .ZN(G27) );
  XOR2_X1 U763 ( .A(G134), .B(n685), .Z(G36) );
  NOR2_X1 U764 ( .A1(n744), .A2(KEYINPUT2), .ZN(n688) );
  XNOR2_X1 U765 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n692) );
  XNOR2_X1 U766 ( .A(n692), .B(KEYINPUT51), .ZN(n706) );
  NAND2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U768 ( .A(n695), .B(KEYINPUT50), .ZN(n702) );
  NOR2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U770 ( .A(KEYINPUT49), .B(n698), .Z(n699) );
  NOR2_X1 U771 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U773 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U774 ( .A(n706), .B(n705), .Z(n707) );
  NOR2_X1 U775 ( .A1(n691), .A2(n707), .ZN(n708) );
  XNOR2_X1 U776 ( .A(KEYINPUT121), .B(n708), .ZN(n719) );
  NOR2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U778 ( .A(KEYINPUT122), .B(n711), .Z(n713) );
  NAND2_X1 U779 ( .A1(n713), .A2(n480), .ZN(n716) );
  OR2_X1 U780 ( .A1(n352), .A2(n714), .ZN(n715) );
  NAND2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U782 ( .A1(n717), .A2(n723), .ZN(n718) );
  NAND2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U784 ( .A(KEYINPUT52), .B(n720), .Z(n721) );
  NOR2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n726) );
  INV_X1 U786 ( .A(n723), .ZN(n724) );
  NOR2_X1 U787 ( .A1(n691), .A2(n724), .ZN(n725) );
  NOR2_X1 U788 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U789 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n729) );
  NAND2_X1 U790 ( .A1(n737), .A2(G469), .ZN(n728) );
  INV_X1 U791 ( .A(KEYINPUT59), .ZN(n731) );
  NAND2_X1 U792 ( .A1(G478), .A2(n737), .ZN(n735) );
  NAND2_X1 U793 ( .A1(G217), .A2(n737), .ZN(n738) );
  XNOR2_X1 U794 ( .A(n741), .B(KEYINPUT126), .ZN(n743) );
  NAND2_X1 U795 ( .A1(n743), .A2(n742), .ZN(n753) );
  NAND2_X1 U796 ( .A1(n744), .A2(n760), .ZN(n745) );
  XNOR2_X1 U797 ( .A(n745), .B(KEYINPUT125), .ZN(n751) );
  XOR2_X1 U798 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n747) );
  NAND2_X1 U799 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U800 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U801 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U802 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U803 ( .A(n753), .B(n752), .ZN(G69) );
  XOR2_X1 U804 ( .A(n754), .B(n755), .Z(n759) );
  XOR2_X1 U805 ( .A(G227), .B(n759), .Z(n756) );
  NAND2_X1 U806 ( .A1(G900), .A2(n756), .ZN(n757) );
  NAND2_X1 U807 ( .A1(n757), .A2(G953), .ZN(n763) );
  XNOR2_X1 U808 ( .A(n759), .B(n758), .ZN(n761) );
  NAND2_X1 U809 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n763), .A2(n762), .ZN(G72) );
  XNOR2_X1 U811 ( .A(G119), .B(n764), .ZN(G21) );
  XOR2_X1 U812 ( .A(n765), .B(G122), .Z(G24) );
  XOR2_X1 U813 ( .A(G140), .B(n766), .Z(G42) );
  XOR2_X1 U814 ( .A(G131), .B(n767), .Z(G33) );
  XOR2_X1 U815 ( .A(G137), .B(n768), .Z(G39) );
endmodule

