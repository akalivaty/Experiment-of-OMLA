//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944;
  XNOR2_X1  g000(.A(G127gat), .B(G155gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G231gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  XNOR2_X1  g003(.A(G15gat), .B(G22gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT88), .ZN(new_n206));
  INV_X1    g005(.A(G15gat), .ZN(new_n207));
  INV_X1    g006(.A(G22gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT88), .ZN(new_n210));
  NAND2_X1  g009(.A1(G15gat), .A2(G22gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(KEYINPUT89), .A2(G1gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(KEYINPUT89), .A2(G1gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT16), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT90), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT90), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n218), .B(KEYINPUT16), .C1(new_n214), .C2(new_n215), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n213), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G8gat), .ZN(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n222), .A3(new_n212), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n221), .B1(new_n220), .B2(new_n223), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT96), .ZN(new_n227));
  AND2_X1   g026(.A1(G71gat), .A2(G78gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(G71gat), .A2(G78gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OR2_X1    g030(.A1(G57gat), .A2(G64gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(G57gat), .A2(G64gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(new_n233), .C1(new_n228), .C2(KEYINPUT9), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n229), .A2(KEYINPUT95), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n227), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(new_n235), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n230), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n236), .A3(KEYINPUT96), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(KEYINPUT21), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G183gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n237), .A2(new_n238), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(KEYINPUT21), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G183gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n226), .A2(new_n250), .A3(new_n243), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT97), .B(G211gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(KEYINPUT98), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n256));
  XOR2_X1   g055(.A(new_n255), .B(new_n256), .Z(new_n257));
  AOI21_X1  g056(.A(new_n249), .B1(new_n245), .B2(new_n251), .ZN(new_n258));
  OR3_X1    g057(.A1(new_n253), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n253), .B2(new_n258), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n204), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n259), .A2(new_n204), .A3(new_n260), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT101), .ZN(new_n265));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266));
  INV_X1    g065(.A(G85gat), .ZN(new_n267));
  INV_X1    g066(.A(G92gat), .ZN(new_n268));
  AOI22_X1  g067(.A1(KEYINPUT8), .A2(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G99gat), .B(G106gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT7), .ZN(new_n271));
  OAI22_X1  g070(.A1(new_n267), .A2(new_n268), .B1(new_n271), .B2(KEYINPUT99), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT99), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n269), .A2(new_n270), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n275), .A2(KEYINPUT100), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(KEYINPUT100), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n265), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n272), .A2(new_n274), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT100), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n279), .A2(new_n280), .A3(new_n270), .A4(new_n269), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n275), .A2(KEYINPUT100), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT101), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n266), .A2(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n268), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n272), .A2(new_n274), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n270), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT102), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n286), .A2(KEYINPUT102), .A3(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n278), .A2(new_n283), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT17), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT14), .ZN(new_n296));
  INV_X1    g095(.A(G29gat), .ZN(new_n297));
  INV_X1    g096(.A(G36gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n299), .A2(new_n300), .B1(G29gat), .B2(G36gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n302));
  XNOR2_X1  g101(.A(G43gat), .B(G50gat), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n301), .A2(new_n302), .B1(KEYINPUT15), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g103(.A(G43gat), .B(G50gat), .Z(new_n305));
  INV_X1    g104(.A(KEYINPUT15), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n301), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n305), .A2(new_n306), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n301), .B(new_n307), .C1(new_n310), .C2(new_n302), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n295), .B(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G190gat), .B(G218gat), .ZN(new_n316));
  OR2_X1    g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G134gat), .B(G162gat), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n318), .B(new_n319), .Z(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n316), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n320), .B1(new_n317), .B2(new_n321), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n264), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT67), .B(G134gat), .Z(new_n327));
  INV_X1    g126(.A(G127gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(G134gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G113gat), .B(G120gat), .ZN(new_n333));
  OAI22_X1  g132(.A1(new_n329), .A2(new_n332), .B1(KEYINPUT1), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G134gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT1), .B1(new_n337), .B2(G127gat), .ZN(new_n338));
  INV_X1    g137(.A(G113gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n340));
  NAND4_X1  g139(.A1(new_n336), .A2(new_n330), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n334), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343));
  INV_X1    g142(.A(G141gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(G148gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(KEYINPUT76), .B(G148gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n345), .B1(new_n346), .B2(new_n344), .ZN(new_n347));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348));
  OR2_X1    g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(KEYINPUT2), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT75), .B(KEYINPUT2), .Z(new_n352));
  XNOR2_X1  g151(.A(G141gat), .B(G148gat), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n348), .B(new_n349), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(new_n343), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n351), .A2(new_n354), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(KEYINPUT3), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n361));
  OAI221_X1 g160(.A(new_n342), .B1(new_n343), .B2(new_n355), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n342), .A2(new_n359), .ZN(new_n363));
  XOR2_X1   g162(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(KEYINPUT4), .B2(new_n363), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n334), .A2(new_n341), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n355), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n342), .A2(new_n359), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n367), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n368), .A2(KEYINPUT5), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  OR2_X1    g176(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n364), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n373), .A2(KEYINPUT5), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n362), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G1gat), .B(G29gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n383), .B(new_n267), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G57gat), .ZN(new_n385));
  XOR2_X1   g184(.A(new_n384), .B(new_n385), .Z(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(KEYINPUT6), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT6), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n382), .B2(new_n386), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n386), .B(KEYINPUT82), .Z(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n377), .B2(new_n381), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n387), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G183gat), .A2(G190gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT24), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(G183gat), .B2(G190gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(G169gat), .A2(G176gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n397), .B(KEYINPUT23), .Z(new_n398));
  NAND3_X1  g197(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(KEYINPUT25), .Z(new_n400));
  NAND2_X1  g199(.A1(new_n250), .A2(KEYINPUT27), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT64), .ZN(new_n402));
  AOI21_X1  g201(.A(G190gat), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n250), .A2(KEYINPUT27), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n403), .B(new_n404), .C1(new_n402), .C2(new_n401), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n406));
  AND2_X1   g205(.A1(new_n404), .A2(new_n401), .ZN(new_n407));
  INV_X1    g206(.A(G190gat), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n408), .A2(KEYINPUT28), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n405), .A2(new_n406), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT66), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT26), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(new_n412), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n411), .B(new_n413), .C1(new_n412), .C2(new_n397), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n413), .A2(new_n411), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n410), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n393), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G197gat), .B(G204gat), .ZN(new_n422));
  AND2_X1   g221(.A1(G211gat), .A2(G218gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n422), .B1(KEYINPUT22), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G211gat), .B(G218gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n400), .A2(new_n417), .A3(G226gat), .A4(G233gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n427), .B1(new_n421), .B2(new_n428), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT72), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(KEYINPUT73), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n426), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(new_n429), .A3(new_n436), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT73), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n435), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n430), .B2(new_n431), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n437), .A2(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n439), .A2(new_n429), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n448), .B(new_n443), .C1(KEYINPUT74), .C2(KEYINPUT30), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n392), .A2(new_n446), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n419), .B1(new_n358), .B2(new_n361), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n426), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n343), .B1(new_n426), .B2(KEYINPUT29), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n359), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(G22gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(G228gat), .A2(G233gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n356), .A2(new_n357), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT29), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n208), .B(new_n456), .C1(new_n464), .C2(new_n427), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n458), .A2(new_n459), .A3(new_n461), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT80), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n459), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n208), .B1(new_n454), .B2(new_n456), .ZN(new_n469));
  INV_X1    g268(.A(new_n465), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT31), .B(G50gat), .Z(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n466), .A2(new_n471), .A3(new_n467), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G78gat), .B(G106gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n474), .A2(new_n478), .A3(new_n476), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n418), .A2(new_n342), .ZN(new_n483));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n400), .A2(new_n369), .A3(new_n417), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(G15gat), .B(G43gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT70), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(G71gat), .ZN(new_n489));
  INV_X1    g288(.A(G99gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n484), .B1(new_n483), .B2(new_n485), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n486), .B(new_n491), .C1(new_n492), .C2(KEYINPUT33), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n483), .A2(new_n485), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT33), .ZN(new_n495));
  INV_X1    g294(.A(new_n491), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n494), .B(new_n484), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT32), .B(new_n499), .C1(new_n494), .C2(new_n484), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT32), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT34), .B1(new_n492), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n500), .A2(new_n493), .A3(new_n497), .A4(new_n502), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT85), .ZN(new_n507));
  INV_X1    g306(.A(new_n386), .ZN(new_n508));
  AOI211_X1 g307(.A(new_n388), .B(new_n508), .C1(new_n377), .C2(new_n381), .ZN(new_n509));
  INV_X1    g308(.A(new_n381), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n374), .A2(KEYINPUT79), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT5), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n510), .B1(new_n514), .B2(new_n368), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT6), .B1(new_n515), .B2(new_n508), .ZN(new_n516));
  INV_X1    g315(.A(new_n391), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n444), .A2(new_n445), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT73), .B1(new_n432), .B2(new_n436), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n440), .A2(new_n441), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n449), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT84), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n452), .A2(new_n482), .A3(new_n507), .A4(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n506), .B1(new_n480), .B2(new_n481), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n382), .A2(new_n386), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n509), .B1(new_n516), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(new_n522), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n524), .B1(new_n451), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n448), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n439), .A2(KEYINPUT37), .A3(new_n429), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n435), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n534), .A2(KEYINPUT38), .B1(new_n448), .B2(new_n443), .ZN(new_n535));
  INV_X1    g334(.A(new_n532), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT38), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n533), .A2(new_n537), .A3(new_n436), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n535), .B(new_n518), .C1(new_n536), .C2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT83), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n362), .A2(new_n378), .A3(new_n379), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(new_n373), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n540), .A3(new_n373), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n370), .A2(new_n367), .A3(new_n371), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n543), .A2(KEYINPUT39), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT39), .ZN(new_n547));
  INV_X1    g346(.A(new_n544), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(new_n542), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n549), .A3(new_n390), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT40), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n546), .A2(new_n549), .A3(KEYINPUT40), .A4(new_n390), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(new_n522), .A3(new_n517), .A4(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n482), .A2(new_n539), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n506), .A2(KEYINPUT71), .A3(KEYINPUT36), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT36), .B1(new_n506), .B2(KEYINPUT71), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n480), .B(new_n481), .C1(new_n527), .C2(new_n522), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n326), .B1(new_n530), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n309), .A2(new_n311), .A3(new_n294), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT91), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n226), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n220), .A2(new_n223), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(G8gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT17), .B1(new_n568), .B2(KEYINPUT91), .ZN(new_n569));
  INV_X1    g368(.A(new_n312), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n564), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT92), .Z(new_n573));
  AOI21_X1  g372(.A(KEYINPUT18), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(KEYINPUT91), .B1(new_n224), .B2(new_n225), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n575), .B2(new_n294), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(new_n577));
  OAI211_X1 g376(.A(KEYINPUT18), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n573), .B(KEYINPUT13), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n568), .A2(KEYINPUT93), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT93), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n584), .A3(new_n567), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n312), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n570), .B1(new_n568), .B2(KEYINPUT93), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G169gat), .B(G197gat), .Z(new_n589));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT12), .Z(new_n594));
  NAND4_X1  g393(.A1(new_n580), .A2(KEYINPUT94), .A3(new_n588), .A4(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n598), .A2(new_n588), .A3(new_n578), .A4(new_n594), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT94), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n580), .A2(new_n588), .ZN(new_n602));
  INV_X1    g401(.A(new_n594), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n595), .A2(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n278), .A2(new_n246), .A3(new_n283), .A4(new_n292), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n288), .A2(KEYINPUT103), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n286), .A2(new_n607), .A3(new_n287), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n606), .B(new_n608), .C1(new_n276), .C2(new_n277), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n247), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(KEYINPUT10), .B1(new_n605), .B2(new_n610), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n239), .A2(KEYINPUT10), .A3(new_n242), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n293), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n612), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT104), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT104), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n622), .B(new_n612), .C1(new_n617), .C2(new_n619), .ZN(new_n623));
  AOI211_X1 g422(.A(new_n613), .B(new_n616), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n620), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n616), .B1(new_n626), .B2(new_n613), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n604), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n561), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n527), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n222), .ZN(G1324gat));
  INV_X1    g432(.A(new_n522), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n635), .A2(KEYINPUT105), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(KEYINPUT105), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT16), .B(G8gat), .Z(new_n638));
  OAI211_X1 g437(.A(new_n636), .B(new_n637), .C1(KEYINPUT42), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n640), .B2(G8gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(KEYINPUT42), .A3(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(G1325gat));
  NOR3_X1   g442(.A1(new_n630), .A2(new_n207), .A3(new_n558), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n561), .A2(new_n629), .A3(new_n507), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n644), .B1(new_n207), .B2(new_n645), .ZN(G1326gat));
  NOR2_X1   g445(.A1(new_n630), .A2(new_n482), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT43), .B(G22gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(G1327gat));
  NAND3_X1  g448(.A1(new_n523), .A2(new_n450), .A3(new_n451), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n480), .A2(new_n481), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT85), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n506), .B(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n451), .B1(new_n525), .B2(new_n528), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n560), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n324), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n629), .A2(new_n264), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n297), .A3(new_n527), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT106), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT45), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n656), .A2(new_n324), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT108), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n657), .A2(KEYINPUT44), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n656), .A2(new_n668), .A3(new_n324), .A4(new_n664), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n658), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(G29gat), .B1(new_n672), .B2(new_n631), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n661), .A2(new_n662), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n663), .A2(new_n673), .A3(new_n674), .ZN(G1328gat));
  OR3_X1    g474(.A1(new_n672), .A2(KEYINPUT110), .A3(new_n634), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT110), .B1(new_n672), .B2(new_n634), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(G36gat), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(G36gat), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n659), .A2(new_n522), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n682), .ZN(G1329gat));
  NOR4_X1   g482(.A1(new_n657), .A2(G43gat), .A3(new_n653), .A4(new_n658), .ZN(new_n684));
  INV_X1    g483(.A(new_n558), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n685), .A3(new_n671), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(G43gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g487(.A(KEYINPUT48), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(KEYINPUT111), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n670), .A2(new_n651), .A3(new_n671), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G50gat), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(KEYINPUT111), .ZN(new_n693));
  NOR4_X1   g492(.A1(new_n657), .A2(G50gat), .A3(new_n482), .A4(new_n658), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AND4_X1   g494(.A1(new_n690), .A2(new_n692), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n694), .B1(new_n691), .B2(G50gat), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n690), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(G1331gat));
  NAND2_X1  g498(.A1(new_n602), .A2(new_n603), .ZN(new_n700));
  INV_X1    g499(.A(new_n601), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n599), .A2(new_n600), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n628), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n561), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n527), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g508(.A(new_n634), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n561), .A2(KEYINPUT112), .A3(new_n705), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT112), .B1(new_n561), .B2(new_n705), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT113), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n713), .A2(KEYINPUT113), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n715), .A2(new_n716), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n717));
  INV_X1    g516(.A(new_n716), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n718), .A2(new_n714), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(G1333gat));
  NOR3_X1   g520(.A1(new_n706), .A2(G71gat), .A3(new_n653), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n685), .B1(new_n711), .B2(new_n712), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n722), .B1(new_n723), .B2(G71gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT50), .ZN(G1334gat));
  OAI21_X1  g524(.A(new_n651), .B1(new_n711), .B2(new_n712), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G78gat), .ZN(G1335gat));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728));
  OR2_X1    g527(.A1(new_n322), .A2(new_n323), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n530), .B2(new_n560), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n264), .A2(new_n604), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n657), .A2(KEYINPUT51), .A3(new_n731), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n733), .A2(new_n734), .A3(new_n704), .ZN(new_n735));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n527), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n731), .A2(new_n704), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n670), .A2(new_n737), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n738), .A2(new_n267), .A3(new_n631), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n736), .A2(new_n739), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n738), .B2(new_n634), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n735), .A2(new_n268), .A3(new_n522), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT52), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n738), .B2(new_n558), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n735), .A2(new_n490), .A3(new_n507), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n670), .A2(new_n651), .A3(new_n737), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G106gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT114), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n733), .A2(new_n734), .ZN(new_n754));
  INV_X1    g553(.A(G106gat), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n754), .A2(new_n755), .A3(new_n628), .A4(new_n651), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n753), .A2(new_n757), .A3(KEYINPUT53), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n752), .B(new_n756), .C1(KEYINPUT114), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1339gat));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762));
  INV_X1    g561(.A(new_n263), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n261), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n729), .A2(new_n764), .A3(new_n604), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n765), .B2(new_n628), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n325), .A2(KEYINPUT115), .A3(new_n604), .A4(new_n704), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n616), .B1(new_n620), .B2(KEYINPUT54), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n621), .A2(new_n623), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT10), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n611), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n612), .ZN(new_n773));
  OR2_X1    g572(.A1(new_n293), .A2(new_n618), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n617), .A2(new_n619), .A3(new_n612), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(KEYINPUT116), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n770), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n770), .A2(KEYINPUT117), .A3(new_n780), .A4(new_n777), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n769), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n624), .B1(new_n785), .B2(KEYINPUT55), .ZN(new_n786));
  INV_X1    g585(.A(new_n769), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n772), .A2(KEYINPUT116), .A3(new_n773), .A4(new_n774), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n621), .B2(new_n623), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT117), .B1(new_n790), .B2(new_n777), .ZN(new_n791));
  INV_X1    g590(.A(new_n784), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n595), .A2(new_n601), .ZN(new_n796));
  INV_X1    g595(.A(new_n593), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n571), .A2(new_n573), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n586), .A2(new_n582), .A3(new_n587), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n795), .A3(new_n324), .A4(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n796), .A2(new_n628), .A3(new_n800), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n604), .B1(new_n793), .B2(new_n794), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(new_n786), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n805), .B2(new_n324), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n768), .B1(new_n806), .B2(new_n264), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(new_n651), .A3(new_n653), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n631), .A2(new_n522), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n339), .B1(new_n811), .B2(new_n703), .ZN(new_n812));
  INV_X1    g611(.A(new_n525), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n809), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n815), .A2(G113gat), .A3(new_n604), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n812), .A2(new_n816), .ZN(G1340gat));
  OAI21_X1  g616(.A(G120gat), .B1(new_n810), .B2(new_n704), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n815), .A2(G120gat), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n704), .ZN(G1341gat));
  OAI21_X1  g619(.A(new_n328), .B1(new_n815), .B2(new_n264), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n764), .A2(G127gat), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n821), .B1(new_n810), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT118), .Z(G1342gat));
  NOR3_X1   g623(.A1(new_n815), .A2(new_n327), .A3(new_n729), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n810), .B2(new_n729), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n826), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  INV_X1    g629(.A(new_n803), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n625), .B1(new_n793), .B2(new_n794), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n703), .B1(new_n785), .B2(KEYINPUT55), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n729), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n764), .B1(new_n835), .B2(new_n802), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n651), .B1(new_n836), .B2(new_n768), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n558), .A2(new_n809), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n840), .A2(G141gat), .A3(new_n604), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(KEYINPUT58), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n805), .B2(new_n324), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n834), .A2(KEYINPUT119), .A3(new_n729), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n845), .A3(new_n802), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n768), .B1(new_n846), .B2(new_n264), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT57), .B1(new_n847), .B2(new_n482), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n807), .A2(new_n482), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n838), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n848), .A2(new_n851), .A3(new_n703), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n842), .B1(new_n344), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n848), .A2(new_n851), .A3(KEYINPUT120), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT120), .B1(new_n848), .B2(new_n851), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n703), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n841), .B1(new_n856), .B2(G141gat), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n853), .B1(new_n857), .B2(new_n858), .ZN(G1344gat));
  OAI21_X1  g658(.A(new_n628), .B1(new_n854), .B2(new_n855), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(new_n346), .ZN(new_n862));
  INV_X1    g661(.A(G148gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n837), .A2(KEYINPUT57), .ZN(new_n864));
  INV_X1    g663(.A(new_n838), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n765), .A2(new_n628), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n850), .B(new_n651), .C1(new_n836), .C2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n864), .A2(new_n628), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n862), .A2(new_n872), .ZN(new_n873));
  OR3_X1    g672(.A1(new_n840), .A2(new_n346), .A3(new_n704), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1345gat));
  AOI21_X1  g674(.A(G155gat), .B1(new_n839), .B2(new_n764), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n854), .A2(new_n855), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n264), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n878), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g678(.A(G162gat), .B1(new_n839), .B2(new_n324), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n877), .A2(new_n729), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(G162gat), .ZN(G1347gat));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n807), .B2(new_n527), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n631), .C1(new_n836), .C2(new_n768), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n813), .B(new_n634), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(G169gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n703), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n634), .A2(new_n527), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n808), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G169gat), .B1(new_n890), .B2(new_n604), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n888), .A2(new_n891), .ZN(G1348gat));
  OAI21_X1  g691(.A(G176gat), .B1(new_n890), .B2(new_n704), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n886), .A2(new_n628), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(G176gat), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT123), .ZN(G1349gat));
  AOI21_X1  g695(.A(new_n813), .B1(new_n884), .B2(new_n885), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n897), .A2(new_n407), .A3(new_n522), .A4(new_n764), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n886), .A2(KEYINPUT124), .A3(new_n407), .A4(new_n764), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G183gat), .B1(new_n890), .B2(new_n264), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT60), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n906), .A3(new_n903), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n890), .B2(new_n729), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT61), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n886), .A2(new_n408), .A3(new_n324), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1351gat));
  NAND2_X1  g711(.A1(new_n884), .A2(new_n885), .ZN(new_n913));
  AND4_X1   g712(.A1(new_n651), .A2(new_n913), .A3(new_n522), .A4(new_n558), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(KEYINPUT125), .ZN(new_n916));
  XOR2_X1   g715(.A(KEYINPUT126), .B(G197gat), .Z(new_n917));
  NOR2_X1   g716(.A1(new_n604), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n864), .A2(new_n867), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n558), .A2(new_n889), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n922), .B2(new_n604), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n919), .A2(new_n923), .ZN(G1352gat));
  INV_X1    g723(.A(G204gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n914), .A2(new_n925), .A3(new_n628), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n920), .A2(new_n628), .A3(new_n921), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n927), .B(new_n928), .C1(new_n925), .C2(new_n929), .ZN(G1353gat));
  NOR2_X1   g729(.A1(new_n264), .A2(G211gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G211gat), .B1(new_n922), .B2(new_n264), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT127), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n920), .A2(new_n939), .A3(new_n921), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n324), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G218gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n729), .A2(G218gat), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n915), .A2(new_n916), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1355gat));
endmodule


