//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n207), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  OR2_X1    g0014(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n207), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n215), .A2(new_n218), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n214), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XOR2_X1   g0037(.A(G58), .B(G77), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n221), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G33), .ZN(new_n247));
  NOR2_X1   g0047(.A1(new_n247), .A2(G20), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT67), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT67), .B1(new_n247), .B2(G20), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G77), .A3(new_n251), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G68), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n246), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(KEYINPUT11), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT68), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT68), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n261), .A2(new_n258), .A3(G13), .A4(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n246), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n222), .A2(G1), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n264), .A2(new_n254), .A3(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n257), .A2(new_n266), .ZN(new_n267));
  OR3_X1    g0067(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n268));
  OAI21_X1  g0068(.A(KEYINPUT12), .B1(new_n263), .B2(G68), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n256), .A2(KEYINPUT11), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT77), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n257), .A2(new_n266), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT77), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(new_n271), .A4(new_n270), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  OAI211_X1 g0079(.A(G232), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  OAI211_X1 g0081(.A(G226), .B(new_n281), .C1(new_n278), .C2(new_n279), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G97), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(new_n221), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(G1), .A2(G13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(G274), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n290), .A2(G238), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT75), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n294), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n294), .B2(new_n296), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n287), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT13), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n302), .B(new_n287), .C1(new_n298), .C2(new_n299), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(G179), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n301), .A2(KEYINPUT76), .A3(new_n303), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n298), .A2(new_n299), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT76), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n307), .A2(new_n308), .A3(new_n302), .A4(new_n287), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(G169), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT14), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(KEYINPUT78), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n305), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n312), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n306), .A2(new_n309), .A3(G169), .A4(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n277), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n317), .B1(new_n300), .B2(KEYINPUT13), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n273), .A2(new_n276), .B1(new_n303), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n306), .A2(G200), .A3(new_n309), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT16), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT3), .B(G33), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(G20), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n278), .A2(new_n279), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n254), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G58), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n254), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G58), .A2(G68), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n253), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n324), .B1(new_n330), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT7), .B1(new_n328), .B2(new_n222), .ZN(new_n338));
  NOR4_X1   g0138(.A1(new_n278), .A2(new_n279), .A3(new_n325), .A4(G20), .ZN(new_n339));
  OAI21_X1  g0139(.A(G68), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n336), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(KEYINPUT16), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n342), .A3(new_n245), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT66), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT8), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n345), .A2(G58), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n331), .A2(KEYINPUT8), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n331), .A2(KEYINPUT8), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(G58), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT66), .ZN(new_n351));
  INV_X1    g0151(.A(new_n265), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n264), .B1(KEYINPUT79), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT79), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n348), .A2(new_n355), .A3(new_n351), .A4(new_n352), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n348), .A2(new_n351), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n260), .A2(new_n262), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n354), .A2(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n290), .A2(new_n295), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n294), .B1(new_n361), .B2(new_n228), .ZN(new_n362));
  OAI211_X1 g0162(.A(G223), .B(new_n281), .C1(new_n278), .C2(new_n279), .ZN(new_n363));
  OAI211_X1 g0163(.A(G226), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n364));
  INV_X1    g0164(.A(G87), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n363), .B(new_n364), .C1(new_n247), .C2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n286), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(KEYINPUT80), .B(G190), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n366), .A2(new_n286), .ZN(new_n371));
  INV_X1    g0171(.A(new_n362), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n343), .A2(new_n360), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n375), .B(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n353), .A2(KEYINPUT79), .ZN(new_n378));
  INV_X1    g0178(.A(new_n264), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n356), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n358), .A2(new_n359), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n340), .A2(new_n341), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n246), .B1(new_n383), .B2(new_n324), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n382), .B1(new_n384), .B2(new_n342), .ZN(new_n385));
  INV_X1    g0185(.A(G179), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n367), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(G169), .B2(new_n367), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT18), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n343), .A2(new_n360), .ZN(new_n390));
  AOI21_X1  g0190(.A(G169), .B1(new_n371), .B2(new_n372), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n386), .B2(new_n367), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n377), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n323), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT9), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT72), .ZN(new_n399));
  INV_X1    g0199(.A(G150), .ZN(new_n400));
  INV_X1    g0200(.A(new_n253), .ZN(new_n401));
  OAI22_X1  g0201(.A1(new_n400), .A2(new_n401), .B1(new_n201), .B2(new_n222), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n250), .A2(new_n251), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(new_n357), .B2(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n404), .A2(new_n246), .ZN(new_n405));
  INV_X1    g0205(.A(G50), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n265), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n263), .A2(new_n246), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G50), .B2(new_n263), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n399), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n404), .A2(new_n246), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n412), .A2(KEYINPUT72), .A3(new_n409), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n398), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n326), .A2(G222), .A3(new_n281), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n326), .A2(G1698), .ZN(new_n416));
  INV_X1    g0216(.A(G223), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n415), .B1(new_n202), .B2(new_n326), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n286), .ZN(new_n419));
  INV_X1    g0219(.A(new_n294), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n286), .A2(new_n293), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(G226), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(G190), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n405), .A2(new_n399), .A3(new_n410), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT72), .B1(new_n412), .B2(new_n409), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(KEYINPUT9), .A3(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n414), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n419), .A2(new_n422), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G200), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n429), .C1(KEYINPUT73), .C2(KEYINPUT10), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n414), .A2(new_n429), .A3(new_n423), .A4(new_n426), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n414), .A2(KEYINPUT73), .A3(new_n423), .A4(new_n426), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT10), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(G169), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n405), .A2(new_n410), .B1(new_n428), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(G179), .B2(new_n428), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n326), .A2(G232), .A3(new_n281), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n326), .A2(G238), .A3(G1698), .ZN(new_n440));
  INV_X1    g0240(.A(G107), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n439), .B(new_n440), .C1(new_n441), .C2(new_n326), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n286), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT69), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n420), .B1(G244), .B2(new_n421), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n443), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g0248(.A(G190), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n346), .A2(new_n347), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT70), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n401), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(new_n451), .B2(new_n401), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT15), .B(G87), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(new_n248), .B1(G20), .B2(G77), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n246), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n264), .A2(new_n202), .A3(new_n265), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n263), .A2(G77), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n443), .A2(new_n445), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(G200), .A3(new_n446), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n449), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G179), .B1(new_n462), .B2(new_n446), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n462), .A2(new_n436), .A3(new_n446), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(KEYINPUT71), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n460), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n386), .B1(new_n447), .B2(new_n448), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT71), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n464), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n435), .A2(KEYINPUT74), .A3(new_n438), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT74), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n430), .A2(new_n434), .A3(new_n438), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n475), .B1(new_n476), .B2(new_n472), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n397), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n292), .A2(G1), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(G274), .B1(new_n285), .B2(new_n221), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT81), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G274), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n486), .B1(new_n288), .B2(new_n289), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT81), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n487), .A2(new_n488), .A3(new_n489), .A4(new_n480), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n489), .A2(new_n480), .B1(new_n288), .B2(new_n289), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n485), .A2(new_n490), .B1(new_n491), .B2(G257), .ZN(new_n492));
  OAI211_X1 g0292(.A(G244), .B(new_n281), .C1(new_n278), .C2(new_n279), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G250), .A2(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(KEYINPUT4), .A2(G244), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(G1698), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n497), .B1(new_n326), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n286), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n492), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G200), .ZN(new_n505));
  INV_X1    g0305(.A(G97), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n359), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n258), .A2(G33), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n263), .A2(G97), .A3(new_n246), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(G107), .B1(new_n338), .B2(new_n339), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT6), .ZN(new_n512));
  AND2_X1   g0312(.A1(G97), .A2(G107), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n512), .B1(new_n513), .B2(new_n204), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n441), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n510), .B1(new_n518), .B2(new_n245), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n492), .A2(new_n503), .A3(G190), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n505), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n485), .A2(new_n490), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n491), .A2(G257), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n290), .B1(new_n495), .B2(new_n501), .ZN(new_n525));
  OAI21_X1  g0325(.A(G169), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n492), .A2(new_n503), .A3(G179), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT82), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n326), .A2(G244), .A3(G1698), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G33), .A2(G116), .ZN(new_n531));
  OAI211_X1 g0331(.A(G238), .B(new_n281), .C1(new_n278), .C2(new_n279), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n286), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT83), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n258), .A2(G45), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G250), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n535), .B1(new_n286), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n290), .A2(KEYINPUT83), .A3(G250), .A4(new_n536), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n538), .A2(new_n539), .B1(new_n487), .B2(new_n480), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(G200), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n222), .B1(new_n283), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G87), .B2(new_n205), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n326), .A2(new_n222), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n222), .A2(G33), .A3(G97), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n547), .A2(KEYINPUT84), .A3(new_n543), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT84), .B1(new_n547), .B2(new_n543), .ZN(new_n549));
  OAI221_X1 g0349(.A(new_n545), .B1(new_n546), .B2(new_n254), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n550), .A2(new_n245), .B1(new_n359), .B2(new_n454), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n263), .A2(new_n246), .A3(new_n508), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G87), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n534), .A2(new_n540), .A3(G190), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n542), .A2(new_n551), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n541), .A2(new_n436), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n455), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n545), .B1(new_n546), .B2(new_n254), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n548), .A2(new_n549), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n245), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n359), .A2(new_n454), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n534), .A2(new_n540), .A3(new_n386), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n555), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n505), .A2(new_n519), .A3(new_n520), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n529), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n222), .B(G87), .C1(new_n278), .C2(new_n279), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT22), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT22), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n326), .A2(new_n573), .A3(new_n222), .A4(G87), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  OR3_X1    g0375(.A1(new_n531), .A2(KEYINPUT86), .A3(G20), .ZN(new_n576));
  OR3_X1    g0376(.A1(new_n222), .A2(KEYINPUT23), .A3(G107), .ZN(new_n577));
  OAI21_X1  g0377(.A(KEYINPUT86), .B1(new_n531), .B2(G20), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT23), .B1(new_n222), .B2(G107), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n575), .B2(new_n580), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n245), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT25), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n263), .B2(G107), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n359), .A2(KEYINPUT25), .A3(new_n441), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(new_n552), .B2(G107), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G257), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n590));
  OAI211_X1 g0390(.A(G250), .B(new_n281), .C1(new_n278), .C2(new_n279), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G294), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT87), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT87), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n590), .A2(new_n591), .A3(new_n595), .A4(new_n592), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n286), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n491), .A2(G264), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n522), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n436), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n589), .B(new_n600), .C1(G179), .C2(new_n599), .ZN(new_n601));
  INV_X1    g0401(.A(G116), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n359), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n263), .A2(G116), .A3(new_n246), .A4(new_n508), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n244), .A2(new_n221), .B1(G20), .B2(new_n602), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n496), .B(new_n222), .C1(G33), .C2(new_n506), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n606), .A2(KEYINPUT20), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT20), .B1(new_n606), .B2(new_n607), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n485), .A2(new_n490), .B1(new_n491), .B2(G270), .ZN(new_n612));
  OAI211_X1 g0412(.A(G264), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n613));
  OAI211_X1 g0413(.A(G257), .B(new_n281), .C1(new_n278), .C2(new_n279), .ZN(new_n614));
  OR2_X1    g0414(.A1(KEYINPUT3), .A2(G33), .ZN(new_n615));
  NAND2_X1  g0415(.A1(KEYINPUT3), .A2(G33), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(G303), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n613), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n286), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n612), .A2(new_n369), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n611), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G200), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n612), .B2(new_n619), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT85), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n623), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(new_n626), .A3(new_n611), .A4(new_n620), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n491), .A2(G270), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n522), .A2(new_n619), .A3(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n603), .B(new_n604), .C1(new_n609), .C2(new_n608), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G179), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n612), .A2(new_n619), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n633), .A2(new_n631), .A3(KEYINPUT21), .A4(G169), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n436), .B1(new_n612), .B2(new_n619), .ZN(new_n636));
  AOI21_X1  g0436(.A(KEYINPUT21), .B1(new_n636), .B2(new_n631), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n599), .A2(G200), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n290), .B1(new_n593), .B2(KEYINPUT87), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n640), .A2(new_n596), .B1(G264), .B2(new_n491), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(G190), .A3(new_n522), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n642), .A3(new_n584), .A4(new_n588), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n601), .A2(new_n628), .A3(new_n638), .A4(new_n643), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n479), .A2(new_n570), .A3(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n438), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT92), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n393), .B1(new_n390), .B2(new_n392), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n389), .A2(KEYINPUT92), .A3(new_n394), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n466), .A2(KEYINPUT71), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n469), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n460), .B1(new_n465), .B2(KEYINPUT71), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n316), .B1(new_n658), .B2(new_n321), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n653), .B1(new_n659), .B2(new_n377), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n646), .B1(new_n660), .B2(new_n435), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n492), .A2(new_n503), .A3(G179), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n436), .B1(new_n492), .B2(new_n503), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT89), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n514), .A2(new_n515), .ZN(new_n665));
  OAI22_X1  g0465(.A1(new_n665), .A2(new_n222), .B1(new_n202), .B2(new_n401), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n441), .B1(new_n327), .B2(new_n329), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n245), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n510), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n526), .A2(new_n671), .A3(new_n527), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n664), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(KEYINPUT90), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n664), .A2(new_n672), .A3(new_n676), .A4(new_n670), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n674), .A2(new_n675), .A3(new_n566), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n564), .A2(KEYINPUT88), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT88), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n556), .A2(new_n562), .A3(new_n680), .A4(new_n563), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n528), .A2(new_n555), .A3(new_n564), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(KEYINPUT26), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n678), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT91), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n678), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n670), .B1(new_n662), .B2(new_n663), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n568), .B1(new_n689), .B2(new_n567), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n567), .A2(new_n568), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n601), .A2(new_n638), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n692), .A2(new_n566), .A3(new_n693), .A4(new_n643), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n661), .B1(new_n479), .B2(new_n696), .ZN(G369));
  NAND3_X1  g0497(.A1(new_n258), .A2(new_n222), .A3(G13), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT27), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n699), .A2(G213), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n589), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n643), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n705), .A2(new_n601), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n601), .A2(new_n703), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n703), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n628), .B(new_n638), .C1(new_n611), .C2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n631), .B(new_n703), .C1(new_n635), .C2(new_n637), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n708), .A2(G330), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n638), .A2(new_n703), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n706), .A2(new_n715), .B1(new_n601), .B2(new_n703), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n713), .A2(new_n717), .ZN(G399));
  INV_X1    g0518(.A(new_n216), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G41), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n220), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n204), .A2(new_n365), .A3(new_n602), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT93), .ZN(new_n723));
  INV_X1    g0523(.A(new_n720), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(G1), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n721), .B1(new_n725), .B2(KEYINPUT94), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n726), .B1(KEYINPUT94), .B2(new_n725), .ZN(new_n727));
  XOR2_X1   g0527(.A(new_n727), .B(KEYINPUT28), .Z(new_n728));
  AOI21_X1  g0528(.A(new_n565), .B1(new_n673), .B2(KEYINPUT90), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(KEYINPUT98), .A3(KEYINPUT26), .A4(new_n677), .ZN(new_n730));
  INV_X1    g0530(.A(new_n682), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n694), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n674), .A2(KEYINPUT26), .A3(new_n566), .A4(new_n677), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT98), .B1(new_n683), .B2(new_n675), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n709), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n695), .A2(new_n709), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n737), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n522), .A2(new_n619), .A3(G179), .A4(new_n629), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(KEYINPUT95), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT95), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n612), .A2(new_n743), .A3(G179), .A4(new_n619), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n597), .A2(new_n598), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n746), .A2(new_n504), .A3(new_n541), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n745), .A2(KEYINPUT30), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g0548(.A(KEYINPUT96), .B(KEYINPUT30), .Z(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(new_n744), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n524), .A2(new_n525), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n534), .A2(new_n540), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n641), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n750), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n633), .A2(new_n541), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n756), .A2(new_n386), .A3(new_n504), .A4(new_n599), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n748), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  AND3_X1   g0558(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT31), .B1(new_n758), .B2(new_n703), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT97), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n504), .A2(new_n541), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n762), .A2(new_n742), .A3(new_n641), .A4(new_n744), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT30), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n749), .B1(new_n745), .B2(new_n747), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n703), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT31), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT97), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n703), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n644), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n690), .A2(new_n691), .A3(new_n565), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n773), .A2(new_n774), .A3(new_n709), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n761), .A2(new_n772), .A3(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n738), .A2(new_n740), .B1(G330), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n728), .B1(new_n777), .B2(G1), .ZN(G364));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n221), .B1(G20), .B2(new_n436), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n719), .A2(new_n326), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n239), .A2(G45), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT100), .Z(new_n787));
  AOI211_X1 g0587(.A(new_n785), .B(new_n787), .C1(new_n292), .C2(new_n220), .ZN(new_n788));
  INV_X1    g0588(.A(G355), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n326), .A2(new_n216), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n790), .B1(G116), .B2(new_n216), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n783), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n222), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(new_n317), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n328), .B1(new_n795), .B2(G107), .ZN(new_n796));
  NAND2_X1  g0596(.A1(G20), .A2(G179), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT101), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G190), .A2(G200), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n798), .A2(new_n369), .A3(new_n622), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n796), .B1(new_n800), .B2(new_n202), .C1(new_n331), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n793), .A2(new_n799), .ZN(new_n803));
  INV_X1    g0603(.A(G159), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT102), .B(KEYINPUT32), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n365), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n317), .A2(G179), .A3(G200), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n222), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n809), .B1(G97), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n798), .A2(new_n317), .A3(G200), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n807), .B(new_n813), .C1(new_n254), .C2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n798), .A2(new_n369), .A3(G200), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n802), .B(new_n815), .C1(G50), .C2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n812), .A2(G294), .B1(new_n795), .B2(G283), .ZN(new_n819));
  INV_X1    g0619(.A(new_n803), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n326), .B1(new_n820), .B2(G329), .ZN(new_n821));
  INV_X1    g0621(.A(G303), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n819), .B(new_n821), .C1(new_n822), .C2(new_n808), .ZN(new_n823));
  INV_X1    g0623(.A(G322), .ZN(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n801), .A2(new_n824), .B1(new_n800), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT103), .B(G326), .Z(new_n827));
  XOR2_X1   g0627(.A(KEYINPUT33), .B(G317), .Z(new_n828));
  OAI22_X1  g0628(.A1(new_n816), .A2(new_n827), .B1(new_n814), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g0629(.A1(new_n823), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n782), .B1(new_n818), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n222), .A2(G13), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n832), .A2(G45), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(G1), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n720), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n792), .A2(new_n831), .A3(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT104), .Z(new_n839));
  INV_X1    g0639(.A(new_n781), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n712), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n712), .A2(G330), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n712), .A2(G330), .ZN(new_n843));
  INV_X1    g0643(.A(new_n837), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n841), .B1(new_n842), .B2(new_n845), .ZN(G396));
  NAND3_X1  g0646(.A1(new_n695), .A2(new_n473), .A3(new_n709), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n529), .A2(new_n566), .A3(new_n569), .A4(new_n643), .ZN(new_n848));
  INV_X1    g0648(.A(new_n693), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(KEYINPUT91), .B2(new_n685), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n703), .B1(new_n851), .B2(new_n688), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n468), .A2(new_n703), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n655), .B2(new_n656), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n472), .B2(new_n853), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n847), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n776), .A2(G330), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n837), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n782), .A2(new_n779), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(G283), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n822), .A2(new_n816), .B1(new_n814), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(G294), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n801), .A2(new_n865), .B1(new_n800), .B2(new_n602), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n328), .B1(new_n803), .B2(new_n825), .C1(new_n811), .C2(new_n506), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n365), .A2(new_n794), .B1(new_n808), .B2(new_n441), .ZN(new_n868));
  NOR4_X1   g0668(.A1(new_n864), .A2(new_n866), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n801), .ZN(new_n870));
  INV_X1    g0670(.A(new_n800), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n870), .A2(G143), .B1(new_n871), .B2(G159), .ZN(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n872), .B1(new_n873), .B2(new_n816), .C1(new_n400), .C2(new_n814), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT34), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n795), .A2(G68), .ZN(new_n876));
  INV_X1    g0676(.A(G132), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n876), .B(new_n326), .C1(new_n877), .C2(new_n803), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n811), .A2(new_n331), .B1(new_n808), .B2(new_n406), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n869), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n782), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n837), .B1(G77), .B2(new_n862), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n855), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n779), .B2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT105), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n860), .A2(new_n886), .ZN(G384));
  OR2_X1    g0687(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(G116), .A3(new_n223), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT36), .Z(new_n891));
  OAI211_X1 g0691(.A(new_n220), .B(G77), .C1(new_n331), .C2(new_n254), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n406), .A2(G68), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n258), .B(G13), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n701), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n390), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT107), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n390), .A2(KEYINPUT107), .A3(new_n896), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n375), .B(KEYINPUT17), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n650), .A2(new_n651), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n390), .A2(new_n392), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n375), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n901), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n904), .A2(new_n375), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n899), .A4(new_n900), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n901), .A2(new_n903), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT108), .B1(new_n910), .B2(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n901), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n909), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT108), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n897), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT37), .B1(new_n905), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n909), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n918), .B1(new_n377), .B2(new_n395), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n920), .A2(KEYINPUT38), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n911), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT39), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n310), .A2(new_n312), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n927), .A2(new_n315), .A3(new_n304), .ZN(new_n928));
  INV_X1    g0728(.A(new_n277), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n930), .A2(new_n703), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT38), .B1(new_n920), .B2(new_n921), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n922), .A2(new_n932), .A3(new_n925), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n926), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n273), .A2(new_n276), .A3(new_n703), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT106), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n930), .A2(new_n938), .A3(new_n321), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n936), .B(KEYINPUT106), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n316), .B2(new_n322), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n657), .A2(new_n703), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n847), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n922), .A2(new_n932), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n653), .A2(new_n896), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n935), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n478), .A2(new_n740), .A3(new_n738), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n661), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT40), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n922), .B2(new_n932), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n775), .A2(new_n769), .A3(new_n771), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n957), .A2(new_n855), .A3(new_n939), .A4(new_n941), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n939), .A2(new_n941), .A3(new_n855), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n769), .A2(new_n771), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n570), .A2(new_n644), .A3(new_n703), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n924), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n959), .B1(new_n965), .B2(KEYINPUT40), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n479), .B2(new_n963), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n947), .A2(new_n964), .A3(new_n955), .ZN(new_n968));
  AOI21_X1  g0768(.A(KEYINPUT38), .B1(new_n912), .B2(new_n913), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n922), .B1(new_n969), .B2(new_n915), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n958), .B1(new_n970), .B2(new_n911), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n968), .B1(new_n971), .B2(new_n955), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n478), .A3(new_n957), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n967), .A2(G330), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n954), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n258), .B2(new_n832), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n954), .A2(new_n974), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n895), .B1(new_n976), .B2(new_n977), .ZN(G367));
  OAI211_X1 g0778(.A(new_n529), .B(new_n569), .C1(new_n519), .C2(new_n709), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n673), .A2(new_n709), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(new_n716), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT44), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n983), .B(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n717), .A2(KEYINPUT45), .A3(new_n981), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n982), .B2(new_n716), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n713), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(new_n713), .A3(new_n989), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT110), .B1(new_n712), .B2(G330), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n843), .B(KEYINPUT110), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n708), .B(new_n714), .ZN(new_n997));
  MUX2_X1   g0797(.A(new_n995), .B(new_n996), .S(new_n997), .Z(new_n998));
  NAND2_X1  g0798(.A1(new_n777), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n777), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n720), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n836), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n689), .B1(new_n982), .B2(new_n601), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n708), .A2(new_n981), .A3(new_n714), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n1006), .A2(new_n709), .B1(KEYINPUT42), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1007), .A2(KEYINPUT42), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n551), .A2(new_n553), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n703), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n731), .A2(KEYINPUT109), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n566), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT109), .B1(new_n731), .B2(new_n1012), .ZN(new_n1015));
  AND2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1016), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT43), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1010), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n713), .A2(new_n982), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1008), .A2(new_n1017), .A3(new_n1016), .A4(new_n1009), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1022), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1005), .A2(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n783), .B1(new_n216), .B2(new_n454), .C1(new_n234), .C2(new_n785), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1028), .A2(new_n837), .ZN(new_n1029));
  INV_X1    g0829(.A(G317), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n328), .B1(new_n803), .B2(new_n1030), .C1(new_n506), .C2(new_n794), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT112), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT111), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n808), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1034), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1032), .B1(new_n1033), .B2(new_n1035), .C1(new_n825), .C2(new_n816), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n870), .A2(G303), .B1(G107), .B2(new_n812), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n814), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1038), .A2(G294), .B1(new_n1035), .B2(new_n1033), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT46), .B1(new_n1034), .B2(G116), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G283), .B2(new_n871), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT113), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n808), .A2(new_n331), .B1(new_n803), .B2(new_n873), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1038), .A2(G159), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n817), .A2(G143), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n794), .A2(new_n202), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n328), .B(new_n1048), .C1(G68), .C2(new_n812), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n406), .B2(new_n800), .C1(new_n400), .C2(new_n801), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1036), .A2(new_n1042), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT47), .Z(new_n1052));
  OAI221_X1 g0852(.A(new_n1029), .B1(new_n882), .B2(new_n1052), .C1(new_n1019), .C2(new_n840), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1027), .A2(new_n1053), .ZN(G387));
  NAND2_X1  g0854(.A1(new_n998), .A2(new_n836), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n708), .A2(new_n840), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n801), .A2(new_n406), .B1(new_n800), .B2(new_n254), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n326), .B1(new_n803), .B2(new_n400), .C1(new_n506), .C2(new_n794), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n811), .A2(new_n454), .B1(new_n808), .B2(new_n202), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n1057), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n804), .B2(new_n816), .C1(new_n358), .C2(new_n814), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n827), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n326), .B1(new_n1062), .B2(new_n820), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n811), .A2(new_n863), .B1(new_n808), .B2(new_n865), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n870), .A2(G317), .B1(new_n871), .B2(G303), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n825), .B2(new_n814), .C1(new_n824), .C2(new_n816), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT49), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1063), .B1(new_n602), .B2(new_n794), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1061), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n782), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n784), .B1(new_n231), .B2(new_n292), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n450), .A2(G50), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT50), .ZN(new_n1077));
  AOI21_X1  g0877(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n723), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1075), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n723), .A2(new_n790), .B1(G107), .B2(new_n216), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT114), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n783), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1074), .A2(new_n837), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n999), .A2(new_n720), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n777), .A2(new_n998), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1055), .B1(new_n1056), .B2(new_n1084), .C1(new_n1085), .C2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(new_n993), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n713), .B1(new_n985), .B2(new_n989), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n982), .A2(new_n781), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n783), .B1(new_n506), .B2(new_n216), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n242), .B2(new_n784), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n328), .B1(new_n803), .B2(new_n824), .C1(new_n441), .C2(new_n794), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G283), .B2(new_n1034), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT115), .Z(new_n1096));
  AOI22_X1  g0896(.A1(new_n871), .A2(G294), .B1(G116), .B2(new_n812), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n822), .C2(new_n814), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n825), .A2(new_n801), .B1(new_n816), .B2(new_n1030), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  OAI22_X1  g0900(.A1(new_n400), .A2(new_n816), .B1(new_n801), .B2(new_n804), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT51), .Z(new_n1102));
  NAND2_X1  g0902(.A1(new_n812), .A2(G77), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n254), .B2(new_n808), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n328), .B1(new_n820), .B2(G143), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n365), .B2(new_n794), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n406), .B2(new_n814), .C1(new_n450), .C2(new_n800), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1098), .A2(new_n1100), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n844), .B(new_n1093), .C1(new_n1109), .C2(new_n782), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1090), .A2(new_n836), .B1(new_n1091), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n994), .A2(new_n999), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n720), .B1(new_n994), .B2(new_n999), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(G390));
  INV_X1    g0914(.A(new_n931), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n709), .B(new_n855), .C1(new_n732), .C2(new_n735), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1116), .A2(new_n945), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n924), .C1(new_n1117), .C2(new_n943), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n776), .A2(new_n942), .A3(G330), .A4(new_n855), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n847), .A2(new_n945), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n931), .B1(new_n1120), .B2(new_n942), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n933), .B1(new_n924), .B2(new_n925), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1118), .B(new_n1119), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(G330), .B1(new_n961), .B2(new_n962), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1125), .A2(new_n960), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n970), .B2(new_n911), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1128), .A2(new_n933), .B1(new_n946), .B2(new_n931), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n1129), .B2(new_n1118), .ZN(new_n1130));
  INV_X1    g0930(.A(G330), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n759), .A2(new_n760), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1132), .B2(new_n775), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n884), .B1(new_n1133), .B2(KEYINPUT117), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT117), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1125), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n942), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n776), .A2(G330), .A3(new_n855), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n943), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n1127), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(KEYINPUT116), .A3(new_n1120), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT116), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1126), .B1(new_n1140), .B2(new_n943), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n944), .B1(new_n852), .B2(new_n473), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1139), .B1(new_n1143), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n478), .A2(new_n1133), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n952), .A2(new_n661), .A3(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1124), .A2(new_n1130), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT116), .B1(new_n1142), .B2(new_n1120), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1145), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1118), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1126), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1150), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1155), .A2(new_n1157), .A3(new_n1123), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1151), .A2(new_n1159), .A3(new_n720), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n836), .A3(new_n1123), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n837), .B1(new_n357), .B2(new_n862), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n808), .A2(new_n400), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  INV_X1    g0964(.A(G128), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n816), .C1(new_n873), .C2(new_n814), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT54), .B(G143), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n870), .A2(G132), .B1(new_n871), .B2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n794), .A2(new_n406), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n328), .B(new_n1170), .C1(G125), .C2(new_n820), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n804), .C2(new_n811), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n870), .A2(G116), .B1(new_n871), .B2(G97), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n326), .B(new_n809), .C1(G294), .C2(new_n820), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1173), .A2(new_n1174), .A3(new_n876), .A4(new_n1103), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n863), .A2(new_n816), .B1(new_n814), .B2(new_n441), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1166), .A2(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1162), .B1(new_n1177), .B2(new_n782), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1122), .B2(new_n780), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1161), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1160), .A2(new_n1181), .ZN(G378));
  AOI21_X1  g0982(.A(new_n701), .B1(new_n424), .B2(new_n425), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n476), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n430), .A2(new_n434), .A3(new_n438), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1184), .A2(new_n1186), .A3(new_n1188), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n780), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n814), .A2(new_n877), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n812), .A2(G150), .B1(new_n1034), .B2(new_n1168), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n800), .B2(new_n873), .C1(new_n1165), .C2(new_n801), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G125), .C2(new_n817), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(KEYINPUT59), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n795), .A2(G159), .ZN(new_n1201));
  AOI211_X1 g1001(.A(G33), .B(G41), .C1(new_n820), .C2(G124), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n870), .A2(G107), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1204), .B(KEYINPUT119), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n331), .A2(new_n794), .B1(new_n808), .B2(new_n202), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n326), .A2(G41), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n863), .B2(new_n803), .C1(new_n254), .C2(new_n811), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1206), .B(new_n1208), .C1(new_n455), .C2(new_n871), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(G116), .A2(new_n817), .B1(new_n1038), .B2(G97), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1205), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G50), .B(new_n1207), .C1(new_n247), .C2(new_n291), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT118), .ZN(new_n1216));
  AND4_X1   g1016(.A1(new_n1203), .A2(new_n1213), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n837), .B1(G50), .B2(new_n862), .C1(new_n1217), .C2(new_n882), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1193), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT121), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n951), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1192), .B1(new_n972), .B2(G330), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n955), .B1(new_n924), .B2(new_n964), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G330), .B(new_n1192), .C1(new_n1224), .C2(new_n959), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1222), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1192), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n966), .B2(new_n1131), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1229), .A2(new_n1221), .A3(new_n951), .A4(new_n1225), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1220), .B1(new_n1231), .B2(new_n1004), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n951), .B1(new_n1226), .B2(new_n1223), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n949), .B1(new_n1122), .B2(new_n931), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1229), .A2(new_n948), .A3(new_n1235), .A4(new_n1225), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT122), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1150), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n952), .A2(new_n1149), .A3(KEYINPUT122), .A4(new_n661), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1159), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n724), .B1(new_n1237), .B2(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1150), .B1(new_n1246), .B2(new_n1152), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1241), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1233), .B1(new_n1248), .B2(new_n1231), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1232), .B1(new_n1244), .B2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(G375));
  OAI21_X1  g1051(.A(new_n837), .B1(G68), .B2(new_n862), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n326), .B1(new_n803), .B2(new_n1165), .C1(new_n331), .C2(new_n794), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n811), .A2(new_n406), .B1(new_n808), .B2(new_n804), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n873), .B2(new_n801), .C1(new_n400), .C2(new_n800), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n877), .A2(new_n816), .B1(new_n814), .B2(new_n1167), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n870), .A2(G283), .B1(new_n871), .B2(G107), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n326), .B(new_n1048), .C1(G303), .C2(new_n820), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n812), .A2(new_n455), .B1(new_n1034), .B2(G97), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n865), .A2(new_n816), .B1(new_n814), .B2(new_n602), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1256), .A2(new_n1257), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1252), .B1(new_n1263), .B2(new_n782), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n942), .B2(new_n780), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1148), .B2(new_n1004), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT123), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(KEYINPUT123), .B(new_n1265), .C1(new_n1148), .C2(new_n1004), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1246), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1002), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(G381));
  OR4_X1    g1074(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1275), .A2(G381), .A3(G387), .A4(G378), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1250), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1277), .B(KEYINPUT124), .Z(G407));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(G378), .A2(G343), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1279), .B1(new_n1250), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G407), .A2(new_n1281), .ZN(G409));
  AND2_X1   g1082(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1002), .A3(new_n1243), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1219), .B1(new_n1285), .B2(new_n836), .ZN(new_n1286));
  AOI21_X1  g1086(.A(G378), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(G378), .B2(new_n1250), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1279), .A2(G343), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT125), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1232), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT57), .B1(new_n1283), .B2(new_n1243), .ZN(new_n1292));
  NOR3_X1   g1092(.A1(new_n1226), .A2(new_n1223), .A3(new_n951), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1229), .A2(new_n1225), .B1(new_n948), .B2(new_n1235), .ZN(new_n1294));
  OAI21_X1  g1094(.A(KEYINPUT57), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n720), .B1(new_n1295), .B2(new_n1248), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G378), .B(new_n1291), .C1(new_n1292), .C2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1157), .A2(new_n1123), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n724), .B1(new_n1271), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1180), .B1(new_n1300), .B2(new_n1159), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1289), .B1(new_n1297), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1289), .A2(G2897), .ZN(new_n1306));
  XOR2_X1   g1106(.A(new_n1306), .B(KEYINPUT126), .Z(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1272), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1148), .A2(KEYINPUT60), .A3(new_n1150), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1271), .A4(new_n720), .ZN(new_n1312));
  AND3_X1   g1112(.A1(new_n1270), .A2(G384), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G384), .B1(new_n1270), .B2(new_n1312), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1308), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1270), .A2(new_n1312), .ZN(new_n1316));
  INV_X1    g1116(.A(G384), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1270), .A2(G384), .A3(new_n1312), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(new_n1319), .A3(new_n1307), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1315), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1290), .A2(new_n1305), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT127), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G390), .B1(new_n1027), .B2(new_n1053), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n836), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1026), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G390), .B(new_n1053), .C1(new_n1326), .C2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1324), .B1(new_n1325), .B2(new_n1329), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(G393), .B(G396), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT61), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1324), .B(new_n1331), .C1(new_n1325), .C2(new_n1329), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1289), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1338));
  AOI211_X1 g1138(.A(new_n1232), .B(new_n1301), .C1(new_n1249), .C2(new_n1244), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1337), .B(new_n1338), .C1(new_n1339), .C2(new_n1287), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1336), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1338), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1323), .A2(new_n1342), .A3(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1303), .A2(new_n1345), .A3(new_n1338), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1334), .B1(new_n1303), .B2(new_n1321), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1345), .B1(new_n1303), .B2(new_n1338), .ZN(new_n1348));
  NOR3_X1   g1148(.A1(new_n1346), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1344), .B1(new_n1349), .B2(new_n1351), .ZN(G405));
  NOR2_X1   g1152(.A1(new_n1250), .A2(G378), .ZN(new_n1353));
  OR3_X1    g1153(.A1(new_n1339), .A2(new_n1353), .A3(new_n1338), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1338), .B1(new_n1339), .B2(new_n1353), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1350), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1354), .A2(new_n1351), .A3(new_n1355), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(G402));
endmodule


