

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XNOR2_X1 U322 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U323 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U324 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n407) );
  XNOR2_X1 U325 ( .A(n408), .B(n407), .ZN(n566) );
  XNOR2_X1 U326 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n323) );
  XNOR2_X1 U327 ( .A(n458), .B(n323), .ZN(n548) );
  XNOR2_X1 U328 ( .A(n451), .B(KEYINPUT58), .ZN(n452) );
  XNOR2_X1 U329 ( .A(n453), .B(n452), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n291) );
  NAND2_X1 U331 ( .A1(G227GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U333 ( .A(n292), .B(G176GAT), .Z(n300) );
  XOR2_X1 U334 ( .A(KEYINPUT17), .B(G183GAT), .Z(n294) );
  XNOR2_X1 U335 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U337 ( .A(KEYINPUT83), .B(n295), .Z(n393) );
  XOR2_X1 U338 ( .A(G99GAT), .B(G15GAT), .Z(n297) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(G43GAT), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n393), .B(n298), .ZN(n299) );
  XNOR2_X1 U342 ( .A(n300), .B(n299), .ZN(n303) );
  XOR2_X1 U343 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n302) );
  XNOR2_X1 U344 ( .A(G113GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n423) );
  XOR2_X1 U346 ( .A(n303), .B(n423), .Z(n305) );
  XOR2_X1 U347 ( .A(G190GAT), .B(G134GAT), .Z(n350) );
  XOR2_X1 U348 ( .A(G120GAT), .B(G71GAT), .Z(n307) );
  XNOR2_X1 U349 ( .A(n350), .B(n307), .ZN(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n526) );
  XNOR2_X1 U351 ( .A(G106GAT), .B(G78GAT), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n306), .B(G148GAT), .ZN(n433) );
  XOR2_X1 U353 ( .A(KEYINPUT13), .B(G57GAT), .Z(n363) );
  XNOR2_X1 U354 ( .A(n307), .B(n363), .ZN(n309) );
  XOR2_X1 U355 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n308) );
  XNOR2_X1 U356 ( .A(n309), .B(n308), .ZN(n315) );
  XOR2_X1 U357 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n311) );
  XNOR2_X1 U358 ( .A(KEYINPUT31), .B(KEYINPUT75), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n311), .B(n310), .ZN(n313) );
  AND2_X1 U360 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  XOR2_X1 U361 ( .A(n433), .B(n316), .Z(n322) );
  XOR2_X1 U362 ( .A(G92GAT), .B(G64GAT), .Z(n318) );
  XNOR2_X1 U363 ( .A(G176GAT), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U365 ( .A(KEYINPUT74), .B(n319), .Z(n392) );
  XNOR2_X1 U366 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n320), .B(KEYINPUT73), .ZN(n355) );
  XNOR2_X1 U368 ( .A(n392), .B(n355), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n458) );
  XNOR2_X1 U370 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n324) );
  XNOR2_X1 U371 ( .A(n324), .B(G29GAT), .ZN(n325) );
  XOR2_X1 U372 ( .A(n325), .B(KEYINPUT7), .Z(n327) );
  XNOR2_X1 U373 ( .A(G43GAT), .B(G50GAT), .ZN(n326) );
  XNOR2_X1 U374 ( .A(n327), .B(n326), .ZN(n346) );
  XOR2_X1 U375 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n329) );
  XNOR2_X1 U376 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n331) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(G22GAT), .ZN(n431) );
  INV_X1 U379 ( .A(n431), .ZN(n330) );
  XNOR2_X1 U380 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U381 ( .A(G169GAT), .B(G8GAT), .Z(n397) );
  XOR2_X1 U382 ( .A(n397), .B(G197GAT), .Z(n333) );
  NAND2_X1 U383 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U385 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U386 ( .A(G15GAT), .B(G1GAT), .Z(n375) );
  XOR2_X1 U387 ( .A(n336), .B(n375), .Z(n338) );
  XNOR2_X1 U388 ( .A(KEYINPUT68), .B(G113GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n346), .B(n339), .ZN(n570) );
  NAND2_X1 U391 ( .A1(n548), .A2(n570), .ZN(n342) );
  XOR2_X1 U392 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n340) );
  XNOR2_X1 U393 ( .A(KEYINPUT112), .B(n340), .ZN(n341) );
  XNOR2_X1 U394 ( .A(n342), .B(n341), .ZN(n381) );
  XOR2_X1 U395 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n344) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(KEYINPUT66), .ZN(n343) );
  XNOR2_X1 U397 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U399 ( .A(G162GAT), .B(KEYINPUT9), .Z(n348) );
  XNOR2_X1 U400 ( .A(G92GAT), .B(G218GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n352) );
  AND2_X1 U403 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U404 ( .A(n352), .B(n351), .ZN(n354) );
  INV_X1 U405 ( .A(KEYINPUT76), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n357) );
  XNOR2_X1 U407 ( .A(n355), .B(KEYINPUT65), .ZN(n356) );
  XNOR2_X1 U408 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U409 ( .A(n359), .B(n358), .ZN(n555) );
  XOR2_X1 U410 ( .A(KEYINPUT78), .B(G78GAT), .Z(n361) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G64GAT), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U413 ( .A(n363), .B(n362), .Z(n365) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G8GAT), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n365), .B(n364), .ZN(n379) );
  XOR2_X1 U416 ( .A(KEYINPUT79), .B(G211GAT), .Z(n367) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U419 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n369) );
  XNOR2_X1 U420 ( .A(G127GAT), .B(G155GAT), .ZN(n368) );
  XNOR2_X1 U421 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U422 ( .A(n371), .B(n370), .Z(n377) );
  XOR2_X1 U423 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n373) );
  XNOR2_X1 U424 ( .A(G183GAT), .B(KEYINPUT77), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U427 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U428 ( .A(n379), .B(n378), .ZN(n561) );
  INV_X1 U429 ( .A(n561), .ZN(n578) );
  NOR2_X1 U430 ( .A1(n555), .A2(n578), .ZN(n380) );
  AND2_X1 U431 ( .A1(n381), .A2(n380), .ZN(n382) );
  XNOR2_X1 U432 ( .A(n382), .B(KEYINPUT47), .ZN(n389) );
  XNOR2_X1 U433 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n383) );
  INV_X1 U434 ( .A(n555), .ZN(n541) );
  XNOR2_X1 U435 ( .A(n383), .B(n541), .ZN(n583) );
  NOR2_X1 U436 ( .A1(n583), .A2(n561), .ZN(n384) );
  XNOR2_X1 U437 ( .A(KEYINPUT45), .B(n384), .ZN(n385) );
  NAND2_X1 U438 ( .A1(n385), .A2(n458), .ZN(n386) );
  XOR2_X1 U439 ( .A(KEYINPUT114), .B(n386), .Z(n387) );
  INV_X1 U440 ( .A(n570), .ZN(n545) );
  XNOR2_X1 U441 ( .A(n545), .B(KEYINPUT70), .ZN(n558) );
  NAND2_X1 U442 ( .A1(n387), .A2(n558), .ZN(n388) );
  NAND2_X1 U443 ( .A1(n389), .A2(n388), .ZN(n391) );
  XOR2_X1 U444 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n390) );
  XNOR2_X1 U445 ( .A(n391), .B(n390), .ZN(n527) );
  XNOR2_X1 U446 ( .A(n393), .B(n392), .ZN(n406) );
  XOR2_X1 U447 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n395) );
  XNOR2_X1 U448 ( .A(G36GAT), .B(G190GAT), .ZN(n394) );
  XNOR2_X1 U449 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U450 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U451 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n402) );
  XOR2_X1 U453 ( .A(KEYINPUT21), .B(G211GAT), .Z(n401) );
  XNOR2_X1 U454 ( .A(G197GAT), .B(G218GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n441) );
  XOR2_X1 U456 ( .A(n402), .B(n441), .Z(n404) );
  XNOR2_X1 U457 ( .A(KEYINPUT92), .B(KEYINPUT94), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U459 ( .A(n406), .B(n405), .ZN(n466) );
  NAND2_X1 U460 ( .A1(n527), .A2(n466), .ZN(n408) );
  XOR2_X1 U461 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n410) );
  XNOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n416) );
  XOR2_X1 U464 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n412) );
  XNOR2_X1 U465 ( .A(G162GAT), .B(G155GAT), .ZN(n411) );
  XNOR2_X1 U466 ( .A(n412), .B(n411), .ZN(n440) );
  XOR2_X1 U467 ( .A(n440), .B(KEYINPUT6), .Z(n414) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n430) );
  XOR2_X1 U471 ( .A(G57GAT), .B(G148GAT), .Z(n418) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G120GAT), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n420) );
  XNOR2_X1 U475 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U477 ( .A(n422), .B(n421), .Z(n428) );
  XOR2_X1 U478 ( .A(G85GAT), .B(n423), .Z(n425) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(G134GAT), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U481 ( .A(G141GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n565) );
  XNOR2_X1 U484 ( .A(G50GAT), .B(G204GAT), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n445) );
  XOR2_X1 U486 ( .A(KEYINPUT85), .B(n433), .Z(n435) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U489 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n437) );
  XNOR2_X1 U490 ( .A(KEYINPUT86), .B(KEYINPUT22), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U492 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n468) );
  INV_X1 U496 ( .A(n468), .ZN(n446) );
  AND2_X1 U497 ( .A1(n565), .A2(n446), .ZN(n447) );
  AND2_X1 U498 ( .A1(n566), .A2(n447), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n448), .B(KEYINPUT55), .ZN(n449) );
  NOR2_X1 U500 ( .A1(n526), .A2(n449), .ZN(n450) );
  XOR2_X1 U501 ( .A(KEYINPUT122), .B(n450), .Z(n562) );
  NOR2_X1 U502 ( .A1(n562), .A2(n541), .ZN(n453) );
  INV_X1 U503 ( .A(G190GAT), .ZN(n451) );
  XOR2_X1 U504 ( .A(n548), .B(KEYINPUT106), .Z(n533) );
  NOR2_X1 U505 ( .A1(n562), .A2(n533), .ZN(n457) );
  XNOR2_X1 U506 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n455) );
  XNOR2_X1 U507 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  INV_X1 U510 ( .A(n458), .ZN(n575) );
  NOR2_X1 U511 ( .A1(n558), .A2(n575), .ZN(n490) );
  NAND2_X1 U512 ( .A1(n541), .A2(n578), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(KEYINPUT81), .ZN(n460) );
  XNOR2_X1 U514 ( .A(KEYINPUT16), .B(n460), .ZN(n474) );
  XNOR2_X1 U515 ( .A(n468), .B(KEYINPUT28), .ZN(n525) );
  XNOR2_X1 U516 ( .A(n466), .B(KEYINPUT27), .ZN(n528) );
  NAND2_X1 U517 ( .A1(n526), .A2(n528), .ZN(n461) );
  NOR2_X1 U518 ( .A1(n525), .A2(n461), .ZN(n462) );
  NOR2_X1 U519 ( .A1(n565), .A2(n462), .ZN(n473) );
  NAND2_X1 U520 ( .A1(n468), .A2(n526), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT96), .ZN(n464) );
  XOR2_X1 U522 ( .A(KEYINPUT26), .B(n464), .Z(n567) );
  NAND2_X1 U523 ( .A1(n567), .A2(n528), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n565), .A2(n465), .ZN(n471) );
  INV_X1 U525 ( .A(n466), .ZN(n515) );
  NOR2_X1 U526 ( .A1(n526), .A2(n515), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U528 ( .A(KEYINPUT25), .B(n469), .Z(n470) );
  NOR2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n488) );
  AND2_X1 U531 ( .A1(n474), .A2(n488), .ZN(n501) );
  NAND2_X1 U532 ( .A1(n490), .A2(n501), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT97), .B(n475), .Z(n484) );
  NOR2_X1 U534 ( .A1(n565), .A2(n484), .ZN(n476) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n476), .Z(n477) );
  XNOR2_X1 U536 ( .A(KEYINPUT34), .B(n477), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n515), .A2(n484), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT98), .B(n478), .Z(n479) );
  XNOR2_X1 U539 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n484), .A2(n526), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n481) );
  XNOR2_X1 U542 ( .A(G15GAT), .B(KEYINPUT100), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  INV_X1 U545 ( .A(n525), .ZN(n521) );
  NOR2_X1 U546 ( .A1(n521), .A2(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(G1327GAT) );
  NOR2_X1 U549 ( .A1(n578), .A2(n583), .ZN(n487) );
  NAND2_X1 U550 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT37), .B(n489), .ZN(n510) );
  NAND2_X1 U552 ( .A1(n510), .A2(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT103), .Z(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n498) );
  NOR2_X1 U555 ( .A1(n565), .A2(n498), .ZN(n493) );
  XNOR2_X1 U556 ( .A(n493), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n498), .A2(n515), .ZN(n495) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  NOR2_X1 U560 ( .A1(n526), .A2(n498), .ZN(n496) );
  XOR2_X1 U561 ( .A(KEYINPUT40), .B(n496), .Z(n497) );
  XNOR2_X1 U562 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NOR2_X1 U563 ( .A1(n521), .A2(n498), .ZN(n499) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n499), .Z(n500) );
  XNOR2_X1 U565 ( .A(KEYINPUT104), .B(n500), .ZN(G1331GAT) );
  NOR2_X1 U566 ( .A1(n533), .A2(n570), .ZN(n511) );
  NAND2_X1 U567 ( .A1(n511), .A2(n501), .ZN(n507) );
  NOR2_X1 U568 ( .A1(n565), .A2(n507), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n515), .A2(n507), .ZN(n505) );
  XOR2_X1 U573 ( .A(G64GAT), .B(n505), .Z(G1333GAT) );
  NOR2_X1 U574 ( .A1(n526), .A2(n507), .ZN(n506) );
  XOR2_X1 U575 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U576 ( .A1(n521), .A2(n507), .ZN(n509) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n509), .B(n508), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n511), .A2(n510), .ZN(n512) );
  XOR2_X1 U580 ( .A(KEYINPUT107), .B(n512), .Z(n520) );
  NOR2_X1 U581 ( .A1(n565), .A2(n520), .ZN(n513) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n513), .Z(n514) );
  XNOR2_X1 U583 ( .A(KEYINPUT108), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U584 ( .A1(n515), .A2(n520), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n526), .A2(n520), .ZN(n518) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(n518), .Z(n519) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n519), .ZN(G1338GAT) );
  NOR2_X1 U590 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n522) );
  XNOR2_X1 U592 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n531) );
  NAND2_X1 U595 ( .A1(n527), .A2(n528), .ZN(n529) );
  NOR2_X1 U596 ( .A1(n565), .A2(n529), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT116), .B(n530), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n531), .A2(n544), .ZN(n540) );
  NOR2_X1 U599 ( .A1(n558), .A2(n540), .ZN(n532) );
  XOR2_X1 U600 ( .A(G113GAT), .B(n532), .Z(G1340GAT) );
  NOR2_X1 U601 ( .A1(n533), .A2(n540), .ZN(n535) );
  XNOR2_X1 U602 ( .A(KEYINPUT117), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U603 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  NOR2_X1 U605 ( .A1(n561), .A2(n540), .ZN(n538) );
  XNOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n539), .Z(G1342GAT) );
  NOR2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n542) );
  XNOR2_X1 U611 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n567), .A2(n544), .ZN(n547) );
  NOR2_X1 U613 ( .A1(n545), .A2(n547), .ZN(n546) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n546), .Z(G1344GAT) );
  XOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT119), .Z(n550) );
  INV_X1 U616 ( .A(n547), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n556), .A2(n548), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U619 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n578), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n558), .A2(n562), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(KEYINPUT123), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(KEYINPUT126), .B(KEYINPUT59), .ZN(n574) );
  XOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .Z(n572) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n569) );
  INV_X1 U635 ( .A(n567), .ZN(n568) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n581) );
  NAND2_X1 U637 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  XOR2_X1 U643 ( .A(G211GAT), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1354GAT) );
  INV_X1 U646 ( .A(n581), .ZN(n582) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U648 ( .A(KEYINPUT62), .B(n584), .Z(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

