

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575;

  NOR2_X1 U317 ( .A1(n462), .A2(n573), .ZN(n463) );
  XNOR2_X1 U318 ( .A(n434), .B(n433), .ZN(n437) );
  XOR2_X1 U319 ( .A(n324), .B(n323), .Z(n505) );
  XOR2_X1 U320 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n285) );
  INV_X1 U321 ( .A(G176GAT), .ZN(n431) );
  XNOR2_X1 U322 ( .A(n432), .B(n431), .ZN(n434) );
  XNOR2_X1 U323 ( .A(n402), .B(KEYINPUT119), .ZN(n403) );
  XNOR2_X1 U324 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U325 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n452) );
  XNOR2_X1 U326 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U327 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U328 ( .A(n453), .B(n452), .ZN(n556) );
  XNOR2_X1 U329 ( .A(n423), .B(n422), .ZN(n442) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n443) );
  XOR2_X1 U331 ( .A(n340), .B(n339), .Z(n535) );
  XNOR2_X1 U332 ( .A(n441), .B(n440), .ZN(n515) );
  XNOR2_X1 U333 ( .A(n443), .B(KEYINPUT58), .ZN(n444) );
  XNOR2_X1 U334 ( .A(n468), .B(G43GAT), .ZN(n469) );
  XNOR2_X1 U335 ( .A(n445), .B(n444), .ZN(G1351GAT) );
  XNOR2_X1 U336 ( .A(n470), .B(n469), .ZN(G1330GAT) );
  XOR2_X1 U337 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n287) );
  XNOR2_X1 U338 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n286) );
  XNOR2_X1 U339 ( .A(n287), .B(n286), .ZN(n305) );
  XOR2_X1 U340 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n289) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(KEYINPUT75), .ZN(n288) );
  XNOR2_X1 U342 ( .A(n289), .B(n288), .ZN(n291) );
  INV_X1 U343 ( .A(G218GAT), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n293) );
  XOR2_X1 U345 ( .A(G43GAT), .B(G134GAT), .Z(n435) );
  XNOR2_X1 U346 ( .A(G190GAT), .B(n435), .ZN(n292) );
  XNOR2_X1 U347 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U348 ( .A(G85GAT), .B(G92GAT), .Z(n370) );
  XOR2_X1 U349 ( .A(n370), .B(KEYINPUT77), .Z(n295) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U352 ( .A(n297), .B(n296), .Z(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT67), .B(KEYINPUT7), .Z(n299) );
  XNOR2_X1 U354 ( .A(G36GAT), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U356 ( .A(KEYINPUT8), .B(n300), .ZN(n339) );
  INV_X1 U357 ( .A(n339), .ZN(n301) );
  XOR2_X1 U358 ( .A(G50GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U359 ( .A(n301), .B(n409), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U361 ( .A(n305), .B(n304), .Z(n471) );
  XOR2_X1 U362 ( .A(G127GAT), .B(KEYINPUT0), .Z(n307) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n427) );
  XOR2_X1 U365 ( .A(n427), .B(G1GAT), .Z(n309) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n324) );
  XOR2_X1 U368 ( .A(G85GAT), .B(G162GAT), .Z(n311) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(G134GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U371 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n313) );
  XNOR2_X1 U372 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U374 ( .A(n315), .B(n314), .Z(n322) );
  XOR2_X1 U375 ( .A(G155GAT), .B(KEYINPUT2), .Z(n317) );
  XNOR2_X1 U376 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n316) );
  XNOR2_X1 U377 ( .A(n317), .B(n316), .ZN(n416) );
  XOR2_X1 U378 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n319) );
  XNOR2_X1 U379 ( .A(G120GAT), .B(G148GAT), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n416), .B(n320), .ZN(n321) );
  XNOR2_X1 U382 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U383 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n326) );
  XNOR2_X1 U384 ( .A(G197GAT), .B(G141GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n338) );
  XOR2_X1 U386 ( .A(G43GAT), .B(G50GAT), .Z(n330) );
  XOR2_X1 U387 ( .A(G8GAT), .B(G1GAT), .Z(n328) );
  XNOR2_X1 U388 ( .A(G15GAT), .B(G22GAT), .ZN(n327) );
  XNOR2_X1 U389 ( .A(n328), .B(n327), .ZN(n341) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(n341), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n332) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XOR2_X1 U394 ( .A(n332), .B(n331), .Z(n334) );
  XNOR2_X1 U395 ( .A(G169GAT), .B(KEYINPUT69), .ZN(n333) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U397 ( .A(n341), .B(KEYINPUT79), .Z(n343) );
  NAND2_X1 U398 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n358) );
  XOR2_X1 U400 ( .A(G211GAT), .B(G127GAT), .Z(n345) );
  XNOR2_X1 U401 ( .A(G183GAT), .B(G71GAT), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n348) );
  XOR2_X1 U403 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n347) );
  XNOR2_X1 U404 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n361) );
  XOR2_X1 U406 ( .A(n348), .B(n361), .Z(n356) );
  XOR2_X1 U407 ( .A(KEYINPUT15), .B(G64GAT), .Z(n350) );
  XNOR2_X1 U408 ( .A(G155GAT), .B(G78GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U410 ( .A(KEYINPUT78), .B(KEYINPUT12), .Z(n352) );
  XNOR2_X1 U411 ( .A(KEYINPUT80), .B(KEYINPUT14), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U414 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U415 ( .A(n358), .B(n357), .Z(n568) );
  XNOR2_X1 U416 ( .A(n471), .B(KEYINPUT36), .ZN(n573) );
  NOR2_X1 U417 ( .A1(n568), .A2(n573), .ZN(n359) );
  XNOR2_X1 U418 ( .A(KEYINPUT45), .B(n359), .ZN(n375) );
  XNOR2_X1 U419 ( .A(G176GAT), .B(G204GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n360), .B(G64GAT), .ZN(n394) );
  XOR2_X1 U421 ( .A(n361), .B(n394), .Z(n366) );
  XNOR2_X1 U422 ( .A(G99GAT), .B(G71GAT), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n362), .B(G120GAT), .ZN(n428) );
  XOR2_X1 U424 ( .A(G78GAT), .B(G148GAT), .Z(n364) );
  XNOR2_X1 U425 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n363) );
  XNOR2_X1 U426 ( .A(n364), .B(n363), .ZN(n414) );
  XNOR2_X1 U427 ( .A(n428), .B(n414), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n374) );
  XOR2_X1 U429 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n368) );
  XNOR2_X1 U430 ( .A(KEYINPUT73), .B(KEYINPUT32), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U432 ( .A(n370), .B(n369), .Z(n372) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U435 ( .A(n374), .B(n373), .Z(n563) );
  NAND2_X1 U436 ( .A1(n375), .A2(n563), .ZN(n376) );
  NOR2_X1 U437 ( .A1(n535), .A2(n376), .ZN(n377) );
  XNOR2_X1 U438 ( .A(KEYINPUT111), .B(n377), .ZN(n384) );
  XOR2_X1 U439 ( .A(KEYINPUT110), .B(KEYINPUT47), .Z(n382) );
  INV_X1 U440 ( .A(n568), .ZN(n541) );
  INV_X1 U441 ( .A(n563), .ZN(n464) );
  XOR2_X1 U442 ( .A(KEYINPUT41), .B(n464), .Z(n537) );
  INV_X1 U443 ( .A(n537), .ZN(n551) );
  INV_X1 U444 ( .A(n535), .ZN(n558) );
  NOR2_X1 U445 ( .A1(n551), .A2(n558), .ZN(n378) );
  XNOR2_X1 U446 ( .A(n378), .B(KEYINPUT46), .ZN(n379) );
  NOR2_X1 U447 ( .A1(n541), .A2(n379), .ZN(n380) );
  NAND2_X1 U448 ( .A1(n380), .A2(n471), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n383) );
  NAND2_X1 U450 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n385), .B(KEYINPUT48), .ZN(n532) );
  XOR2_X1 U452 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n387) );
  XNOR2_X1 U453 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n386) );
  XNOR2_X1 U454 ( .A(n387), .B(n386), .ZN(n389) );
  INV_X1 U455 ( .A(KEYINPUT18), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U457 ( .A(G169GAT), .B(G183GAT), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n439) );
  XOR2_X1 U459 ( .A(G92GAT), .B(G8GAT), .Z(n393) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n395) );
  XOR2_X1 U462 ( .A(n395), .B(n394), .Z(n400) );
  XOR2_X1 U463 ( .A(KEYINPUT90), .B(G218GAT), .Z(n397) );
  XNOR2_X1 U464 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U466 ( .A(G197GAT), .B(n398), .Z(n417) );
  XNOR2_X1 U467 ( .A(G36GAT), .B(n417), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n439), .B(n401), .ZN(n508) );
  NAND2_X1 U470 ( .A1(n532), .A2(n508), .ZN(n404) );
  XOR2_X1 U471 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n402) );
  NOR2_X1 U472 ( .A1(n505), .A2(n405), .ZN(n557) );
  XOR2_X1 U473 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n407) );
  XNOR2_X1 U474 ( .A(G22GAT), .B(KEYINPUT92), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U476 ( .A(n409), .B(n408), .Z(n411) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U478 ( .A(n411), .B(n410), .ZN(n421) );
  XOR2_X1 U479 ( .A(G204GAT), .B(KEYINPUT23), .Z(n413) );
  XNOR2_X1 U480 ( .A(KEYINPUT89), .B(KEYINPUT91), .ZN(n412) );
  XNOR2_X1 U481 ( .A(n413), .B(n412), .ZN(n415) );
  XOR2_X1 U482 ( .A(n415), .B(n414), .Z(n419) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n451) );
  NAND2_X1 U486 ( .A1(n557), .A2(n451), .ZN(n423) );
  XOR2_X1 U487 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n422) );
  XOR2_X1 U488 ( .A(KEYINPUT87), .B(KEYINPUT84), .Z(n425) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U491 ( .A(n426), .B(KEYINPUT83), .Z(n430) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n441) );
  XNOR2_X1 U494 ( .A(KEYINPUT85), .B(KEYINPUT64), .ZN(n432) );
  XOR2_X1 U495 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n433) );
  XNOR2_X1 U496 ( .A(G15GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n440) );
  NAND2_X1 U499 ( .A1(n442), .A2(n515), .ZN(n554) );
  NOR2_X1 U500 ( .A1(n471), .A2(n554), .ZN(n445) );
  XOR2_X1 U501 ( .A(KEYINPUT38), .B(KEYINPUT104), .Z(n467) );
  XNOR2_X1 U502 ( .A(n515), .B(KEYINPUT88), .ZN(n448) );
  XNOR2_X1 U503 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n446) );
  XNOR2_X1 U504 ( .A(n446), .B(n508), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n505), .A2(n454), .ZN(n534) );
  XOR2_X1 U506 ( .A(KEYINPUT28), .B(n451), .Z(n512) );
  NOR2_X1 U507 ( .A1(n534), .A2(n512), .ZN(n516) );
  XNOR2_X1 U508 ( .A(n516), .B(KEYINPUT95), .ZN(n447) );
  NOR2_X1 U509 ( .A1(n448), .A2(n447), .ZN(n460) );
  NAND2_X1 U510 ( .A1(n515), .A2(n508), .ZN(n449) );
  NAND2_X1 U511 ( .A1(n451), .A2(n449), .ZN(n450) );
  XNOR2_X1 U512 ( .A(n450), .B(KEYINPUT25), .ZN(n456) );
  NOR2_X1 U513 ( .A1(n515), .A2(n451), .ZN(n453) );
  AND2_X1 U514 ( .A1(n556), .A2(n454), .ZN(n455) );
  NOR2_X1 U515 ( .A1(n456), .A2(n455), .ZN(n457) );
  OR2_X1 U516 ( .A1(n505), .A2(n457), .ZN(n458) );
  XNOR2_X1 U517 ( .A(KEYINPUT97), .B(n458), .ZN(n459) );
  NOR2_X1 U518 ( .A1(n460), .A2(n459), .ZN(n474) );
  NOR2_X1 U519 ( .A1(n474), .A2(n541), .ZN(n461) );
  XOR2_X1 U520 ( .A(KEYINPUT102), .B(n461), .Z(n462) );
  XNOR2_X1 U521 ( .A(n463), .B(n285), .ZN(n503) );
  NOR2_X1 U522 ( .A1(n464), .A2(n558), .ZN(n465) );
  XOR2_X1 U523 ( .A(n465), .B(KEYINPUT74), .Z(n476) );
  OR2_X1 U524 ( .A1(n503), .A2(n476), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n467), .B(n466), .ZN(n490) );
  NAND2_X1 U526 ( .A1(n490), .A2(n515), .ZN(n470) );
  XOR2_X1 U527 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n468) );
  INV_X1 U528 ( .A(n471), .ZN(n545) );
  NOR2_X1 U529 ( .A1(n568), .A2(n545), .ZN(n472) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n472), .Z(n473) );
  NOR2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(n475), .Z(n493) );
  NOR2_X1 U533 ( .A1(n476), .A2(n493), .ZN(n483) );
  NAND2_X1 U534 ( .A1(n505), .A2(n483), .ZN(n477) );
  XNOR2_X1 U535 ( .A(KEYINPUT34), .B(n477), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U537 ( .A1(n508), .A2(n483), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U540 ( .A1(n483), .A2(n515), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U542 ( .A(G15GAT), .B(n482), .Z(G1326GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n485) );
  NAND2_X1 U544 ( .A1(n483), .A2(n512), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U546 ( .A(G22GAT), .B(n486), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .Z(n488) );
  NAND2_X1 U548 ( .A1(n490), .A2(n505), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  NAND2_X1 U550 ( .A1(n508), .A2(n490), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U552 ( .A1(n512), .A2(n490), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U554 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n495) );
  NOR2_X1 U555 ( .A1(n535), .A2(n551), .ZN(n492) );
  XOR2_X1 U556 ( .A(KEYINPUT106), .B(n492), .Z(n504) );
  NOR2_X1 U557 ( .A1(n504), .A2(n493), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n505), .A2(n499), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1332GAT) );
  XOR2_X1 U560 ( .A(G64GAT), .B(KEYINPUT107), .Z(n497) );
  NAND2_X1 U561 ( .A1(n499), .A2(n508), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(G1333GAT) );
  NAND2_X1 U563 ( .A1(n515), .A2(n499), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n498), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n501) );
  NAND2_X1 U566 ( .A1(n499), .A2(n512), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(n502), .ZN(G1335GAT) );
  XOR2_X1 U569 ( .A(G85GAT), .B(KEYINPUT109), .Z(n507) );
  NOR2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n511) );
  NAND2_X1 U571 ( .A1(n511), .A2(n505), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(G1336GAT) );
  NAND2_X1 U573 ( .A1(n508), .A2(n511), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n511), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT44), .ZN(n514) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(n514), .ZN(G1339GAT) );
  INV_X1 U580 ( .A(n515), .ZN(n518) );
  NAND2_X1 U581 ( .A1(n532), .A2(n516), .ZN(n517) );
  NOR2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(KEYINPUT112), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n535), .A2(n529), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G113GAT), .B(n520), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n522) );
  NAND2_X1 U587 ( .A1(n529), .A2(n537), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U589 ( .A(G120GAT), .B(n523), .Z(G1341GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n525) );
  XNOR2_X1 U591 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n529), .A2(n541), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n526), .B(KEYINPUT114), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(G134GAT), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U597 ( .A1(n529), .A2(n545), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1343GAT) );
  NAND2_X1 U599 ( .A1(n532), .A2(n556), .ZN(n533) );
  NOR2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n544), .A2(n535), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n539) );
  NAND2_X1 U604 ( .A1(n544), .A2(n537), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(n540), .ZN(G1345GAT) );
  XOR2_X1 U607 ( .A(G155GAT), .B(KEYINPUT117), .Z(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n541), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1346GAT) );
  NAND2_X1 U610 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n546), .B(KEYINPUT118), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G162GAT), .B(n547), .ZN(G1347GAT) );
  NOR2_X1 U613 ( .A1(n558), .A2(n554), .ZN(n548) );
  XOR2_X1 U614 ( .A(G169GAT), .B(n548), .Z(G1348GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n550) );
  XNOR2_X1 U616 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n551), .A2(n554), .ZN(n552) );
  XOR2_X1 U619 ( .A(n553), .B(n552), .Z(G1349GAT) );
  NOR2_X1 U620 ( .A1(n568), .A2(n554), .ZN(n555) );
  XOR2_X1 U621 ( .A(G183GAT), .B(n555), .Z(G1350GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n572) );
  NOR2_X1 U623 ( .A1(n558), .A2(n572), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U626 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1352GAT) );
  NOR2_X1 U628 ( .A1(n572), .A2(n563), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n565) );
  XNOR2_X1 U630 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1353GAT) );
  NOR2_X1 U633 ( .A1(n568), .A2(n572), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT126), .B(KEYINPUT127), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G211GAT), .B(n571), .ZN(G1354GAT) );
  NOR2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U638 ( .A(KEYINPUT62), .B(n574), .Z(n575) );
  XNOR2_X1 U639 ( .A(G218GAT), .B(n575), .ZN(G1355GAT) );
endmodule

