

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U323 ( .A(n438), .B(n437), .ZN(n550) );
  INV_X1 U324 ( .A(n570), .ZN(n439) );
  NOR2_X1 U325 ( .A1(n570), .A2(n569), .ZN(n572) );
  NOR2_X1 U326 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X2 U327 ( .A(KEYINPUT81), .B(n550), .ZN(n570) );
  XNOR2_X1 U328 ( .A(n339), .B(KEYINPUT74), .ZN(n426) );
  XNOR2_X1 U329 ( .A(G99GAT), .B(G85GAT), .ZN(n339) );
  XNOR2_X1 U330 ( .A(G190GAT), .B(G218GAT), .ZN(n391) );
  XNOR2_X1 U331 ( .A(n313), .B(n312), .ZN(n560) );
  XOR2_X1 U332 ( .A(KEYINPUT93), .B(KEYINPUT89), .Z(n291) );
  INV_X1 U333 ( .A(G71GAT), .ZN(n304) );
  INV_X1 U334 ( .A(KEYINPUT103), .ZN(n404) );
  XNOR2_X1 U335 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U336 ( .A(n404), .B(KEYINPUT26), .ZN(n405) );
  XNOR2_X1 U337 ( .A(n307), .B(n306), .ZN(n311) );
  XNOR2_X1 U338 ( .A(n406), .B(n405), .ZN(n576) );
  XOR2_X1 U339 ( .A(KEYINPUT38), .B(n464), .Z(n488) );
  XNOR2_X1 U340 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U341 ( .A(n468), .B(n467), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U343 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n399) );
  XOR2_X1 U345 ( .A(n399), .B(G134GAT), .Z(n295) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U347 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U348 ( .A(G190GAT), .B(n296), .ZN(n313) );
  XOR2_X1 U349 ( .A(KEYINPUT92), .B(KEYINPUT20), .Z(n298) );
  XNOR2_X1 U350 ( .A(G183GAT), .B(KEYINPUT91), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n301) );
  XNOR2_X1 U352 ( .A(G120GAT), .B(KEYINPUT90), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n291), .B(n299), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U355 ( .A(G176GAT), .B(G99GAT), .Z(n303) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U358 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n309) );
  XNOR2_X1 U359 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n364) );
  XNOR2_X1 U361 ( .A(n364), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n315) );
  XNOR2_X1 U364 ( .A(G1GAT), .B(KEYINPUT30), .ZN(n314) );
  XNOR2_X1 U365 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U366 ( .A(G29GAT), .B(G36GAT), .Z(n317) );
  XOR2_X1 U367 ( .A(G15GAT), .B(G22GAT), .Z(n457) );
  XNOR2_X1 U368 ( .A(n457), .B(KEYINPUT70), .ZN(n316) );
  XNOR2_X1 U369 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U370 ( .A(n319), .B(n318), .Z(n321) );
  NAND2_X1 U371 ( .A1(G229GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n325) );
  XOR2_X1 U373 ( .A(G197GAT), .B(G113GAT), .Z(n323) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(G50GAT), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U376 ( .A(n325), .B(n324), .Z(n333) );
  XOR2_X1 U377 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n327) );
  XNOR2_X1 U378 ( .A(KEYINPUT8), .B(G43GAT), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U380 ( .A(KEYINPUT7), .B(n328), .Z(n437) );
  XOR2_X1 U381 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n330) );
  XNOR2_X1 U382 ( .A(G141GAT), .B(G8GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n437), .B(n331), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n578) );
  XOR2_X1 U386 ( .A(KEYINPUT76), .B(KEYINPUT75), .Z(n335) );
  XNOR2_X1 U387 ( .A(KEYINPUT72), .B(KEYINPUT31), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n351) );
  XOR2_X1 U389 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n337) );
  NAND2_X1 U390 ( .A1(G230GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U392 ( .A(n338), .B(KEYINPUT73), .Z(n343) );
  XOR2_X1 U393 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n341) );
  XNOR2_X1 U394 ( .A(G71GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n449) );
  XNOR2_X1 U396 ( .A(n426), .B(n449), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U398 ( .A(G176GAT), .B(G64GAT), .Z(n396) );
  XOR2_X1 U399 ( .A(G92GAT), .B(n396), .Z(n345) );
  XOR2_X1 U400 ( .A(G120GAT), .B(G57GAT), .Z(n359) );
  XNOR2_X1 U401 ( .A(G106GAT), .B(n359), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U403 ( .A(n347), .B(n346), .Z(n349) );
  XNOR2_X1 U404 ( .A(G204GAT), .B(G148GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U406 ( .A(n351), .B(n350), .Z(n582) );
  NOR2_X1 U407 ( .A1(n578), .A2(n582), .ZN(n473) );
  XNOR2_X1 U408 ( .A(G155GAT), .B(KEYINPUT98), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n352), .B(KEYINPUT3), .ZN(n353) );
  XOR2_X1 U410 ( .A(n353), .B(KEYINPUT2), .Z(n355) );
  XNOR2_X1 U411 ( .A(G141GAT), .B(G148GAT), .ZN(n354) );
  XOR2_X1 U412 ( .A(n355), .B(n354), .Z(n385) );
  XOR2_X1 U413 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n357) );
  XNOR2_X1 U414 ( .A(G85GAT), .B(KEYINPUT6), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U416 ( .A(n385), .B(n358), .Z(n368) );
  XOR2_X1 U417 ( .A(G1GAT), .B(G127GAT), .Z(n445) );
  XOR2_X1 U418 ( .A(n445), .B(n359), .Z(n366) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(G134GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n360), .B(G162GAT), .ZN(n418) );
  XOR2_X1 U421 ( .A(n418), .B(KEYINPUT5), .Z(n362) );
  NAND2_X1 U422 ( .A1(G225GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U426 ( .A(n368), .B(n367), .ZN(n412) );
  XNOR2_X1 U427 ( .A(G211GAT), .B(KEYINPUT97), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n369), .B(KEYINPUT96), .ZN(n370) );
  XOR2_X1 U429 ( .A(n370), .B(KEYINPUT21), .Z(n372) );
  XNOR2_X1 U430 ( .A(G197GAT), .B(G204GAT), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n398) );
  XOR2_X1 U432 ( .A(KEYINPUT95), .B(KEYINPUT22), .Z(n374) );
  XNOR2_X1 U433 ( .A(G218GAT), .B(G162GAT), .ZN(n373) );
  XNOR2_X1 U434 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U435 ( .A(KEYINPUT23), .B(KEYINPUT99), .Z(n376) );
  XNOR2_X1 U436 ( .A(G22GAT), .B(G78GAT), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U438 ( .A(n378), .B(n377), .Z(n383) );
  XOR2_X1 U439 ( .A(G50GAT), .B(G106GAT), .Z(n425) );
  XOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n380) );
  NAND2_X1 U441 ( .A1(G228GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n425), .B(n381), .ZN(n382) );
  XNOR2_X1 U444 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n398), .B(n384), .ZN(n386) );
  XNOR2_X1 U446 ( .A(n386), .B(n385), .ZN(n553) );
  XOR2_X1 U447 ( .A(G8GAT), .B(G183GAT), .Z(n446) );
  INV_X1 U448 ( .A(G92GAT), .ZN(n387) );
  NAND2_X1 U449 ( .A1(KEYINPUT79), .A2(n387), .ZN(n390) );
  INV_X1 U450 ( .A(KEYINPUT79), .ZN(n388) );
  NAND2_X1 U451 ( .A1(n388), .A2(G92GAT), .ZN(n389) );
  NAND2_X1 U452 ( .A1(n390), .A2(n389), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U454 ( .A(G36GAT), .B(n393), .Z(n433) );
  XOR2_X1 U455 ( .A(n446), .B(n433), .Z(n395) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U458 ( .A(n397), .B(n396), .Z(n401) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U460 ( .A(n401), .B(n400), .ZN(n554) );
  NAND2_X1 U461 ( .A1(n560), .A2(n554), .ZN(n402) );
  NAND2_X1 U462 ( .A1(n553), .A2(n402), .ZN(n403) );
  XOR2_X1 U463 ( .A(KEYINPUT25), .B(n403), .Z(n408) );
  NOR2_X1 U464 ( .A1(n560), .A2(n553), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n554), .B(KEYINPUT27), .ZN(n413) );
  NAND2_X1 U466 ( .A1(n576), .A2(n413), .ZN(n407) );
  NAND2_X1 U467 ( .A1(n408), .A2(n407), .ZN(n409) );
  XOR2_X1 U468 ( .A(KEYINPUT104), .B(n409), .Z(n410) );
  NOR2_X1 U469 ( .A1(n412), .A2(n410), .ZN(n411) );
  XOR2_X1 U470 ( .A(KEYINPUT105), .B(n411), .Z(n417) );
  XNOR2_X1 U471 ( .A(KEYINPUT100), .B(n412), .ZN(n552) );
  NAND2_X1 U472 ( .A1(n413), .A2(n552), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n414), .B(KEYINPUT101), .ZN(n538) );
  XNOR2_X1 U474 ( .A(KEYINPUT28), .B(n553), .ZN(n480) );
  NAND2_X1 U475 ( .A1(n538), .A2(n480), .ZN(n525) );
  NOR2_X1 U476 ( .A1(n560), .A2(n525), .ZN(n415) );
  XNOR2_X1 U477 ( .A(KEYINPUT102), .B(n415), .ZN(n416) );
  NOR2_X1 U478 ( .A1(n417), .A2(n416), .ZN(n472) );
  NAND2_X1 U479 ( .A1(n418), .A2(KEYINPUT64), .ZN(n422) );
  INV_X1 U480 ( .A(n418), .ZN(n420) );
  INV_X1 U481 ( .A(KEYINPUT64), .ZN(n419) );
  NAND2_X1 U482 ( .A1(n420), .A2(n419), .ZN(n421) );
  NAND2_X1 U483 ( .A1(n422), .A2(n421), .ZN(n424) );
  AND2_X1 U484 ( .A1(G232GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U486 ( .A(KEYINPUT9), .B(KEYINPUT78), .Z(n428) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n436) );
  XOR2_X1 U490 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n432) );
  XNOR2_X1 U491 ( .A(KEYINPUT80), .B(KEYINPUT77), .ZN(n431) );
  XNOR2_X1 U492 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U493 ( .A(n434), .B(n433), .Z(n435) );
  XNOR2_X1 U494 ( .A(n436), .B(n435), .ZN(n438) );
  NAND2_X1 U495 ( .A1(KEYINPUT36), .A2(n570), .ZN(n442) );
  INV_X1 U496 ( .A(KEYINPUT36), .ZN(n440) );
  NAND2_X1 U497 ( .A1(n440), .A2(n439), .ZN(n441) );
  NAND2_X1 U498 ( .A1(n442), .A2(n441), .ZN(n512) );
  NOR2_X1 U499 ( .A1(n472), .A2(n512), .ZN(n462) );
  XOR2_X1 U500 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n444) );
  XNOR2_X1 U501 ( .A(G57GAT), .B(G64GAT), .ZN(n443) );
  XNOR2_X1 U502 ( .A(n444), .B(n443), .ZN(n461) );
  XOR2_X1 U503 ( .A(n446), .B(n445), .Z(n448) );
  XNOR2_X1 U504 ( .A(G211GAT), .B(G155GAT), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n453) );
  XOR2_X1 U506 ( .A(KEYINPUT84), .B(n449), .Z(n451) );
  NAND2_X1 U507 ( .A1(G231GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U509 ( .A(n453), .B(n452), .Z(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT85), .B(KEYINPUT82), .Z(n455) );
  XNOR2_X1 U511 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n461), .B(n460), .ZN(n587) );
  NAND2_X1 U516 ( .A1(n462), .A2(n587), .ZN(n463) );
  XNOR2_X1 U517 ( .A(KEYINPUT37), .B(n463), .ZN(n500) );
  NAND2_X1 U518 ( .A1(n473), .A2(n500), .ZN(n464) );
  NAND2_X1 U519 ( .A1(n560), .A2(n488), .ZN(n468) );
  XOR2_X1 U520 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n466) );
  XNOR2_X1 U521 ( .A(G43GAT), .B(KEYINPUT109), .ZN(n465) );
  INV_X1 U522 ( .A(n587), .ZN(n547) );
  NAND2_X1 U523 ( .A1(n547), .A2(n570), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT16), .ZN(n470) );
  XNOR2_X1 U525 ( .A(n470), .B(KEYINPUT86), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n491) );
  AND2_X1 U527 ( .A1(n473), .A2(n491), .ZN(n481) );
  NAND2_X1 U528 ( .A1(n552), .A2(n481), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT34), .ZN(n475) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n481), .A2(n554), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(KEYINPUT106), .ZN(n477) );
  XNOR2_X1 U533 ( .A(G8GAT), .B(n477), .ZN(G1325GAT) );
  XOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .Z(n479) );
  NAND2_X1 U535 ( .A1(n481), .A2(n560), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n479), .B(n478), .ZN(G1326GAT) );
  XOR2_X1 U537 ( .A(G22GAT), .B(KEYINPUT107), .Z(n483) );
  INV_X1 U538 ( .A(n480), .ZN(n507) );
  NAND2_X1 U539 ( .A1(n481), .A2(n507), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(G1327GAT) );
  XOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT39), .Z(n485) );
  NAND2_X1 U542 ( .A1(n488), .A2(n552), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  NAND2_X1 U544 ( .A1(n488), .A2(n554), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(KEYINPUT108), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G36GAT), .B(n487), .ZN(G1329GAT) );
  XOR2_X1 U547 ( .A(G50GAT), .B(KEYINPUT111), .Z(n490) );
  NAND2_X1 U548 ( .A1(n488), .A2(n507), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1331GAT) );
  INV_X1 U550 ( .A(n578), .ZN(n540) );
  XNOR2_X1 U551 ( .A(n582), .B(KEYINPUT41), .ZN(n564) );
  NOR2_X1 U552 ( .A1(n540), .A2(n564), .ZN(n501) );
  AND2_X1 U553 ( .A1(n501), .A2(n491), .ZN(n497) );
  NAND2_X1 U554 ( .A1(n497), .A2(n552), .ZN(n492) );
  XNOR2_X1 U555 ( .A(KEYINPUT42), .B(n492), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(n493), .ZN(G1332GAT) );
  NAND2_X1 U557 ( .A1(n497), .A2(n554), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(KEYINPUT112), .ZN(n495) );
  XNOR2_X1 U559 ( .A(G64GAT), .B(n495), .ZN(G1333GAT) );
  NAND2_X1 U560 ( .A1(n497), .A2(n560), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U562 ( .A(G78GAT), .B(KEYINPUT43), .Z(n499) );
  NAND2_X1 U563 ( .A1(n497), .A2(n507), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(G1335GAT) );
  NAND2_X1 U565 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(KEYINPUT113), .ZN(n508) );
  NAND2_X1 U567 ( .A1(n552), .A2(n508), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n503), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n554), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n504), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U571 ( .A1(n508), .A2(n560), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(KEYINPUT114), .ZN(n506) );
  XNOR2_X1 U573 ( .A(G99GAT), .B(n506), .ZN(G1338GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n510) );
  NAND2_X1 U575 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(G106GAT), .B(n511), .ZN(G1339GAT) );
  NOR2_X1 U578 ( .A1(n512), .A2(n587), .ZN(n513) );
  XOR2_X1 U579 ( .A(KEYINPUT45), .B(n513), .Z(n514) );
  NOR2_X1 U580 ( .A1(n582), .A2(n514), .ZN(n515) );
  XNOR2_X1 U581 ( .A(KEYINPUT116), .B(n515), .ZN(n516) );
  NAND2_X1 U582 ( .A1(n516), .A2(n578), .ZN(n522) );
  OR2_X1 U583 ( .A1(n550), .A2(n547), .ZN(n519) );
  NOR2_X1 U584 ( .A1(n578), .A2(n564), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n517), .B(KEYINPUT46), .ZN(n518) );
  NOR2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(KEYINPUT47), .B(n520), .ZN(n521) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(KEYINPUT48), .ZN(n524) );
  XNOR2_X1 U590 ( .A(KEYINPUT117), .B(n524), .ZN(n556) );
  NOR2_X1 U591 ( .A1(n556), .A2(n525), .ZN(n526) );
  NAND2_X1 U592 ( .A1(n526), .A2(n560), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(KEYINPUT118), .ZN(n534) );
  NOR2_X1 U594 ( .A1(n578), .A2(n534), .ZN(n528) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n528), .Z(G1340GAT) );
  NOR2_X1 U596 ( .A1(n534), .A2(n564), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n534), .A2(n587), .ZN(n532) );
  XNOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n531) );
  XNOR2_X1 U601 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  XNOR2_X1 U603 ( .A(KEYINPUT120), .B(KEYINPUT51), .ZN(n536) );
  NOR2_X1 U604 ( .A1(n570), .A2(n534), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(n537), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n538), .A2(n576), .ZN(n539) );
  NOR2_X1 U608 ( .A1(n556), .A2(n539), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n540), .A2(n549), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n541), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT121), .Z(n544) );
  INV_X1 U612 ( .A(n564), .ZN(n542) );
  NAND2_X1 U613 ( .A1(n549), .A2(n542), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n549), .A2(n547), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U621 ( .A(n552), .ZN(n575) );
  AND2_X1 U622 ( .A1(n575), .A2(n553), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT122), .B(n554), .Z(n555) );
  XNOR2_X1 U624 ( .A(KEYINPUT54), .B(n557), .ZN(n574) );
  NAND2_X1 U625 ( .A1(n558), .A2(n574), .ZN(n559) );
  XNOR2_X1 U626 ( .A(KEYINPUT55), .B(n559), .ZN(n561) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n569) );
  NOR2_X1 U628 ( .A1(n578), .A2(n569), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  NOR2_X1 U631 ( .A1(n564), .A2(n569), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(n567), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n587), .A2(n569), .ZN(n568) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  XNOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(G190GAT), .B(n573), .Z(G1351GAT) );
  AND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n591) );
  NOR2_X1 U642 ( .A1(n578), .A2(n591), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U647 ( .A(n591), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G204GAT), .B(n586), .Z(G1353GAT) );
  NOR2_X1 U651 ( .A1(n587), .A2(n591), .ZN(n588) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n588), .Z(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(n593) );
  NOR2_X1 U656 ( .A1(n512), .A2(n591), .ZN(n592) );
  XOR2_X1 U657 ( .A(n593), .B(n592), .Z(G1355GAT) );
endmodule

