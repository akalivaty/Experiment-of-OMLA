//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n568, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n600, new_n601,
    new_n602, new_n603, new_n605, new_n608, new_n609, new_n610, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n645, new_n646, new_n647, new_n648, new_n651, new_n653, new_n654,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n456), .A2(G2106), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(KEYINPUT68), .A3(new_n472), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n468), .A2(new_n473), .A3(G125), .ZN(new_n474));
  AND2_X1   g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G137), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(G137), .B(new_n480), .C1(new_n466), .C2(new_n467), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT69), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n470), .A2(G2105), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n479), .A2(new_n482), .B1(G101), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n476), .A2(new_n484), .ZN(G160));
  NAND2_X1  g060(.A1(new_n477), .A2(G136), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n480), .B1(new_n471), .B2(new_n472), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n480), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n486), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT70), .Z(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n468), .A2(new_n473), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n480), .C1(new_n466), .C2(new_n467), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n480), .A2(G114), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n502), .A2(new_n504), .A3(new_n505), .A4(G2104), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n501), .A2(new_n506), .B1(new_n487), .B2(G126), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n498), .A2(new_n507), .A3(KEYINPUT72), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT72), .B1(new_n498), .B2(new_n507), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT73), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT73), .A2(G651), .ZN(new_n513));
  OAI21_X1  g088(.A(KEYINPUT6), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT74), .B1(new_n519), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT5), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n520), .A2(new_n523), .B1(new_n519), .B2(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n511), .A2(new_n518), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(KEYINPUT73), .A2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT73), .A2(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n528), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n527), .A2(new_n533), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XOR2_X1   g110(.A(new_n535), .B(KEYINPUT7), .Z(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n536), .B1(new_n524), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n525), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n518), .A2(KEYINPUT75), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n517), .A2(new_n542), .A3(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n540), .B1(new_n544), .B2(G51), .ZN(G168));
  NAND2_X1  g120(.A1(new_n524), .A2(G64), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n532), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n515), .B1(new_n531), .B2(KEYINPUT6), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n519), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n521), .B1(KEYINPUT5), .B2(new_n522), .ZN(new_n551));
  NOR3_X1   g126(.A1(new_n519), .A2(KEYINPUT74), .A3(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n548), .A2(KEYINPUT76), .B1(new_n554), .B2(G90), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n546), .A2(new_n547), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(new_n531), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n542), .B1(new_n517), .B2(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(G52), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n555), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G171));
  AOI22_X1  g139(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G81), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n532), .B1(new_n525), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n544), .B2(G43), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  NAND4_X1  g144(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  AOI22_X1  g148(.A1(new_n524), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G651), .ZN(new_n575));
  INV_X1    g150(.A(G91), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n574), .A2(new_n575), .B1(new_n525), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(G53), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n517), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n582), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT77), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n580), .B1(new_n514), .B2(new_n516), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n579), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT9), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(new_n586), .B2(new_n585), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n583), .B(new_n584), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n582), .A2(KEYINPUT77), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n593), .B1(new_n529), .B2(new_n530), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n585), .B(new_n581), .C1(new_n594), .C2(new_n515), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT9), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n584), .B1(new_n597), .B2(new_n583), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n578), .B1(new_n591), .B2(new_n598), .ZN(G299));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n563), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n555), .A2(new_n559), .A3(KEYINPUT80), .A4(new_n562), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G301));
  NAND2_X1  g179(.A1(new_n544), .A2(G51), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n605), .B(new_n538), .C1(new_n539), .C2(new_n525), .ZN(G286));
  INV_X1    g181(.A(G166), .ZN(G303));
  OAI21_X1  g182(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n517), .A2(G49), .A3(G543), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n554), .A2(G87), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G288));
  AOI22_X1  g187(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(new_n532), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n517), .A2(new_n524), .A3(G86), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n517), .A2(G48), .A3(G543), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(G305));
  NAND2_X1  g193(.A1(new_n544), .A2(G47), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n554), .A2(G85), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n619), .B(new_n620), .C1(new_n532), .C2(new_n621), .ZN(G290));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NOR2_X1   g198(.A1(G301), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n554), .A2(G92), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT10), .Z(new_n626));
  NAND2_X1  g201(.A1(G79), .A2(G543), .ZN(new_n627));
  INV_X1    g202(.A(G66), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n553), .B2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT81), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g206(.A(KEYINPUT81), .B(new_n627), .C1(new_n553), .C2(new_n628), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(new_n632), .A3(G651), .ZN(new_n633));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n634));
  OAI21_X1  g209(.A(G54), .B1(new_n560), .B2(new_n561), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n634), .B1(new_n633), .B2(new_n635), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n626), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n626), .B(KEYINPUT83), .C1(new_n636), .C2(new_n637), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n624), .B1(new_n623), .B2(new_n642), .ZN(G284));
  AOI21_X1  g218(.A(new_n624), .B1(new_n623), .B2(new_n642), .ZN(G321));
  NAND2_X1  g219(.A1(G286), .A2(G868), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n583), .B1(new_n587), .B2(new_n589), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT79), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n577), .B1(new_n647), .B2(new_n590), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n645), .B1(new_n648), .B2(G868), .ZN(G297));
  OAI21_X1  g224(.A(new_n645), .B1(new_n648), .B2(G868), .ZN(G280));
  INV_X1    g225(.A(G559), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n642), .B1(new_n651), .B2(G860), .ZN(G148));
  NAND2_X1  g227(.A1(new_n642), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(G868), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g230(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g231(.A1(new_n468), .A2(new_n473), .A3(new_n483), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT12), .Z(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT13), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n477), .A2(G135), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n487), .A2(G123), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n480), .A2(G111), .ZN(new_n663));
  OAI21_X1  g238(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n664));
  OAI211_X1 g239(.A(new_n661), .B(new_n662), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n667), .ZN(G156));
  XNOR2_X1  g243(.A(G2427), .B(G2438), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2430), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT15), .B(G2435), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(KEYINPUT14), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT85), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2451), .B(G2454), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT16), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2443), .B(G2446), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n675), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1341), .B(G1348), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n683), .A3(G14), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G401));
  XNOR2_X1  g260(.A(G2072), .B(G2078), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT17), .ZN(new_n687));
  XOR2_X1   g262(.A(G2084), .B(G2090), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G2067), .B(G2678), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n687), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT86), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n693), .B(new_n689), .C1(new_n686), .C2(new_n690), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n688), .A2(new_n686), .A3(new_n690), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT18), .Z(new_n696));
  NAND3_X1  g271(.A1(new_n692), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G2096), .B(G2100), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G227));
  XOR2_X1   g274(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n700));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1956), .B(G2474), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1961), .B(G1966), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT20), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n703), .A2(new_n704), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n705), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n707), .B(new_n709), .C1(new_n702), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT88), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(G1991), .B(G1996), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(G229));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G20), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT23), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n648), .B2(new_n719), .ZN(new_n722));
  INV_X1    g297(.A(G1956), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT97), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G29), .B2(G32), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n477), .A2(G141), .B1(G105), .B2(new_n483), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n487), .A2(G129), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT26), .Z(new_n730));
  NAND3_X1  g305(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(new_n726), .B(new_n725), .S(new_n733), .Z(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  OR2_X1    g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  NAND2_X1  g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n737), .A2(new_n732), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n665), .B2(new_n732), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT100), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n732), .A2(G26), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT28), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n477), .A2(G140), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n487), .A2(G128), .ZN(new_n746));
  OR2_X1    g321(.A1(G104), .A2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n747), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2067), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR3_X1   g327(.A1(new_n736), .A2(new_n742), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G29), .A2(G35), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G162), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT29), .B(G2090), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G34), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G160), .B2(G29), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n757), .B1(G2084), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n761), .A2(G2084), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n755), .B2(new_n756), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n719), .A2(G19), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT93), .ZN(new_n766));
  INV_X1    g341(.A(new_n568), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1341), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n753), .A2(new_n762), .A3(new_n764), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT25), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n477), .A2(G139), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n468), .A2(new_n473), .A3(G127), .ZN(new_n776));
  INV_X1    g351(.A(G115), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n470), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n775), .B1(new_n778), .B2(G2105), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G29), .B2(G33), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(new_n442), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n442), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT96), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n771), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(G168), .A2(G16), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G21), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(KEYINPUT98), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(KEYINPUT98), .B2(new_n787), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  INV_X1    g366(.A(G1966), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n732), .A2(G27), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G164), .B2(new_n732), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT104), .B(G2078), .Z(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n768), .A2(new_n769), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G5), .A2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT102), .Z(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n563), .B2(new_n719), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT103), .B(G1961), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AOI211_X1 g378(.A(new_n798), .B(new_n803), .C1(new_n795), .C2(new_n797), .ZN(new_n804));
  AND4_X1   g379(.A1(new_n724), .A2(new_n786), .A3(new_n793), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n791), .A2(new_n792), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(KEYINPUT101), .Z(new_n807));
  NOR2_X1   g382(.A1(G4), .A2(G16), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n642), .B2(G16), .ZN(new_n809));
  INV_X1    g384(.A(G1348), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n805), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(G16), .A2(G24), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G290), .B2(new_n719), .ZN(new_n814));
  INV_X1    g389(.A(G1986), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT35), .B(G1991), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT90), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT91), .Z(new_n819));
  OAI21_X1  g394(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NOR3_X1   g396(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n822));
  OAI221_X1 g397(.A(G2104), .B1(G107), .B2(new_n480), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n477), .A2(G131), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n487), .A2(G119), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  MUX2_X1   g401(.A(G25), .B(new_n826), .S(G29), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n819), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n814), .A2(new_n815), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n816), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  MUX2_X1   g405(.A(G23), .B(G288), .S(G16), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT92), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT33), .B(G1976), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n719), .A2(G22), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G166), .B2(new_n719), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G1971), .Z(new_n839));
  MUX2_X1   g414(.A(G6), .B(G305), .S(G16), .Z(new_n840));
  XOR2_X1   g415(.A(KEYINPUT32), .B(G1981), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n835), .A2(new_n836), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n830), .B1(new_n843), .B2(KEYINPUT34), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(KEYINPUT34), .B2(new_n843), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT36), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n845), .A2(KEYINPUT36), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n812), .B1(new_n846), .B2(new_n847), .ZN(G311));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n846), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n849), .A2(new_n811), .A3(new_n807), .A4(new_n805), .ZN(G150));
  AOI22_X1  g425(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G93), .ZN(new_n852));
  OAI22_X1  g427(.A1(new_n851), .A2(new_n532), .B1(new_n525), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n544), .B2(G55), .ZN(new_n854));
  INV_X1    g429(.A(G860), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n642), .A2(G559), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n568), .B(new_n854), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n858), .B(KEYINPUT38), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n568), .B(new_n854), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n866), .A2(KEYINPUT105), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT105), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n855), .B1(new_n866), .B2(new_n867), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n857), .B1(new_n870), .B2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n826), .B(KEYINPUT107), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n658), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n477), .A2(G142), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n487), .A2(G130), .ZN(new_n877));
  OR2_X1    g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(G2104), .C1(G118), .C2(new_n480), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n658), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n873), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n875), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n875), .B2(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n886));
  OR3_X1    g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n886), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n779), .A2(KEYINPUT106), .A3(new_n731), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n731), .B1(new_n779), .B2(KEYINPUT106), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n498), .A2(new_n507), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n891), .A2(new_n892), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n749), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n894), .A2(new_n895), .A3(new_n749), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n887), .B(new_n888), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n887), .A2(new_n888), .ZN(new_n900));
  INV_X1    g475(.A(new_n898), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n896), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g478(.A(G162), .B(new_n665), .Z(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(G160), .Z(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n897), .A2(new_n898), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n907), .B2(new_n900), .ZN(new_n908));
  OAI22_X1  g483(.A1(new_n897), .A2(new_n898), .B1(new_n884), .B2(new_n885), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT109), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n905), .ZN(new_n911));
  AND4_X1   g486(.A1(KEYINPUT109), .A2(new_n902), .A3(new_n909), .A4(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n906), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(G395));
  NAND2_X1  g490(.A1(new_n653), .A2(new_n861), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n642), .A2(new_n651), .A3(new_n864), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n638), .A2(G299), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n638), .A2(G299), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n922), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(KEYINPUT41), .A3(new_n920), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n918), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n916), .B(new_n917), .C1(new_n921), .C2(new_n922), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT42), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(G305), .ZN(new_n931));
  XOR2_X1   g506(.A(G166), .B(G288), .Z(new_n932));
  OR2_X1    g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n927), .A2(new_n937), .A3(new_n928), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n930), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n930), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(new_n854), .A2(G868), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(G295));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n942), .ZN(G331));
  AOI21_X1  g519(.A(G286), .B1(new_n601), .B2(new_n602), .ZN(new_n945));
  NOR2_X1   g520(.A1(G171), .A2(G168), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n861), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n864), .B1(new_n945), .B2(new_n946), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n920), .A3(new_n949), .A4(new_n924), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n945), .A2(new_n864), .A3(new_n946), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n953), .B(new_n864), .C1(new_n945), .C2(new_n946), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n935), .B(new_n950), .C1(new_n955), .C2(new_n926), .ZN(new_n956));
  INV_X1    g531(.A(G37), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n935), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n933), .A2(KEYINPUT112), .A3(new_n934), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n948), .A2(new_n920), .A3(new_n924), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n963), .B1(new_n952), .B2(new_n954), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n948), .A2(new_n949), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n965), .A2(new_n923), .A3(new_n925), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n962), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n958), .A2(KEYINPUT43), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n950), .B1(new_n955), .B2(new_n926), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n962), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT43), .B1(new_n958), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT44), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n974), .A2(new_n967), .A3(new_n957), .A4(new_n956), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n958), .B2(new_n970), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n972), .A2(new_n977), .ZN(G397));
  AND3_X1   g553(.A1(new_n476), .A2(G40), .A3(new_n484), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n498), .B2(new_n507), .ZN(new_n980));
  XOR2_X1   g555(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n731), .B(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n749), .B(new_n751), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OR3_X1    g563(.A1(new_n988), .A2(new_n826), .A3(new_n818), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n749), .A2(G2067), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OR3_X1    g566(.A1(G290), .A2(new_n984), .A3(G1986), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT48), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n988), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n826), .B(new_n818), .Z(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n984), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n992), .A2(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n991), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n998), .A2(KEYINPUT46), .A3(new_n985), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT46), .B1(new_n998), .B2(new_n985), .ZN(new_n1002));
  INV_X1    g577(.A(new_n731), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n984), .B1(new_n1003), .B2(new_n987), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1000), .B1(new_n1006), .B2(KEYINPUT127), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(KEYINPUT127), .B2(new_n1006), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n979), .B(new_n1009), .C1(KEYINPUT45), .C2(new_n980), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n476), .A2(G40), .A3(new_n484), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT120), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1014), .B(new_n982), .C1(new_n508), .C2(new_n509), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n792), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n508), .B2(new_n509), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1012), .B1(new_n1018), .B2(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(G2084), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n892), .A2(new_n1014), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT115), .B1(new_n1021), .B2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n980), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1019), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1017), .A2(G168), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT51), .B1(new_n1028), .B2(G8), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(G168), .B1(new_n1017), .B2(new_n1027), .ZN(new_n1031));
  AND2_X1   g606(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1028), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1030), .B(KEYINPUT62), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT62), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1033), .A2(new_n1031), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(new_n1029), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(G2078), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1010), .A2(new_n1013), .A3(new_n1015), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1961), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1038), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1045));
  INV_X1    g620(.A(G1961), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(KEYINPUT124), .A3(new_n1041), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1050), .B(G1384), .C1(new_n498), .C2(new_n507), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1051), .B1(new_n1018), .B2(new_n981), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n979), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1039), .B1(new_n1053), .B2(G2078), .ZN(new_n1054));
  AOI21_X1  g629(.A(G301), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1056));
  NAND3_X1  g631(.A1(G303), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1056), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(G166), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G2090), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1019), .A2(new_n1062), .A3(new_n1026), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT114), .B(G1971), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1052), .B2(new_n979), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(new_n1061), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(G8), .B1(new_n1012), .B2(new_n1021), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n614), .A2(new_n1068), .A3(new_n617), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n613), .A2(new_n532), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n615), .A2(new_n616), .ZN(new_n1071));
  OAI21_X1  g646(.A(G1981), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT49), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1067), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(KEYINPUT49), .A3(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1067), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n610), .A2(KEYINPUT117), .A3(G1976), .A4(new_n611), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n610), .A2(G1976), .A3(new_n611), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1976), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT52), .B1(G288), .B2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1078), .A2(new_n1079), .A3(new_n1082), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1079), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT52), .B1(new_n1086), .B2(new_n1067), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1077), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1064), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1053), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1024), .B1(new_n892), .B2(new_n1014), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(new_n1012), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1024), .B(new_n1014), .C1(new_n508), .C2(new_n509), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n1062), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1059), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1066), .B(new_n1088), .C1(new_n1095), .C2(new_n1061), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1034), .A2(new_n1037), .A3(new_n1055), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1017), .A2(new_n1027), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(G8), .A3(G168), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1063), .A2(new_n1065), .A3(new_n1061), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1088), .A3(new_n1066), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1101), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1067), .B(KEYINPUT118), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n610), .A2(new_n1083), .A3(new_n611), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1069), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1077), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1066), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1110), .B(KEYINPUT119), .C1(new_n1066), .C2(new_n1111), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1104), .A2(new_n1105), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1098), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n476), .A2(new_n484), .A3(G40), .A4(new_n985), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1051), .B(new_n1119), .C1(new_n1018), .C2(new_n981), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT58), .B(G1341), .Z(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1012), .B2(new_n1021), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1018), .A2(new_n981), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1051), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1119), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(new_n1129), .A3(new_n1122), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT59), .B1(new_n1131), .B2(new_n568), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1133), .B(new_n767), .C1(new_n1124), .C2(new_n1130), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1125), .A2(new_n979), .A3(new_n1126), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n723), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n646), .A2(new_n578), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n648), .B2(new_n1141), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1145), .A2(new_n1137), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1144), .A2(KEYINPUT61), .A3(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n642), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1045), .A2(new_n810), .B1(new_n751), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1153), .A2(KEYINPUT60), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n642), .A2(KEYINPUT60), .A3(new_n1153), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1135), .A2(new_n1150), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1144), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1146), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1118), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT54), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT53), .B1(new_n443), .B2(KEYINPUT126), .ZN(new_n1164));
  AOI211_X1 g739(.A(new_n1164), .B(new_n1051), .C1(KEYINPUT126), .C2(new_n443), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n983), .A2(new_n1012), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1166), .A2(KEYINPUT125), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(KEYINPUT125), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1054), .A2(new_n1047), .A3(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1170), .A2(new_n603), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1163), .B1(new_n1055), .B2(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1036), .A2(new_n1096), .A3(new_n1029), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1049), .A2(G301), .A3(new_n1054), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1163), .B1(new_n1170), .B2(G171), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1172), .A2(new_n1173), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1162), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1159), .A2(new_n1118), .A3(new_n1161), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1117), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(G290), .B(new_n815), .ZN(new_n1181));
  INV_X1    g756(.A(new_n997), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n984), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1008), .B1(new_n1180), .B2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g759(.A1(G229), .A2(new_n463), .A3(G401), .A4(G227), .ZN(new_n1186));
  OAI211_X1 g760(.A(new_n1186), .B(new_n913), .C1(new_n975), .C2(new_n976), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


