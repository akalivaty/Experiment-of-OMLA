

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747;

  OR2_X1 U369 ( .A1(n556), .A2(n555), .ZN(n452) );
  NAND2_X1 U370 ( .A1(n368), .A2(n420), .ZN(n419) );
  XNOR2_X1 U371 ( .A(n458), .B(n456), .ZN(n563) );
  OR2_X1 U372 ( .A1(n638), .A2(G902), .ZN(n440) );
  XNOR2_X1 U373 ( .A(G137), .B(n511), .ZN(n462) );
  XNOR2_X1 U374 ( .A(n509), .B(n448), .ZN(n529) );
  NOR2_X1 U375 ( .A1(G953), .A2(G237), .ZN(n539) );
  XNOR2_X1 U376 ( .A(n449), .B(G128), .ZN(n509) );
  INV_X1 U377 ( .A(G143), .ZN(n449) );
  NAND2_X2 U378 ( .A1(n629), .A2(n628), .ZN(n714) );
  XNOR2_X1 U379 ( .A(n348), .B(n615), .ZN(n622) );
  NAND2_X1 U380 ( .A1(n406), .A2(n355), .ZN(n348) );
  XNOR2_X1 U381 ( .A(G113), .B(G143), .ZN(n533) );
  XOR2_X2 U382 ( .A(KEYINPUT4), .B(KEYINPUT69), .Z(n511) );
  NOR2_X1 U383 ( .A1(n707), .A2(n720), .ZN(n708) );
  NOR2_X1 U384 ( .A1(G953), .A2(n700), .ZN(n701) );
  AND2_X1 U385 ( .A1(n714), .A2(G210), .ZN(n634) );
  AND2_X1 U386 ( .A1(n369), .A2(n353), .ZN(n696) );
  NOR2_X1 U387 ( .A1(n721), .A2(n586), .ZN(n624) );
  AND2_X1 U388 ( .A1(n433), .A2(n665), .ZN(n733) );
  XNOR2_X1 U389 ( .A(n376), .B(n361), .ZN(n721) );
  AND2_X1 U390 ( .A1(n389), .A2(n391), .ZN(n385) );
  NOR2_X1 U391 ( .A1(n416), .A2(n421), .ZN(n604) );
  NOR2_X1 U392 ( .A1(n556), .A2(n402), .ZN(n573) );
  XNOR2_X1 U393 ( .A(n428), .B(n494), .ZN(n678) );
  NAND2_X1 U394 ( .A1(n566), .A2(n565), .ZN(n656) );
  XNOR2_X1 U395 ( .A(n451), .B(KEYINPUT32), .ZN(n450) );
  XNOR2_X1 U396 ( .A(n446), .B(G107), .ZN(n513) );
  XNOR2_X1 U397 ( .A(G116), .B(KEYINPUT72), .ZN(n480) );
  INV_X1 U398 ( .A(KEYINPUT65), .ZN(n451) );
  XNOR2_X2 U399 ( .A(n732), .B(n463), .ZN(n375) );
  XNOR2_X2 U400 ( .A(n529), .B(n462), .ZN(n732) );
  XNOR2_X1 U401 ( .A(n367), .B(G146), .ZN(n503) );
  INV_X1 U402 ( .A(G125), .ZN(n367) );
  NAND2_X1 U403 ( .A1(G214), .A2(n517), .ZN(n679) );
  NOR2_X1 U404 ( .A1(n702), .A2(G902), .ZN(n466) );
  XNOR2_X1 U405 ( .A(n415), .B(n476), .ZN(n571) );
  NOR2_X1 U406 ( .A1(n716), .A2(G902), .ZN(n415) );
  INV_X1 U407 ( .A(G146), .ZN(n463) );
  AND2_X1 U408 ( .A1(n425), .A2(n423), .ZN(n420) );
  NOR2_X1 U409 ( .A1(n445), .A2(n436), .ZN(n435) );
  OR2_X1 U410 ( .A1(G237), .A2(G902), .ZN(n517) );
  AND2_X1 U411 ( .A1(n399), .A2(n398), .ZN(n379) );
  XNOR2_X1 U412 ( .A(n576), .B(KEYINPUT105), .ZN(n398) );
  XNOR2_X1 U413 ( .A(KEYINPUT15), .B(G902), .ZN(n516) );
  XNOR2_X1 U414 ( .A(n562), .B(n430), .ZN(n429) );
  INV_X1 U415 ( .A(KEYINPUT106), .ZN(n430) );
  NAND2_X1 U416 ( .A1(n371), .A2(n667), .ZN(n670) );
  XNOR2_X1 U417 ( .A(G131), .B(KEYINPUT5), .ZN(n488) );
  INV_X1 U418 ( .A(KEYINPUT98), .ZN(n487) );
  XOR2_X1 U419 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n486) );
  XNOR2_X1 U420 ( .A(n515), .B(n727), .ZN(n630) );
  XNOR2_X1 U421 ( .A(n508), .B(n507), .ZN(n512) );
  XNOR2_X1 U422 ( .A(n426), .B(n605), .ZN(n607) );
  NOR2_X1 U423 ( .A1(n683), .A2(n682), .ZN(n426) );
  INV_X1 U424 ( .A(n656), .ZN(n418) );
  OR2_X1 U425 ( .A1(n425), .A2(n423), .ZN(n422) );
  BUF_X1 U426 ( .A(n618), .Z(n402) );
  NAND2_X1 U427 ( .A1(n387), .A2(n386), .ZN(n391) );
  AND2_X1 U428 ( .A1(n397), .A2(n453), .ZN(n386) );
  AND2_X1 U429 ( .A1(n396), .A2(n393), .ZN(n384) );
  NAND2_X1 U430 ( .A1(n387), .A2(n397), .ZN(n396) );
  XNOR2_X1 U431 ( .A(n551), .B(KEYINPUT22), .ZN(n556) );
  BUF_X1 U432 ( .A(n614), .Z(n400) );
  AND2_X1 U433 ( .A1(n373), .A2(n352), .ZN(n606) );
  XNOR2_X1 U434 ( .A(n374), .B(n360), .ZN(n373) );
  BUF_X1 U435 ( .A(n571), .Z(n365) );
  XNOR2_X1 U436 ( .A(n597), .B(n439), .ZN(n570) );
  INV_X1 U437 ( .A(KEYINPUT6), .ZN(n439) );
  XNOR2_X1 U438 ( .A(n514), .B(n380), .ZN(n727) );
  XNOR2_X1 U439 ( .A(n513), .B(n381), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n382), .B(G122), .ZN(n381) );
  INV_X1 U441 ( .A(KEYINPUT16), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n471), .B(n542), .ZN(n716) );
  XNOR2_X1 U443 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U444 ( .A(n411), .B(n408), .ZN(n470) );
  XNOR2_X1 U445 ( .A(n527), .B(n403), .ZN(n710) );
  XNOR2_X1 U446 ( .A(n404), .B(n528), .ZN(n403) );
  XOR2_X1 U447 ( .A(KEYINPUT9), .B(KEYINPUT101), .Z(n526) );
  XNOR2_X1 U448 ( .A(n465), .B(n455), .ZN(n454) );
  INV_X1 U449 ( .A(n513), .ZN(n455) );
  XNOR2_X1 U450 ( .A(n432), .B(n543), .ZN(n465) );
  INV_X1 U451 ( .A(n653), .ZN(n445) );
  XNOR2_X1 U452 ( .A(n438), .B(n437), .ZN(n436) );
  INV_X1 U453 ( .A(KEYINPUT47), .ZN(n437) );
  NOR2_X1 U454 ( .A1(n654), .A2(n684), .ZN(n438) );
  INV_X1 U455 ( .A(KEYINPUT46), .ZN(n444) );
  XNOR2_X1 U456 ( .A(n400), .B(n447), .ZN(n680) );
  INV_X1 U457 ( .A(KEYINPUT38), .ZN(n447) );
  NAND2_X1 U458 ( .A1(G234), .A2(G237), .ZN(n495) );
  INV_X1 U459 ( .A(KEYINPUT89), .ZN(n378) );
  XNOR2_X1 U460 ( .A(G101), .B(G119), .ZN(n482) );
  INV_X1 U461 ( .A(G134), .ZN(n448) );
  XNOR2_X1 U462 ( .A(KEYINPUT100), .B(KEYINPUT11), .ZN(n535) );
  XOR2_X1 U463 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n536) );
  XOR2_X1 U464 ( .A(G104), .B(G122), .Z(n534) );
  XNOR2_X1 U465 ( .A(n503), .B(n504), .ZN(n508) );
  XNOR2_X1 U466 ( .A(n506), .B(n505), .ZN(n507) );
  INV_X1 U467 ( .A(KEYINPUT18), .ZN(n505) );
  XNOR2_X1 U468 ( .A(n623), .B(KEYINPUT87), .ZN(n433) );
  NAND2_X1 U469 ( .A1(n680), .A2(n679), .ZN(n683) );
  AND2_X1 U470 ( .A1(n680), .A2(n372), .ZN(n425) );
  XNOR2_X1 U471 ( .A(n588), .B(KEYINPUT71), .ZN(n596) );
  NOR2_X1 U472 ( .A1(n521), .A2(KEYINPUT34), .ZN(n397) );
  XNOR2_X1 U473 ( .A(n427), .B(n356), .ZN(n614) );
  NAND2_X1 U474 ( .A1(n630), .A2(n516), .ZN(n427) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n411) );
  XNOR2_X1 U476 ( .A(G119), .B(G137), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n414), .B(G128), .ZN(n413) );
  INV_X1 U478 ( .A(G110), .ZN(n414) );
  XNOR2_X1 U479 ( .A(n410), .B(n409), .ZN(n408) );
  XNOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT73), .ZN(n410) );
  XNOR2_X1 U481 ( .A(G140), .B(KEYINPUT24), .ZN(n409) );
  XOR2_X1 U482 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n468) );
  INV_X1 U483 ( .A(n529), .ZN(n404) );
  XNOR2_X1 U484 ( .A(G116), .B(G122), .ZN(n522) );
  XOR2_X1 U485 ( .A(KEYINPUT7), .B(G107), .Z(n523) );
  INV_X1 U486 ( .A(n721), .ZN(n370) );
  XNOR2_X1 U487 ( .A(n464), .B(G101), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n431), .B(G140), .ZN(n543) );
  INV_X1 U489 ( .A(G131), .ZN(n431) );
  XNOR2_X1 U490 ( .A(G104), .B(G110), .ZN(n446) );
  XNOR2_X1 U491 ( .A(n493), .B(KEYINPUT33), .ZN(n494) );
  INV_X1 U492 ( .A(n607), .ZN(n693) );
  XOR2_X1 U493 ( .A(G478), .B(n532), .Z(n565) );
  NOR2_X1 U494 ( .A1(n670), .A2(n595), .ZN(n560) );
  XNOR2_X1 U495 ( .A(n457), .B(KEYINPUT0), .ZN(n456) );
  INV_X1 U496 ( .A(KEYINPUT68), .ZN(n457) );
  XNOR2_X1 U497 ( .A(n375), .B(n351), .ZN(n638) );
  XOR2_X1 U498 ( .A(n632), .B(n631), .Z(n633) );
  XNOR2_X1 U499 ( .A(n609), .B(n608), .ZN(n746) );
  XNOR2_X1 U500 ( .A(KEYINPUT115), .B(KEYINPUT42), .ZN(n608) );
  NAND2_X1 U501 ( .A1(n417), .A2(n419), .ZN(n600) );
  INV_X1 U502 ( .A(n421), .ZN(n417) );
  NOR2_X1 U503 ( .A1(n620), .A2(n617), .ZN(n593) );
  NAND2_X2 U504 ( .A1(n385), .A2(n383), .ZN(n743) );
  NAND2_X1 U505 ( .A1(n384), .A2(n388), .ZN(n383) );
  AND2_X1 U506 ( .A1(n357), .A2(n612), .ZN(n388) );
  XNOR2_X1 U507 ( .A(n574), .B(KEYINPUT104), .ZN(n744) );
  XNOR2_X1 U508 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U509 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U510 ( .A(n702), .B(n364), .ZN(n442) );
  AND2_X1 U511 ( .A1(n733), .A2(n626), .ZN(n349) );
  XOR2_X1 U512 ( .A(KEYINPUT108), .B(n547), .Z(n612) );
  AND2_X1 U513 ( .A1(n365), .A2(n549), .ZN(n350) );
  XNOR2_X1 U514 ( .A(n375), .B(n454), .ZN(n702) );
  INV_X1 U515 ( .A(n587), .ZN(n372) );
  XOR2_X1 U516 ( .A(n514), .B(n491), .Z(n351) );
  XOR2_X1 U517 ( .A(n595), .B(KEYINPUT110), .Z(n352) );
  OR2_X1 U518 ( .A1(n692), .A2(n691), .ZN(n353) );
  AND2_X1 U519 ( .A1(n571), .A2(n372), .ZN(n354) );
  AND2_X1 U520 ( .A1(n664), .A2(n435), .ZN(n355) );
  AND2_X1 U521 ( .A1(G210), .A2(n517), .ZN(n356) );
  AND2_X1 U522 ( .A1(n395), .A2(n392), .ZN(n357) );
  AND2_X1 U523 ( .A1(n370), .A2(n625), .ZN(n358) );
  XOR2_X1 U524 ( .A(n584), .B(KEYINPUT39), .Z(n359) );
  XNOR2_X1 U525 ( .A(KEYINPUT35), .B(KEYINPUT86), .ZN(n453) );
  XOR2_X1 U526 ( .A(n598), .B(KEYINPUT28), .Z(n360) );
  XOR2_X1 U527 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n361) );
  XOR2_X1 U528 ( .A(n638), .B(KEYINPUT62), .Z(n362) );
  NAND2_X1 U529 ( .A1(KEYINPUT90), .A2(n558), .ZN(n363) );
  XNOR2_X1 U530 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n364) );
  NOR2_X1 U531 ( .A1(G952), .A2(n735), .ZN(n720) );
  NOR2_X1 U532 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U533 ( .A1(n552), .A2(n553), .ZN(n554) );
  NAND2_X1 U534 ( .A1(n366), .A2(n610), .ZN(n407) );
  INV_X1 U535 ( .A(n742), .ZN(n366) );
  XNOR2_X1 U536 ( .A(n604), .B(n603), .ZN(n742) );
  XNOR2_X1 U537 ( .A(n591), .B(KEYINPUT109), .ZN(n592) );
  INV_X1 U538 ( .A(n583), .ZN(n368) );
  NAND2_X1 U539 ( .A1(n581), .A2(n582), .ZN(n583) );
  NAND2_X1 U540 ( .A1(n349), .A2(n370), .ZN(n369) );
  NAND2_X1 U541 ( .A1(n349), .A2(n358), .ZN(n629) );
  INV_X1 U542 ( .A(n571), .ZN(n371) );
  NAND2_X1 U543 ( .A1(n596), .A2(n597), .ZN(n374) );
  NAND2_X1 U544 ( .A1(n379), .A2(n377), .ZN(n376) );
  XNOR2_X1 U545 ( .A(n548), .B(n378), .ZN(n377) );
  INV_X1 U546 ( .A(n678), .ZN(n387) );
  AND2_X1 U547 ( .A1(n612), .A2(n395), .ZN(n394) );
  NAND2_X1 U548 ( .A1(n678), .A2(KEYINPUT34), .ZN(n393) );
  NAND2_X1 U549 ( .A1(n390), .A2(n453), .ZN(n389) );
  NAND2_X1 U550 ( .A1(n394), .A2(n393), .ZN(n390) );
  INV_X1 U551 ( .A(n453), .ZN(n392) );
  NAND2_X1 U552 ( .A1(n521), .A2(KEYINPUT34), .ZN(n395) );
  NAND2_X1 U553 ( .A1(n401), .A2(n559), .ZN(n399) );
  XNOR2_X1 U554 ( .A(n595), .B(n460), .ZN(n618) );
  XNOR2_X1 U555 ( .A(n519), .B(n518), .ZN(n599) );
  NAND2_X1 U556 ( .A1(n479), .A2(n618), .ZN(n562) );
  NAND2_X1 U557 ( .A1(n599), .A2(n520), .ZN(n458) );
  NAND2_X1 U558 ( .A1(n597), .A2(n679), .ZN(n580) );
  XNOR2_X2 U559 ( .A(n440), .B(n492), .ZN(n597) );
  NAND2_X1 U560 ( .A1(n419), .A2(n418), .ZN(n416) );
  XNOR2_X1 U561 ( .A(n407), .B(n444), .ZN(n406) );
  XNOR2_X1 U562 ( .A(n405), .B(n363), .ZN(n401) );
  NAND2_X1 U563 ( .A1(n744), .A2(n575), .ZN(n576) );
  AND2_X1 U564 ( .A1(n573), .A2(n365), .ZN(n557) );
  NAND2_X1 U565 ( .A1(n745), .A2(n650), .ZN(n405) );
  NAND2_X1 U566 ( .A1(n424), .A2(n422), .ZN(n421) );
  INV_X1 U567 ( .A(n359), .ZN(n423) );
  NAND2_X1 U568 ( .A1(n583), .A2(n359), .ZN(n424) );
  NOR2_X1 U569 ( .A1(n583), .A2(n587), .ZN(n611) );
  INV_X1 U570 ( .A(n400), .ZN(n620) );
  NAND2_X1 U571 ( .A1(n429), .A2(n570), .ZN(n428) );
  NAND2_X1 U572 ( .A1(n624), .A2(n433), .ZN(n626) );
  NAND2_X1 U573 ( .A1(n434), .A2(n402), .ZN(n664) );
  XNOR2_X1 U574 ( .A(n593), .B(KEYINPUT36), .ZN(n434) );
  AND2_X1 U575 ( .A1(n441), .A2(n640), .ZN(G54) );
  XNOR2_X1 U576 ( .A(n443), .B(n442), .ZN(n441) );
  NAND2_X1 U577 ( .A1(n714), .A2(G469), .ZN(n443) );
  XNOR2_X2 U578 ( .A(n452), .B(n450), .ZN(n745) );
  NAND2_X1 U579 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U580 ( .A(n639), .B(n362), .ZN(n641) );
  XNOR2_X1 U581 ( .A(n511), .B(n510), .ZN(n459) );
  XOR2_X1 U582 ( .A(KEYINPUT66), .B(KEYINPUT1), .Z(n460) );
  XOR2_X1 U583 ( .A(n705), .B(n704), .Z(n461) );
  INV_X1 U584 ( .A(n402), .ZN(n552) );
  XNOR2_X1 U585 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U586 ( .A(n490), .B(n489), .ZN(n491) );
  INV_X1 U587 ( .A(n670), .ZN(n479) );
  INV_X1 U588 ( .A(KEYINPUT111), .ZN(n598) );
  XNOR2_X1 U589 ( .A(n512), .B(n459), .ZN(n515) );
  INV_X1 U590 ( .A(KEYINPUT123), .ZN(n709) );
  XNOR2_X1 U591 ( .A(n602), .B(n601), .ZN(n603) );
  INV_X1 U592 ( .A(n720), .ZN(n640) );
  XNOR2_X1 U593 ( .A(n706), .B(n461), .ZN(n707) );
  XNOR2_X1 U594 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U595 ( .A(n642), .B(KEYINPUT63), .ZN(G57) );
  INV_X2 U596 ( .A(G953), .ZN(n735) );
  INV_X1 U597 ( .A(n516), .ZN(n625) );
  NAND2_X1 U598 ( .A1(G227), .A2(n735), .ZN(n464) );
  XNOR2_X2 U599 ( .A(n466), .B(G469), .ZN(n595) );
  XOR2_X1 U600 ( .A(KEYINPUT10), .B(n503), .Z(n542) );
  NAND2_X1 U601 ( .A1(G234), .A2(n735), .ZN(n467) );
  XNOR2_X1 U602 ( .A(n468), .B(n467), .ZN(n524) );
  NAND2_X1 U603 ( .A1(G221), .A2(n524), .ZN(n469) );
  XOR2_X1 U604 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n475) );
  NAND2_X1 U605 ( .A1(n516), .A2(G234), .ZN(n473) );
  XNOR2_X1 U606 ( .A(KEYINPUT20), .B(KEYINPUT96), .ZN(n472) );
  XNOR2_X1 U607 ( .A(n473), .B(n472), .ZN(n477) );
  NAND2_X1 U608 ( .A1(G217), .A2(n477), .ZN(n474) );
  XNOR2_X1 U609 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U610 ( .A1(n477), .A2(G221), .ZN(n478) );
  XNOR2_X1 U611 ( .A(KEYINPUT21), .B(n478), .ZN(n549) );
  INV_X1 U612 ( .A(n549), .ZN(n667) );
  XNOR2_X1 U613 ( .A(n480), .B(G113), .ZN(n484) );
  INV_X1 U614 ( .A(KEYINPUT3), .ZN(n481) );
  XNOR2_X1 U615 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U616 ( .A(n483), .B(n484), .ZN(n514) );
  NAND2_X1 U617 ( .A1(n539), .A2(G210), .ZN(n485) );
  XNOR2_X1 U618 ( .A(n486), .B(n485), .ZN(n490) );
  XNOR2_X1 U619 ( .A(G472), .B(KEYINPUT76), .ZN(n492) );
  XNOR2_X1 U620 ( .A(KEYINPUT107), .B(KEYINPUT74), .ZN(n493) );
  XNOR2_X1 U621 ( .A(n495), .B(KEYINPUT92), .ZN(n496) );
  XNOR2_X1 U622 ( .A(KEYINPUT14), .B(n496), .ZN(n498) );
  NAND2_X1 U623 ( .A1(G952), .A2(n498), .ZN(n692) );
  NOR2_X1 U624 ( .A1(G953), .A2(n692), .ZN(n497) );
  XOR2_X1 U625 ( .A(KEYINPUT93), .B(n497), .Z(n579) );
  AND2_X1 U626 ( .A1(n498), .A2(G953), .ZN(n499) );
  NAND2_X1 U627 ( .A1(G902), .A2(n499), .ZN(n577) );
  NOR2_X1 U628 ( .A1(G898), .A2(n577), .ZN(n500) );
  XNOR2_X1 U629 ( .A(n500), .B(KEYINPUT94), .ZN(n501) );
  NOR2_X1 U630 ( .A1(n579), .A2(n501), .ZN(n502) );
  XNOR2_X1 U631 ( .A(KEYINPUT95), .B(n502), .ZN(n520) );
  XNOR2_X1 U632 ( .A(KEYINPUT17), .B(KEYINPUT81), .ZN(n504) );
  NAND2_X1 U633 ( .A1(G224), .A2(n735), .ZN(n506) );
  INV_X1 U634 ( .A(n509), .ZN(n510) );
  NAND2_X1 U635 ( .A1(n614), .A2(n679), .ZN(n519) );
  XOR2_X1 U636 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n518) );
  INV_X1 U637 ( .A(n563), .ZN(n521) );
  XNOR2_X1 U638 ( .A(n523), .B(n522), .ZN(n528) );
  NAND2_X1 U639 ( .A1(G217), .A2(n524), .ZN(n525) );
  XNOR2_X1 U640 ( .A(n526), .B(n525), .ZN(n527) );
  NOR2_X1 U641 ( .A1(G902), .A2(n710), .ZN(n531) );
  XNOR2_X1 U642 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n530) );
  XNOR2_X1 U643 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U644 ( .A(n565), .ZN(n567) );
  XNOR2_X1 U645 ( .A(KEYINPUT13), .B(G475), .ZN(n546) );
  XNOR2_X1 U646 ( .A(n534), .B(n533), .ZN(n538) );
  XNOR2_X1 U647 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U648 ( .A(n538), .B(n537), .Z(n541) );
  NAND2_X1 U649 ( .A1(G214), .A2(n539), .ZN(n540) );
  XNOR2_X1 U650 ( .A(n541), .B(n540), .ZN(n544) );
  XNOR2_X1 U651 ( .A(n543), .B(n542), .ZN(n731) );
  XNOR2_X1 U652 ( .A(n731), .B(n544), .ZN(n703) );
  NOR2_X1 U653 ( .A1(G902), .A2(n703), .ZN(n545) );
  XOR2_X1 U654 ( .A(n546), .B(n545), .Z(n568) );
  INV_X1 U655 ( .A(n568), .ZN(n566) );
  NAND2_X1 U656 ( .A1(n567), .A2(n566), .ZN(n547) );
  NAND2_X1 U657 ( .A1(n743), .A2(KEYINPUT44), .ZN(n548) );
  INV_X1 U658 ( .A(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U659 ( .A1(n743), .A2(n558), .ZN(n559) );
  NAND2_X1 U660 ( .A1(n568), .A2(n565), .ZN(n682) );
  NOR2_X1 U661 ( .A1(n682), .A2(n549), .ZN(n550) );
  NAND2_X1 U662 ( .A1(n563), .A2(n550), .ZN(n551) );
  INV_X1 U663 ( .A(n570), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n589), .A2(n365), .ZN(n553) );
  XOR2_X1 U665 ( .A(KEYINPUT82), .B(n554), .Z(n555) );
  INV_X1 U666 ( .A(n597), .ZN(n669) );
  NAND2_X1 U667 ( .A1(n669), .A2(n557), .ZN(n650) );
  XOR2_X1 U668 ( .A(n560), .B(KEYINPUT97), .Z(n582) );
  AND2_X1 U669 ( .A1(n582), .A2(n563), .ZN(n561) );
  NAND2_X1 U670 ( .A1(n669), .A2(n561), .ZN(n644) );
  NOR2_X1 U671 ( .A1(n562), .A2(n669), .ZN(n675) );
  NAND2_X1 U672 ( .A1(n563), .A2(n675), .ZN(n564) );
  XOR2_X1 U673 ( .A(KEYINPUT31), .B(n564), .Z(n660) );
  NAND2_X1 U674 ( .A1(n644), .A2(n660), .ZN(n569) );
  NAND2_X1 U675 ( .A1(n568), .A2(n567), .ZN(n661) );
  NAND2_X1 U676 ( .A1(n656), .A2(n661), .ZN(n594) );
  NAND2_X1 U677 ( .A1(n569), .A2(n594), .ZN(n575) );
  NOR2_X1 U678 ( .A1(n365), .A2(n570), .ZN(n572) );
  NAND2_X1 U679 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U680 ( .A1(G900), .A2(n577), .ZN(n578) );
  NOR2_X1 U681 ( .A1(n579), .A2(n578), .ZN(n587) );
  XOR2_X1 U682 ( .A(KEYINPUT30), .B(n580), .Z(n581) );
  INV_X1 U683 ( .A(KEYINPUT75), .ZN(n584) );
  OR2_X1 U684 ( .A1(n600), .A2(n661), .ZN(n665) );
  NAND2_X1 U685 ( .A1(KEYINPUT2), .A2(n665), .ZN(n585) );
  XOR2_X1 U686 ( .A(KEYINPUT83), .B(n585), .Z(n586) );
  NAND2_X1 U687 ( .A1(n667), .A2(n354), .ZN(n588) );
  NOR2_X1 U688 ( .A1(n589), .A2(n656), .ZN(n590) );
  NAND2_X1 U689 ( .A1(n596), .A2(n590), .ZN(n591) );
  NAND2_X1 U690 ( .A1(n592), .A2(n679), .ZN(n617) );
  INV_X1 U691 ( .A(n594), .ZN(n684) );
  NAND2_X1 U692 ( .A1(n606), .A2(n599), .ZN(n654) );
  XNOR2_X1 U693 ( .A(KEYINPUT113), .B(KEYINPUT112), .ZN(n602) );
  INV_X1 U694 ( .A(KEYINPUT40), .ZN(n601) );
  XOR2_X1 U695 ( .A(KEYINPUT114), .B(KEYINPUT41), .Z(n605) );
  NAND2_X1 U696 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U697 ( .A(n746), .ZN(n610) );
  AND2_X1 U698 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n400), .A2(n613), .ZN(n653) );
  XOR2_X1 U700 ( .A(KEYINPUT70), .B(KEYINPUT48), .Z(n615) );
  NOR2_X1 U701 ( .A1(n402), .A2(n617), .ZN(n619) );
  XOR2_X1 U702 ( .A(KEYINPUT43), .B(n619), .Z(n621) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n666) );
  NAND2_X1 U704 ( .A1(n622), .A2(n666), .ZN(n623) );
  XOR2_X1 U705 ( .A(n625), .B(KEYINPUT85), .Z(n627) );
  AND2_X1 U706 ( .A1(n626), .A2(KEYINPUT2), .ZN(n698) );
  NAND2_X1 U707 ( .A1(n627), .A2(n698), .ZN(n628) );
  XOR2_X1 U708 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n632) );
  XNOR2_X1 U709 ( .A(n630), .B(KEYINPUT91), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n720), .A2(n635), .ZN(n637) );
  XNOR2_X1 U712 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(G51) );
  NAND2_X1 U714 ( .A1(n714), .A2(G472), .ZN(n639) );
  NOR2_X1 U715 ( .A1(n656), .A2(n644), .ZN(n643) );
  XOR2_X1 U716 ( .A(G104), .B(n643), .Z(G6) );
  NOR2_X1 U717 ( .A1(n661), .A2(n644), .ZN(n649) );
  XOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n646) );
  XNOR2_X1 U719 ( .A(G107), .B(KEYINPUT116), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U721 ( .A(KEYINPUT26), .B(n647), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(G9) );
  XNOR2_X1 U723 ( .A(G110), .B(n650), .ZN(G12) );
  NOR2_X1 U724 ( .A1(n661), .A2(n654), .ZN(n652) );
  XNOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n652), .B(n651), .ZN(G30) );
  XNOR2_X1 U727 ( .A(G143), .B(n653), .ZN(G45) );
  NOR2_X1 U728 ( .A1(n656), .A2(n654), .ZN(n655) );
  XOR2_X1 U729 ( .A(G146), .B(n655), .Z(G48) );
  NOR2_X1 U730 ( .A1(n656), .A2(n660), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(G113), .B(n659), .ZN(G15) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U735 ( .A(G116), .B(n662), .Z(G18) );
  XOR2_X1 U736 ( .A(G125), .B(KEYINPUT37), .Z(n663) );
  XNOR2_X1 U737 ( .A(n664), .B(n663), .ZN(G27) );
  XNOR2_X1 U738 ( .A(G134), .B(n665), .ZN(G36) );
  XNOR2_X1 U739 ( .A(G140), .B(n666), .ZN(G42) );
  XNOR2_X1 U740 ( .A(n350), .B(KEYINPUT49), .ZN(n668) );
  NAND2_X1 U741 ( .A1(n669), .A2(n668), .ZN(n673) );
  NAND2_X1 U742 ( .A1(n552), .A2(n670), .ZN(n671) );
  XOR2_X1 U743 ( .A(KEYINPUT50), .B(n671), .Z(n672) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U746 ( .A(KEYINPUT51), .B(n676), .Z(n677) );
  NOR2_X1 U747 ( .A1(n693), .A2(n677), .ZN(n689) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n686) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n678), .A2(n687), .ZN(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U754 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n693), .A2(n678), .ZN(n694) );
  XOR2_X1 U756 ( .A(KEYINPUT120), .B(n694), .Z(n695) );
  NAND2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U758 ( .A(n699), .B(KEYINPUT121), .ZN(n700) );
  XNOR2_X1 U759 ( .A(KEYINPUT53), .B(n701), .ZN(G75) );
  NAND2_X1 U760 ( .A1(G475), .A2(n714), .ZN(n706) );
  XOR2_X1 U761 ( .A(KEYINPUT67), .B(KEYINPUT122), .Z(n705) );
  XNOR2_X1 U762 ( .A(n703), .B(KEYINPUT59), .ZN(n704) );
  XNOR2_X1 U763 ( .A(KEYINPUT60), .B(n708), .ZN(G60) );
  NAND2_X1 U764 ( .A1(n714), .A2(G478), .ZN(n712) );
  XNOR2_X1 U765 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U766 ( .A1(n720), .A2(n713), .ZN(G63) );
  NAND2_X1 U767 ( .A1(G217), .A2(n714), .ZN(n718) );
  XOR2_X1 U768 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n715) );
  NOR2_X1 U769 ( .A1(n720), .A2(n719), .ZN(G66) );
  OR2_X1 U770 ( .A1(G953), .A2(n721), .ZN(n725) );
  NAND2_X1 U771 ( .A1(G953), .A2(G224), .ZN(n722) );
  XNOR2_X1 U772 ( .A(KEYINPUT61), .B(n722), .ZN(n723) );
  NAND2_X1 U773 ( .A1(n723), .A2(G898), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n725), .A2(n724), .ZN(n729) );
  NOR2_X1 U775 ( .A1(G898), .A2(n735), .ZN(n726) );
  NOR2_X1 U776 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U777 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U778 ( .A(KEYINPUT126), .B(n730), .ZN(G69) );
  XOR2_X1 U779 ( .A(n732), .B(n731), .Z(n737) );
  INV_X1 U780 ( .A(n737), .ZN(n734) );
  XOR2_X1 U781 ( .A(n734), .B(n733), .Z(n736) );
  NAND2_X1 U782 ( .A1(n736), .A2(n735), .ZN(n741) );
  XOR2_X1 U783 ( .A(G227), .B(n737), .Z(n738) );
  NAND2_X1 U784 ( .A1(n738), .A2(G900), .ZN(n739) );
  NAND2_X1 U785 ( .A1(n739), .A2(G953), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n741), .A2(n740), .ZN(G72) );
  XOR2_X1 U787 ( .A(n742), .B(G131), .Z(G33) );
  XOR2_X1 U788 ( .A(n743), .B(G122), .Z(G24) );
  XNOR2_X1 U789 ( .A(n744), .B(G101), .ZN(G3) );
  XNOR2_X1 U790 ( .A(n745), .B(G119), .ZN(G21) );
  XNOR2_X1 U791 ( .A(G137), .B(KEYINPUT127), .ZN(n747) );
  XNOR2_X1 U792 ( .A(n747), .B(n746), .ZN(G39) );
endmodule

