//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1204, new_n1205, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  INV_X1    g0006(.A(G244), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  OAI22_X1  g0009(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n202), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G116), .C2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G1), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(G50), .B1(G58), .B2(G68), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT64), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n221), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OR2_X1    g0031(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n223), .A2(G13), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n233), .B(G250), .C1(G257), .C2(G264), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  NAND4_X1  g0035(.A1(new_n226), .A2(new_n231), .A3(new_n232), .A4(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G226), .B(G232), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G250), .B(G257), .Z(new_n243));
  XNOR2_X1  g0043(.A(G264), .B(G270), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G58), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n229), .ZN(new_n257));
  NAND3_X1  g0057(.A1(KEYINPUT67), .A2(G33), .A3(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n220), .B1(G41), .B2(G45), .ZN(new_n260));
  AND3_X1   g0060(.A1(new_n259), .A2(KEYINPUT68), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT68), .B1(new_n259), .B2(new_n260), .ZN(new_n262));
  OAI21_X1  g0062(.A(G238), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT74), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n217), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT69), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n267), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(KEYINPUT69), .A3(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G232), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n272), .A2(new_n276), .B1(new_n277), .B2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n212), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n268), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n257), .A2(new_n254), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n263), .B(new_n266), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT13), .ZN(new_n284));
  INV_X1    g0084(.A(new_n282), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n272), .A2(new_n276), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n277), .A2(G1698), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n286), .A2(new_n280), .A3(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n288), .B2(new_n268), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT13), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(new_n266), .A4(new_n263), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT14), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n284), .A2(G179), .A3(new_n291), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT14), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n292), .A2(new_n296), .A3(G169), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT12), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n220), .A2(G13), .A3(G20), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(G68), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(KEYINPUT12), .A3(new_n213), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n229), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G1), .B2(new_n221), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n301), .B(new_n303), .C1(new_n307), .C2(new_n213), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT76), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n221), .A2(G33), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n312), .A2(new_n206), .B1(new_n221), .B2(G68), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT75), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G20), .A2(G33), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G50), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(KEYINPUT75), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n311), .B1(new_n319), .B2(new_n306), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(KEYINPUT11), .A3(new_n305), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n310), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n298), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT77), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n284), .A2(G190), .A3(new_n291), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G200), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n284), .B2(new_n291), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n325), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n329), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(KEYINPUT77), .A3(new_n326), .A4(new_n322), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n324), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  INV_X1    g0135(.A(new_n265), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n270), .A2(new_n271), .A3(new_n269), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT69), .B1(new_n274), .B2(new_n275), .ZN(new_n338));
  OAI21_X1  g0138(.A(G1698), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT70), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n286), .A2(KEYINPUT70), .A3(G1698), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(G238), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n286), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G107), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n286), .A2(G232), .A3(new_n279), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n336), .B1(new_n347), .B2(new_n285), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n261), .A2(new_n262), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G244), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT71), .B1(new_n348), .B2(new_n350), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n335), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G20), .A2(G77), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT8), .B(G58), .ZN(new_n355));
  INV_X1    g0155(.A(new_n315), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n354), .B1(new_n355), .B2(new_n356), .C1(new_n312), .C2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n305), .B1(new_n206), .B2(new_n302), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(new_n206), .B2(new_n307), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n347), .A2(new_n285), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n265), .A3(new_n350), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT71), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n350), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n353), .A2(new_n360), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n259), .A2(G232), .A3(new_n260), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  OAI211_X1 g0171(.A(G223), .B(new_n279), .C1(new_n270), .C2(new_n271), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT79), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n274), .A2(new_n275), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n375), .A2(KEYINPUT79), .A3(G223), .A4(new_n279), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(G226), .A3(G1698), .ZN(new_n377));
  AND4_X1   g0177(.A1(new_n371), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n265), .B(new_n370), .C1(new_n378), .C2(new_n282), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n328), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(G190), .B2(new_n379), .ZN(new_n381));
  XNOR2_X1  g0181(.A(G58), .B(G68), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n382), .A2(G20), .B1(G159), .B2(new_n315), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n270), .A2(new_n271), .A3(new_n384), .A4(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n272), .A2(new_n276), .A3(new_n221), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(new_n384), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n383), .B1(new_n387), .B2(new_n213), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n270), .A2(new_n271), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT7), .B1(new_n391), .B2(new_n221), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n392), .B2(new_n385), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n383), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n393), .A2(KEYINPUT78), .A3(new_n383), .A4(KEYINPUT16), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n390), .A2(new_n305), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(new_n355), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n307), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n399), .B2(new_n302), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n381), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT17), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n381), .A2(KEYINPUT17), .A3(new_n398), .A4(new_n401), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n398), .A2(new_n401), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n379), .A2(G169), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n335), .B2(new_n379), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n406), .A2(KEYINPUT18), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT18), .B1(new_n406), .B2(new_n408), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n404), .B(new_n405), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  OR3_X1    g0211(.A1(new_n334), .A2(new_n369), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n341), .A2(G223), .A3(new_n342), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n286), .A2(G222), .A3(new_n279), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n413), .B(new_n414), .C1(new_n206), .C2(new_n286), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n285), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n349), .A2(G226), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n416), .A2(G190), .A3(new_n265), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n203), .A2(G20), .ZN(new_n419));
  INV_X1    g0219(.A(G150), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n419), .B1(new_n420), .B2(new_n356), .C1(new_n355), .C2(new_n312), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n305), .B1(new_n202), .B2(new_n302), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n307), .A2(new_n202), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT9), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT9), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n426), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n418), .A2(KEYINPUT73), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n416), .A2(new_n265), .A3(new_n417), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(G200), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT73), .B1(new_n418), .B2(new_n428), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT10), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n425), .A2(KEYINPUT72), .A3(new_n427), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT72), .B1(new_n425), .B2(new_n427), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT10), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(new_n418), .A3(new_n431), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g0239(.A1(new_n430), .A2(new_n365), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n424), .B1(new_n430), .B2(G179), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n439), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(G190), .B1(new_n351), .B2(new_n352), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n364), .A2(G200), .A3(new_n366), .ZN(new_n446));
  INV_X1    g0246(.A(new_n360), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n302), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n267), .A2(G1), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n302), .A2(new_n305), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G116), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n221), .C1(G33), .C2(new_n217), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(new_n305), .C1(new_n221), .C2(G116), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT20), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n451), .B(new_n454), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  XOR2_X1   g0262(.A(KEYINPUT82), .B(G303), .Z(new_n463));
  NAND3_X1  g0263(.A1(new_n463), .A2(new_n272), .A3(new_n276), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n218), .A2(new_n279), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n375), .B(new_n465), .C1(G264), .C2(new_n279), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n282), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  INV_X1    g0269(.A(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT5), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G41), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n469), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n264), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n259), .A2(new_n474), .A3(G270), .ZN(new_n476));
  OR3_X1    g0276(.A1(new_n467), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n462), .A2(new_n477), .A3(new_n335), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(G169), .A3(new_n461), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT21), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n467), .A2(new_n475), .A3(new_n476), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n365), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT21), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(new_n461), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n478), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n468), .A2(new_n264), .A3(G1), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n214), .A2(new_n279), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n207), .A2(G1698), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n270), .C2(new_n271), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n267), .B2(new_n450), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n486), .B1(new_n490), .B2(new_n285), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n259), .B(G250), .C1(G1), .C2(new_n468), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(G190), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n375), .A2(new_n221), .A3(G68), .ZN(new_n494));
  INV_X1    g0294(.A(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n208), .A2(new_n217), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(KEYINPUT19), .B(new_n496), .C1(new_n268), .C2(G20), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n312), .B2(new_n217), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n305), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n357), .A2(new_n302), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n453), .A2(G87), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n491), .A2(new_n492), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(G200), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n491), .A2(G179), .A3(new_n492), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n490), .A2(new_n285), .ZN(new_n508));
  INV_X1    g0308(.A(new_n486), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n508), .A2(new_n509), .A3(new_n492), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n507), .B1(new_n510), .B2(new_n365), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n357), .B(KEYINPUT81), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n453), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(new_n502), .A3(new_n501), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n493), .A2(new_n506), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n481), .A2(G190), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n517), .B(new_n462), .C1(new_n328), .C2(new_n481), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n485), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n375), .A2(G244), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n520), .A2(new_n521), .B1(G33), .B2(G283), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n286), .A2(KEYINPUT4), .A3(G244), .A4(new_n279), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n521), .B1(new_n286), .B2(G250), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n522), .B(new_n523), .C1(new_n524), .C2(new_n279), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n285), .ZN(new_n526));
  INV_X1    g0326(.A(new_n475), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n259), .A2(new_n474), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G257), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n315), .A2(G77), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n387), .B2(new_n495), .ZN(new_n533));
  OR2_X1    g0333(.A1(KEYINPUT6), .A2(G97), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT80), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n536), .B1(new_n534), .B2(new_n535), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n495), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n539), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G107), .A3(new_n537), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n221), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n305), .B1(new_n533), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n300), .A2(G97), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n453), .A2(G97), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n525), .A2(new_n285), .B1(G257), .B2(new_n528), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(G190), .A3(new_n527), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n531), .A2(new_n547), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n530), .A2(new_n365), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n335), .A3(new_n527), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT25), .B1(new_n302), .B2(new_n495), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n302), .A2(KEYINPUT25), .A3(new_n495), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n558), .A2(new_n559), .B1(new_n453), .B2(G107), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT84), .ZN(new_n561));
  XNOR2_X1  g0361(.A(KEYINPUT83), .B(KEYINPUT24), .ZN(new_n562));
  AOI21_X1  g0362(.A(G20), .B1(new_n272), .B2(new_n276), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT22), .B1(new_n563), .B2(G87), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n221), .B2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n495), .A2(KEYINPUT23), .A3(G20), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(KEYINPUT22), .B(new_n221), .C1(new_n270), .C2(new_n271), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n565), .B(new_n569), .C1(new_n570), .C2(new_n208), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n562), .B1(new_n564), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n221), .B(G87), .C1(new_n337), .C2(new_n338), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT22), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n562), .ZN(new_n576));
  INV_X1    g0376(.A(new_n571), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n561), .B1(new_n579), .B2(new_n305), .ZN(new_n580));
  AOI211_X1 g0380(.A(KEYINPUT84), .B(new_n306), .C1(new_n572), .C2(new_n578), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n560), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n209), .A2(new_n279), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n218), .A2(G1698), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n270), .C2(new_n271), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G294), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n285), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n585), .B2(new_n587), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n527), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n259), .A2(new_n474), .A3(G264), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT86), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n259), .A2(new_n474), .A3(KEYINPUT86), .A4(G264), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(G169), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT87), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n591), .ZN(new_n600));
  AOI21_X1  g0400(.A(KEYINPUT88), .B1(new_n594), .B2(new_n595), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n594), .A2(KEYINPUT88), .A3(new_n595), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(G179), .A4(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(KEYINPUT87), .B(G169), .C1(new_n591), .C2(new_n596), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n582), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n560), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n564), .A2(new_n562), .A3(new_n571), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n576), .B1(new_n575), .B2(new_n577), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n305), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT84), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n579), .A2(new_n561), .A3(new_n305), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n594), .A2(KEYINPUT88), .A3(new_n595), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n601), .ZN(new_n616));
  AOI21_X1  g0416(.A(G200), .B1(new_n616), .B2(new_n600), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT89), .ZN(new_n618));
  INV_X1    g0418(.A(G190), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n594), .A2(new_n595), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n600), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n585), .A2(new_n587), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT85), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(new_n285), .A3(new_n588), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(new_n620), .A3(new_n619), .A4(new_n527), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT89), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n614), .B1(new_n617), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n519), .A2(new_n556), .A3(new_n607), .A4(new_n628), .ZN(new_n629));
  NOR4_X1   g0429(.A1(new_n412), .A2(new_n444), .A3(new_n449), .A4(new_n629), .ZN(G372));
  NOR3_X1   g0430(.A1(new_n412), .A2(new_n444), .A3(new_n449), .ZN(new_n631));
  INV_X1    g0431(.A(new_n504), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n505), .A2(G200), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n632), .A2(new_n633), .A3(new_n493), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT90), .ZN(new_n635));
  AND4_X1   g0435(.A1(G179), .A2(new_n508), .A3(new_n509), .A4(new_n492), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n365), .B1(new_n491), .B2(new_n492), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(KEYINPUT90), .B(new_n507), .C1(new_n510), .C2(new_n365), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n634), .B1(new_n640), .B2(new_n515), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n627), .A2(new_n617), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n582), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n551), .A2(new_n555), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n599), .A2(new_n604), .A3(new_n605), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n485), .B1(new_n614), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT91), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n607), .A2(KEYINPUT91), .A3(new_n485), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n645), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n640), .A2(new_n515), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n516), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(KEYINPUT26), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n553), .A2(new_n554), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n641), .A2(new_n655), .A3(new_n656), .A4(new_n552), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n631), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n409), .A2(new_n410), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n369), .A2(new_n333), .B1(new_n323), .B2(new_n298), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n404), .A2(new_n405), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n661), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n442), .B1(new_n665), .B2(new_n439), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n660), .A2(new_n666), .ZN(G369));
  NOR2_X1   g0467(.A1(new_n582), .A2(new_n642), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n607), .B2(new_n485), .ZN(new_n669));
  INV_X1    g0469(.A(G13), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n220), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n669), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n485), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n462), .A2(new_n678), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n461), .A2(new_n677), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n485), .A2(new_n518), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n684), .B2(KEYINPUT92), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(KEYINPUT92), .B2(new_n682), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n607), .A2(new_n678), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n668), .B1(new_n582), .B2(new_n606), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n582), .A2(new_n677), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n679), .B1(new_n687), .B2(new_n691), .ZN(G399));
  NAND3_X1  g0492(.A1(new_n641), .A2(new_n655), .A3(new_n552), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n652), .B1(new_n693), .B2(KEYINPUT26), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n669), .A2(new_n556), .ZN(new_n695));
  OAI221_X1 g0495(.A(new_n694), .B1(KEYINPUT26), .B2(new_n653), .C1(new_n695), .C2(new_n634), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n696), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n677), .B1(new_n651), .B2(new_n658), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n510), .A2(G179), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n530), .A2(new_n477), .A3(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n615), .A2(new_n591), .A3(new_n601), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n526), .A2(new_n529), .A3(new_n481), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n636), .A2(new_n600), .A3(new_n602), .A4(new_n603), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT95), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT96), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT30), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n703), .A2(new_n549), .A3(new_n636), .A4(new_n481), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT96), .B1(new_n710), .B2(KEYINPUT95), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT30), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n710), .B2(KEYINPUT96), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n704), .B(new_n709), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n677), .ZN(new_n715));
  OAI211_X1 g0515(.A(KEYINPUT31), .B(new_n715), .C1(new_n629), .C2(new_n677), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n700), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n220), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT93), .ZN(new_n723));
  INV_X1    g0523(.A(new_n233), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(G41), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n233), .A2(KEYINPUT93), .A3(new_n470), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n496), .A2(G116), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(G1), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n227), .B2(new_n727), .ZN(new_n730));
  XOR2_X1   g0530(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n731));
  XNOR2_X1  g0531(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n722), .A2(new_n732), .ZN(G364));
  INV_X1    g0533(.A(new_n727), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n220), .B1(new_n671), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n229), .B1(G20), .B2(new_n365), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n335), .A2(G200), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT98), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(new_n221), .A3(new_n619), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G87), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n742), .A2(new_n221), .A3(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n744), .B(new_n286), .C1(new_n746), .C2(new_n495), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT99), .Z(new_n748));
  NOR2_X1   g0548(.A1(new_n221), .A2(new_n619), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n335), .A2(new_n328), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n335), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(G50), .A2(new_n752), .B1(new_n755), .B2(G58), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n221), .A2(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n750), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n753), .A2(new_n757), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n756), .B1(new_n213), .B2(new_n758), .C1(new_n206), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n221), .B1(new_n761), .B2(G190), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(G97), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n757), .A2(new_n761), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n748), .A2(new_n764), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G294), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n344), .B1(new_n771), .B2(new_n762), .ZN(new_n772));
  INV_X1    g0572(.A(new_n765), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G329), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  INV_X1    g0575(.A(G322), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n774), .B1(new_n775), .B2(new_n759), .C1(new_n776), .C2(new_n754), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n772), .B(new_n777), .C1(G326), .C2(new_n752), .ZN(new_n778));
  INV_X1    g0578(.A(new_n758), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT100), .B(KEYINPUT33), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(G317), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n745), .A2(G283), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  INV_X1    g0583(.A(new_n743), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n778), .B(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n739), .B1(new_n770), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n738), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n724), .A2(new_n375), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(new_n228), .B2(new_n468), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n249), .B2(new_n468), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n286), .A2(new_n233), .A3(G355), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(G116), .C2(new_n233), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n786), .B1(new_n790), .B2(new_n796), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n789), .B(KEYINPUT101), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n737), .B(new_n797), .C1(new_n686), .C2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n737), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n687), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n686), .A2(G330), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G396));
  AND4_X1   g0604(.A1(new_n360), .A2(new_n353), .A3(new_n367), .A4(new_n678), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n360), .A2(new_n677), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT103), .Z(new_n807));
  NAND2_X1  g0607(.A1(new_n448), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n805), .B1(new_n368), .B2(new_n808), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n698), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n698), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n720), .ZN(new_n813));
  INV_X1    g0613(.A(G330), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n718), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(new_n810), .A3(new_n811), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n816), .A3(new_n801), .ZN(new_n817));
  INV_X1    g0617(.A(G58), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n375), .B1(new_n762), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n746), .A2(new_n213), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(G50), .C2(new_n743), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G143), .A2(new_n755), .B1(new_n779), .B2(G150), .ZN(new_n822));
  INV_X1    g0622(.A(G137), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(new_n823), .B2(new_n751), .C1(new_n766), .C2(new_n759), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT34), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n821), .B(new_n825), .C1(new_n826), .C2(new_n765), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n758), .A2(new_n828), .B1(new_n762), .B2(new_n217), .ZN(new_n829));
  INV_X1    g0629(.A(new_n759), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n286), .B(new_n829), .C1(G116), .C2(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n751), .A2(new_n783), .B1(new_n754), .B2(new_n771), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n745), .B2(G87), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n773), .A2(G311), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n743), .A2(G107), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n831), .A2(new_n833), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n739), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n738), .A2(new_n787), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n801), .B(new_n837), .C1(new_n206), .C2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT102), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n788), .B2(new_n809), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n817), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n842), .A2(KEYINPUT104), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(KEYINPUT104), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(G384));
  NAND2_X1  g0646(.A1(new_n406), .A2(new_n408), .ZN(new_n847));
  INV_X1    g0647(.A(new_n675), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n406), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n402), .A2(new_n847), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n396), .A2(new_n305), .A3(new_n397), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT16), .B1(new_n393), .B2(new_n383), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n401), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n848), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n402), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n408), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n851), .B1(new_n857), .B2(new_n850), .ZN(new_n858));
  INV_X1    g0658(.A(new_n855), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n411), .A2(KEYINPUT106), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT106), .B1(new_n411), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT38), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n858), .B(KEYINPUT38), .C1(new_n860), .C2(new_n861), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n323), .A2(new_n677), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n334), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n324), .A2(new_n333), .A3(new_n867), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT105), .ZN(new_n872));
  INV_X1    g0672(.A(new_n805), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n811), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n808), .A2(new_n368), .ZN(new_n875));
  AOI211_X1 g0675(.A(KEYINPUT105), .B(new_n805), .C1(new_n698), .C2(new_n875), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n866), .B(new_n871), .C1(new_n874), .C2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n661), .A2(new_n848), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT107), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n402), .A2(new_n847), .A3(new_n849), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT37), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(KEYINPUT108), .A3(new_n851), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT108), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(new_n885), .A3(KEYINPUT37), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n849), .B1(new_n663), .B2(new_n661), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n863), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n865), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n864), .A2(KEYINPUT39), .A3(new_n865), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n324), .A2(new_n677), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n877), .A2(KEYINPUT107), .A3(new_n878), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n881), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n631), .A2(new_n697), .A3(new_n699), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n666), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n875), .A2(new_n873), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n324), .A2(new_n333), .A3(new_n867), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n867), .B1(new_n324), .B2(new_n333), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n890), .A2(new_n906), .A3(new_n719), .A4(KEYINPUT40), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n871), .A2(new_n809), .A3(new_n716), .A4(new_n717), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT40), .B1(new_n866), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n631), .A2(new_n719), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n912), .B(new_n913), .Z(new_n914));
  NOR2_X1   g0714(.A1(new_n914), .A2(new_n814), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n901), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n220), .B2(new_n671), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n540), .A2(new_n542), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n450), .B1(new_n918), .B2(KEYINPUT35), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n230), .C1(KEYINPUT35), .C2(new_n918), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  OAI21_X1  g0721(.A(G77), .B1(new_n818), .B2(new_n213), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n922), .A2(new_n227), .B1(G50), .B2(new_n213), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G1), .A3(new_n670), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n917), .A2(new_n921), .A3(new_n924), .ZN(G367));
  NAND3_X1  g0725(.A1(new_n689), .A2(new_n680), .A3(new_n678), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n554), .A2(new_n677), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n556), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT42), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n555), .B1(new_n928), .B2(new_n607), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n678), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT111), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(KEYINPUT111), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT112), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT109), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n641), .B1(new_n632), .B2(new_n678), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n652), .A2(new_n504), .A3(new_n677), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT110), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n934), .A2(new_n935), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n941), .A2(new_n942), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n687), .A2(new_n691), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n928), .B1(new_n555), .B2(new_n678), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n945), .A2(new_n948), .A3(new_n949), .A4(new_n946), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n936), .B2(new_n944), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n727), .B(KEYINPUT41), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n949), .A2(new_n679), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT45), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n679), .A2(new_n556), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n948), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n691), .B1(new_n485), .B2(new_n677), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n926), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(new_n687), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n721), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n955), .B1(new_n966), .B2(new_n721), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n735), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n944), .A2(new_n936), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n951), .A2(new_n969), .A3(new_n952), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n954), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(G143), .ZN(new_n972));
  OAI22_X1  g0772(.A1(new_n751), .A2(new_n972), .B1(new_n759), .B2(new_n202), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n746), .A2(new_n206), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G58), .C2(new_n743), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n823), .A2(new_n765), .B1(new_n762), .B2(new_n213), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n976), .B(new_n344), .C1(G159), .C2(new_n779), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(new_n420), .C2(new_n754), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G311), .A2(new_n752), .B1(new_n779), .B2(G294), .ZN(new_n979));
  INV_X1    g0779(.A(new_n463), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n979), .B1(new_n828), .B2(new_n759), .C1(new_n980), .C2(new_n754), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n375), .B(new_n981), .C1(G107), .C2(new_n763), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n743), .A2(G116), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n217), .C2(new_n746), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n765), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n978), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n801), .B1(new_n989), .B2(new_n738), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n790), .B1(new_n233), .B2(new_n357), .C1(new_n792), .C2(new_n245), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n941), .A2(new_n798), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n971), .A2(new_n993), .ZN(G387));
  AOI21_X1  g0794(.A(new_n727), .B1(new_n721), .B2(new_n964), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n965), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G311), .A2(new_n779), .B1(new_n755), .B2(G317), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n776), .B2(new_n751), .C1(new_n980), .C2(new_n759), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT48), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n828), .B2(new_n762), .C1(new_n771), .C2(new_n784), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n773), .A2(G326), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n375), .B1(new_n745), .B2(G116), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n765), .A2(new_n420), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n206), .A2(new_n784), .B1(new_n746), .B2(new_n217), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n375), .B1(new_n759), .B2(new_n213), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n751), .A2(new_n766), .B1(new_n758), .B2(new_n355), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n512), .A2(new_n762), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(G50), .B2(new_n755), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(KEYINPUT113), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1006), .B1(new_n1007), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n801), .B1(new_n1017), .B2(new_n738), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n728), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n399), .A2(new_n202), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n1021), .B(new_n468), .C1(KEYINPUT50), .C2(new_n1020), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G68), .B2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n791), .B1(new_n242), .B2(new_n468), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n286), .A2(new_n1019), .A3(new_n233), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n233), .A2(G107), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n790), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n691), .A2(new_n798), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1018), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n996), .B(new_n1030), .C1(new_n735), .C2(new_n964), .ZN(G393));
  XNOR2_X1  g0831(.A(new_n961), .B(KEYINPUT115), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n736), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n391), .B1(new_n773), .B2(G143), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n784), .B2(new_n213), .C1(new_n208), .C2(new_n746), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT116), .Z(new_n1036));
  NAND2_X1  g0836(.A1(new_n830), .A2(new_n399), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n751), .A2(new_n420), .B1(new_n754), .B2(new_n766), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT51), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n779), .A2(G50), .B1(new_n763), .B2(G77), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n751), .A2(new_n986), .B1(new_n754), .B2(new_n775), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n746), .B2(new_n495), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G283), .B2(new_n743), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n980), .A2(new_n758), .B1(new_n771), .B2(new_n759), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n344), .B1(new_n450), .B2(new_n762), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G322), .C2(new_n773), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1046), .B(new_n1049), .C1(new_n1043), .C2(new_n1042), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n801), .B1(new_n1051), .B2(new_n738), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n790), .B1(new_n217), .B2(new_n233), .C1(new_n792), .C2(new_n252), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n789), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1053), .C1(new_n949), .C2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n727), .B1(new_n961), .B2(new_n965), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n961), .B2(new_n965), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1033), .A2(new_n1055), .A3(new_n1057), .ZN(G390));
  AOI21_X1  g0858(.A(new_n805), .B1(new_n698), .B2(new_n875), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(new_n872), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n815), .A2(new_n906), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n871), .B1(new_n815), .B2(new_n809), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n905), .B1(new_n720), .B2(new_n902), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n696), .A2(new_n678), .A3(new_n875), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n873), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1068), .A3(new_n1061), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1064), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n631), .A2(G330), .A3(new_n719), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n899), .A2(new_n1071), .A3(new_n666), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT117), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n736), .B1(new_n1074), .B2(new_n734), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n871), .B1(new_n874), .B2(new_n876), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n895), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1076), .A2(new_n1077), .B1(new_n892), .B2(new_n893), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n889), .A2(new_n865), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n895), .B(new_n1079), .C1(new_n1067), .C2(new_n871), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1062), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1077), .B(new_n890), .C1(new_n1068), .C2(new_n905), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n895), .B1(new_n1060), .B2(new_n871), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n1061), .C1(new_n1083), .C2(new_n894), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1075), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1081), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n727), .B2(new_n1074), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT54), .B(G143), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n754), .A2(new_n826), .B1(new_n759), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n344), .B1(G125), .B2(new_n773), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1091), .B1(new_n1092), .B2(new_n751), .C1(new_n766), .C2(new_n762), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1090), .B(new_n1093), .C1(G50), .C2(new_n745), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n743), .A2(G150), .ZN(new_n1095));
  XOR2_X1   g0895(.A(new_n1095), .B(KEYINPUT53), .Z(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n1096), .C1(new_n823), .C2(new_n758), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT118), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n820), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n771), .A2(new_n765), .B1(new_n762), .B2(new_n206), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n286), .B(new_n1100), .C1(G107), .C2(new_n779), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n751), .A2(new_n828), .B1(new_n759), .B2(new_n217), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G116), .B2(new_n755), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n744), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1098), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n801), .B1(new_n1105), .B2(new_n738), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n838), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1106), .B1(new_n399), .B2(new_n1107), .C1(new_n894), .C2(new_n788), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1088), .A2(new_n1108), .ZN(G378));
  NAND3_X1  g0909(.A1(new_n1084), .A2(new_n1081), .A3(new_n1070), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1073), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n444), .A2(KEYINPUT55), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT55), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n439), .A2(new_n1113), .A3(new_n443), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n424), .A2(new_n848), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1112), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1115), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1113), .B1(new_n439), .B2(new_n443), .ZN(new_n1118));
  AOI211_X1 g0918(.A(KEYINPUT55), .B(new_n442), .C1(new_n434), .C2(new_n438), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1116), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n912), .A2(KEYINPUT122), .A3(G330), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n909), .B1(new_n865), .B2(new_n864), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n907), .C1(new_n1128), .C2(KEYINPUT40), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT122), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1116), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1122), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1134), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1127), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n881), .A2(new_n896), .A3(new_n897), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n911), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1139), .A2(KEYINPUT122), .A3(G330), .A4(new_n907), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(new_n1134), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n898), .B1(new_n1142), .B2(new_n1127), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1111), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT57), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(KEYINPUT57), .B(new_n1111), .C1(new_n1138), .C2(new_n1143), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(new_n734), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n898), .A2(new_n1142), .A3(new_n1127), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n735), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n391), .B1(new_n784), .B2(new_n206), .C1(new_n818), .C2(new_n746), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n512), .A2(new_n759), .B1(new_n217), .B2(new_n758), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT119), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G116), .A2(new_n752), .B1(new_n755), .B2(G107), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n213), .B2(new_n762), .C1(new_n828), .C2(new_n765), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1152), .A2(new_n1154), .A3(G41), .A4(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT58), .Z(new_n1158));
  OAI21_X1  g0958(.A(new_n202), .B1(new_n270), .B2(G41), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G33), .B1(new_n773), .B2(G124), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n470), .B(new_n1160), .C1(new_n746), .C2(new_n766), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT120), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n762), .A2(new_n420), .ZN(new_n1163));
  INV_X1    g0963(.A(G125), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n751), .A2(new_n1164), .B1(new_n754), .B2(new_n1092), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1163), .B(new_n1165), .C1(G132), .C2(new_n779), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n823), .B2(new_n759), .C1(new_n784), .C2(new_n1089), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT59), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1158), .B(new_n1159), .C1(new_n1162), .C2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n801), .B1(new_n1169), .B2(new_n738), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(G50), .B2(new_n1107), .C1(new_n1134), .C2(new_n788), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1151), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1148), .A2(new_n1173), .ZN(G375));
  NAND2_X1  g0974(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1064), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n955), .A3(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n754), .A2(new_n823), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n751), .A2(new_n826), .B1(new_n758), .B2(new_n1089), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1178), .B(new_n1179), .C1(G128), .C2(new_n773), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n743), .A2(G159), .B1(new_n745), .B2(G58), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n830), .A2(G150), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n391), .B1(new_n763), .B2(G50), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n751), .A2(new_n771), .B1(new_n758), .B2(new_n450), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n344), .B1(new_n495), .B2(new_n759), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G303), .C2(new_n773), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n974), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n743), .A2(G97), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n755), .A2(G283), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1184), .B1(new_n1191), .B2(new_n1012), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n801), .B1(new_n1192), .B2(new_n738), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1193), .B1(new_n871), .B2(new_n788), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n213), .B2(new_n838), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(new_n1070), .B2(new_n736), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1177), .A2(new_n1196), .ZN(G381));
  INV_X1    g0997(.A(G390), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n971), .A2(new_n993), .A3(new_n1198), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1199), .A2(G396), .A3(G393), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(G375), .A2(G378), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(G381), .A2(G384), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(G407));
  INV_X1    g1003(.A(G213), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1201), .B2(new_n676), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(G407), .ZN(G409));
  XOR2_X1   g1006(.A(G393), .B(G396), .Z(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(G387), .A2(G390), .ZN(new_n1209));
  AND3_X1   g1009(.A1(new_n1209), .A2(new_n1199), .A3(KEYINPUT125), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT125), .B1(new_n1209), .B2(new_n1199), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1208), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1208), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT62), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n736), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT123), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1171), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT123), .B1(new_n1151), .B2(new_n1172), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n955), .B(new_n1111), .C1(new_n1138), .C2(new_n1143), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(G378), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1148), .A2(G378), .A3(new_n1173), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1204), .A2(G343), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT126), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(KEYINPUT126), .A3(new_n1228), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT60), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1176), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1064), .A2(new_n1069), .A3(KEYINPUT60), .A4(new_n1072), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1235), .A2(new_n1175), .A3(new_n734), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n1196), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(G384), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n845), .A3(new_n1196), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1239), .A2(KEYINPUT124), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT124), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1216), .B1(new_n1233), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1227), .A2(G2897), .ZN(new_n1247));
  MUX2_X1   g1047(.A(new_n1246), .B(new_n1243), .S(new_n1247), .Z(new_n1248));
  NAND3_X1  g1048(.A1(new_n1231), .A2(new_n1232), .A3(new_n1248), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1227), .B(new_n1243), .C1(new_n1224), .C2(new_n1225), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1250), .B2(new_n1216), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1215), .B1(new_n1245), .B2(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1233), .A2(KEYINPUT63), .A3(new_n1244), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1229), .A2(new_n1248), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT63), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n1255), .A2(new_n1256), .B1(new_n1229), .B2(new_n1243), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT61), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1254), .A2(new_n1257), .A3(new_n1258), .A4(new_n1214), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1253), .A2(new_n1259), .ZN(G405));
  NAND2_X1  g1060(.A1(new_n1225), .A2(KEYINPUT127), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G378), .B1(new_n1148), .B2(new_n1173), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1240), .B(new_n1239), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1265), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1244), .A3(new_n1263), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(new_n1215), .ZN(G402));
endmodule


