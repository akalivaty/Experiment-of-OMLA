//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n965, new_n966;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OAI221_X1 g004(.A(new_n204), .B1(KEYINPUT92), .B2(new_n205), .C1(G1gat), .C2(new_n202), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(KEYINPUT92), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n206), .B(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G71gat), .A2(G78gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(G71gat), .A2(G78gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n212), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n212), .B(new_n215), .C1(new_n210), .C2(new_n213), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n209), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G183gat), .ZN(new_n222));
  INV_X1    g021(.A(G183gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n209), .A2(new_n223), .A3(new_n220), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G231gat), .ZN(new_n226));
  INV_X1    g025(.A(G233gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n222), .A2(G231gat), .A3(G233gat), .A4(new_n224), .ZN(new_n229));
  XOR2_X1   g028(.A(G127gat), .B(G155gat), .Z(new_n230));
  XNOR2_X1  g029(.A(new_n230), .B(KEYINPUT20), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(new_n228), .B2(new_n229), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n236));
  INV_X1    g035(.A(G211gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n235), .B(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  OR3_X1    g039(.A1(new_n233), .A2(new_n234), .A3(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n233), .B2(new_n234), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G232gat), .A2(G233gat), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n244), .B(KEYINPUT97), .Z(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n246), .A2(KEYINPUT41), .ZN(new_n247));
  XOR2_X1   g046(.A(G134gat), .B(G162gat), .Z(new_n248));
  XOR2_X1   g047(.A(new_n247), .B(new_n248), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(G29gat), .ZN(new_n251));
  INV_X1    g050(.A(G36gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT14), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT14), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G29gat), .B2(G36gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G29gat), .A2(G36gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G50gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G43gat), .ZN(new_n260));
  INV_X1    g059(.A(G43gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G50gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT15), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(KEYINPUT89), .B1(new_n261), .B2(G50gat), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n267), .A2(new_n264), .B1(new_n260), .B2(new_n262), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n258), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT90), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT90), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n271), .B(new_n258), .C1(new_n266), .C2(new_n268), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n257), .A2(KEYINPUT15), .A3(new_n260), .A4(new_n262), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT17), .ZN(new_n277));
  INV_X1    g076(.A(new_n274), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(new_n270), .B2(new_n272), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G85gat), .A2(G92gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT7), .ZN(new_n284));
  OR2_X1    g083(.A1(G85gat), .A2(G92gat), .ZN(new_n285));
  INV_X1    g084(.A(G99gat), .ZN(new_n286));
  INV_X1    g085(.A(G106gat), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT8), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(new_n285), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G99gat), .B(G106gat), .Z(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n292), .A2(new_n285), .A3(new_n284), .A4(new_n288), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n282), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n246), .A2(KEYINPUT41), .ZN(new_n296));
  INV_X1    g095(.A(new_n294), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G190gat), .B(G218gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n250), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n303), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n249), .A3(new_n301), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n243), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(KEYINPUT27), .B(G183gat), .ZN(new_n309));
  INV_X1    g108(.A(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT28), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  INV_X1    g114(.A(G176gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT66), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(KEYINPUT26), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(KEYINPUT26), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n318), .B(new_n319), .C1(new_n315), .C2(new_n316), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  OR2_X1    g120(.A1(new_n314), .A2(KEYINPUT24), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n314), .A2(KEYINPUT24), .ZN(new_n323));
  NOR2_X1   g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324));
  OAI221_X1 g123(.A(new_n322), .B1(new_n315), .B2(new_n316), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n326), .A2(KEYINPUT65), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(KEYINPUT65), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n327), .A2(new_n328), .B1(G169gat), .B2(G176gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT23), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT25), .B1(new_n325), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n325), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT64), .B(G176gat), .Z(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT23), .A3(new_n315), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n333), .A2(new_n334), .A3(new_n329), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340));
  INV_X1    g139(.A(G120gat), .ZN(new_n341));
  OR2_X1    g140(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G113gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(KEYINPUT68), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT68), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G120gat), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n345), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n339), .B(new_n340), .C1(new_n344), .C2(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT1), .B1(G113gat), .B2(G120gat), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(G113gat), .B2(G120gat), .ZN(new_n352));
  OR2_X1    g151(.A1(G127gat), .A2(G134gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT67), .B(G127gat), .ZN(new_n354));
  INV_X1    g153(.A(G134gat), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n352), .B(new_n353), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G227gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(new_n227), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n357), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n321), .A2(new_n362), .A3(new_n337), .A4(new_n332), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(G71gat), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT70), .B(G99gat), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n361), .B1(new_n358), .B2(new_n363), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(KEYINPUT33), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT32), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n363), .ZN(new_n377));
  AOI221_X4 g176(.A(new_n374), .B1(KEYINPUT33), .B2(new_n371), .C1(new_n377), .C2(new_n360), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n367), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n360), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT32), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n383), .A3(new_n371), .ZN(new_n384));
  INV_X1    g183(.A(new_n378), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n366), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT88), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n379), .A2(new_n386), .A3(KEYINPUT88), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n357), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n350), .A2(KEYINPUT76), .A3(new_n356), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G155gat), .A2(G162gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT2), .ZN(new_n399));
  INV_X1    g198(.A(G155gat), .ZN(new_n400));
  INV_X1    g199(.A(G162gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n398), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n398), .B(new_n402), .C1(new_n396), .C2(KEYINPUT2), .ZN(new_n405));
  AND2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT3), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n350), .A2(new_n356), .A3(new_n405), .A4(new_n404), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT78), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT78), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n406), .A2(new_n415), .A3(new_n350), .A4(new_n356), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT4), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n418));
  AND2_X1   g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n411), .B(new_n412), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n414), .A2(new_n416), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n406), .B1(new_n393), .B2(new_n394), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(KEYINPUT5), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(G57gat), .B(G85gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G1gat), .B(G29gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT4), .ZN(new_n432));
  OAI22_X1  g231(.A1(new_n422), .A2(new_n432), .B1(new_n413), .B2(new_n418), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n411), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n425), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n425), .A2(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n430), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n438), .B(new_n440), .ZN(new_n441));
  XOR2_X1   g240(.A(G8gat), .B(G36gat), .Z(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(G92gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT75), .B(G64gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  AND2_X1   g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n338), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT22), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT74), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT74), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT22), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(G197gat), .A2(G204gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(G197gat), .A2(G204gat), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT73), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT73), .ZN(new_n456));
  INV_X1    g255(.A(G197gat), .ZN(new_n457));
  INV_X1    g256(.A(G204gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G197gat), .A2(G204gat), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n452), .B1(new_n455), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(G218gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n237), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(G211gat), .A2(G218gat), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT73), .B1(new_n453), .B2(new_n454), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n459), .A2(new_n456), .A3(new_n460), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n449), .A2(new_n451), .A3(new_n465), .ZN(new_n472));
  INV_X1    g271(.A(new_n464), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n338), .B1(KEYINPUT29), .B2(new_n446), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n447), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n447), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n445), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  INV_X1    g281(.A(new_n445), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n483), .A3(new_n478), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n484), .A3(KEYINPUT30), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT30), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n482), .A2(new_n486), .A3(new_n483), .A4(new_n478), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n441), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G50gat), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n476), .B1(new_n410), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G228gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(new_n227), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT3), .B1(new_n476), .B2(new_n493), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n495), .B(new_n497), .C1(new_n498), .C2(new_n406), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT86), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n475), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n471), .A2(new_n474), .A3(KEYINPUT84), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(new_n468), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n504), .A2(new_n505), .A3(new_n493), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n504), .B2(new_n493), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT3), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n495), .B1(new_n508), .B2(new_n406), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n497), .B(KEYINPUT83), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n500), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n471), .A2(new_n474), .A3(KEYINPUT84), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT84), .B1(new_n471), .B2(new_n474), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n466), .B1(new_n471), .B2(new_n452), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT85), .B1(new_n515), .B2(KEYINPUT29), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n504), .A2(new_n505), .A3(new_n493), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n409), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n494), .B1(new_n518), .B2(new_n407), .ZN(new_n519));
  INV_X1    g318(.A(new_n510), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n519), .A2(KEYINPUT86), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n499), .B1(new_n511), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(G22gat), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT86), .B1(new_n519), .B2(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n504), .A2(new_n493), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT3), .B1(new_n525), .B2(KEYINPUT85), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n406), .B1(new_n526), .B2(new_n517), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n500), .B(new_n510), .C1(new_n527), .C2(new_n494), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(G22gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n499), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT82), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n492), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n530), .B1(new_n529), .B2(new_n499), .ZN(new_n535));
  INV_X1    g334(.A(new_n499), .ZN(new_n536));
  AOI211_X1 g335(.A(G22gat), .B(new_n536), .C1(new_n524), .C2(new_n528), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n533), .B(new_n492), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n391), .B(new_n489), .C1(new_n534), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT35), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n533), .B1(new_n535), .B2(new_n537), .ZN(new_n542));
  INV_X1    g341(.A(new_n492), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n367), .B(new_n545), .C1(new_n376), .C2(new_n378), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n367), .A2(new_n545), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n379), .A2(new_n386), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n544), .A2(new_n538), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n439), .A2(KEYINPUT6), .A3(new_n430), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n438), .A2(KEYINPUT80), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT81), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n440), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n439), .A2(KEYINPUT81), .A3(new_n430), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n436), .A2(new_n555), .A3(new_n437), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n551), .A2(new_n553), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  AOI211_X1 g356(.A(new_n541), .B(new_n488), .C1(new_n550), .C2(new_n557), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n540), .A2(new_n541), .B1(new_n549), .B2(new_n558), .ZN(new_n559));
  OR3_X1    g358(.A1(new_n479), .A2(KEYINPUT37), .A3(new_n480), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT37), .B1(new_n479), .B2(new_n480), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n445), .A3(new_n561), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n479), .A2(new_n445), .A3(new_n480), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n562), .B1(KEYINPUT38), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n564), .B(new_n441), .C1(KEYINPUT38), .C2(new_n562), .ZN(new_n565));
  OR3_X1    g364(.A1(new_n423), .A2(new_n422), .A3(new_n421), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT39), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT87), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n433), .A2(new_n411), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(new_n421), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT87), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n566), .A2(new_n571), .A3(KEYINPUT39), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n570), .A2(KEYINPUT39), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(new_n431), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n573), .A2(KEYINPUT40), .A3(new_n574), .A4(new_n431), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n488), .A2(new_n577), .A3(new_n440), .A4(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n565), .B(new_n579), .C1(new_n534), .C2(new_n539), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n557), .A2(new_n550), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n538), .B(new_n544), .C1(new_n581), .C2(new_n488), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n387), .A2(KEYINPUT36), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n548), .A2(KEYINPUT36), .A3(new_n546), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n580), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n308), .B1(new_n559), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT93), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n206), .B(new_n207), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n275), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n209), .A2(new_n279), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n593), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n594), .B1(new_n276), .B2(new_n281), .ZN(new_n598));
  INV_X1    g397(.A(new_n595), .ZN(new_n599));
  NOR3_X1   g398(.A1(new_n598), .A2(new_n599), .A3(new_n590), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n597), .B1(new_n600), .B2(KEYINPUT18), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n282), .B2(new_n209), .ZN(new_n602));
  INV_X1    g401(.A(new_n590), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT18), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G113gat), .B(G141gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n457), .ZN(new_n608));
  XNOR2_X1  g407(.A(KEYINPUT11), .B(G169gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT12), .Z(new_n611));
  OAI211_X1 g410(.A(new_n601), .B(new_n606), .C1(KEYINPUT94), .C2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT17), .B1(new_n275), .B2(KEYINPUT91), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n279), .A2(new_n280), .A3(new_n277), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n209), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n615), .A2(KEYINPUT18), .A3(new_n595), .A4(new_n603), .ZN(new_n616));
  INV_X1    g415(.A(new_n597), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(KEYINPUT94), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n611), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n616), .A2(new_n617), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT18), .B1(new_n602), .B2(new_n603), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n612), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT98), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n294), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT98), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT98), .B1(new_n217), .B2(new_n218), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n625), .B(new_n626), .C1(new_n629), .C2(new_n294), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n297), .A2(KEYINPUT10), .A3(new_n219), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n625), .B1(new_n629), .B2(new_n294), .ZN(new_n635));
  INV_X1    g434(.A(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT99), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n639), .A3(new_n636), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n634), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n634), .A2(new_n638), .A3(new_n646), .A4(new_n640), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n623), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n588), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n581), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g451(.A1(new_n540), .A2(new_n541), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n549), .A2(new_n558), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n587), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n243), .A2(new_n307), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n655), .A2(new_n649), .A3(new_n488), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT100), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n588), .A2(new_n659), .A3(new_n649), .A4(new_n488), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n658), .A2(G8gat), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n658), .A2(new_n660), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT16), .B(G8gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n650), .A2(KEYINPUT42), .A3(new_n488), .A4(new_n666), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n663), .A2(new_n669), .A3(new_n670), .ZN(G1325gat));
  AOI21_X1  g470(.A(G15gat), .B1(new_n650), .B2(new_n391), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n586), .A2(KEYINPUT103), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n583), .A2(KEYINPUT103), .A3(new_n584), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n676), .A2(G15gat), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n672), .B1(new_n650), .B2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n534), .A2(new_n539), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n650), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(G22gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n650), .A2(new_n530), .A3(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n683), .B(new_n685), .ZN(G1327gat));
  AOI21_X1  g485(.A(new_n307), .B1(new_n559), .B2(new_n587), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n243), .A2(new_n623), .A3(new_n648), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n251), .A3(new_n581), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  INV_X1    g490(.A(new_n307), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n655), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n688), .ZN(new_n697));
  INV_X1    g496(.A(new_n581), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n691), .A2(new_n699), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n689), .A2(new_n252), .A3(new_n488), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n702));
  INV_X1    g501(.A(new_n488), .ZN(new_n703));
  OAI21_X1  g502(.A(G36gat), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n701), .A2(KEYINPUT46), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n705), .A2(KEYINPUT105), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n701), .A2(new_n707), .A3(KEYINPUT46), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n702), .B(new_n704), .C1(new_n706), .C2(new_n708), .ZN(G1329gat));
  OAI21_X1  g508(.A(G43gat), .B1(new_n697), .B2(new_n586), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n689), .A2(new_n261), .A3(new_n391), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT47), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G43gat), .B1(new_n697), .B2(new_n675), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n713), .A2(new_n711), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT48), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n687), .A2(new_n679), .A3(new_n688), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n259), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n679), .A2(G50gat), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n717), .B(new_n719), .C1(new_n697), .C2(new_n720), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n716), .A2(KEYINPUT48), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(G1331gat));
  INV_X1    g522(.A(new_n623), .ZN(new_n724));
  INV_X1    g523(.A(new_n648), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n655), .A2(new_n656), .A3(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n698), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g528(.A(KEYINPUT49), .B(G64gat), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n588), .A2(KEYINPUT107), .A3(new_n726), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT107), .B1(new_n588), .B2(new_n726), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n488), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n588), .A2(KEYINPUT107), .A3(new_n726), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n703), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n733), .B(new_n734), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n488), .B1(new_n731), .B2(new_n732), .ZN(new_n742));
  INV_X1    g541(.A(new_n739), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n734), .B1(new_n744), .B2(new_n733), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n741), .A2(new_n745), .ZN(G1333gat));
  INV_X1    g545(.A(G71gat), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n588), .A2(new_n747), .A3(new_n391), .A4(new_n726), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n675), .B1(new_n736), .B2(new_n737), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n747), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1334gat));
  OAI21_X1  g551(.A(new_n679), .B1(new_n731), .B2(new_n732), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  INV_X1    g553(.A(new_n243), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n623), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT110), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(new_n648), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n695), .A2(new_n696), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n698), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n698), .A2(G85gat), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n687), .A2(KEYINPUT51), .A3(new_n757), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n687), .B2(new_n757), .ZN(new_n763));
  OAI211_X1 g562(.A(new_n648), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n760), .A2(KEYINPUT111), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(G1336gat));
  NAND4_X1  g568(.A1(new_n695), .A2(new_n488), .A3(new_n696), .A4(new_n758), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G92gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT112), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n703), .A2(G92gat), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n648), .B(new_n773), .C1(new_n762), .C2(new_n763), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n772), .A2(new_n775), .A3(KEYINPUT52), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n771), .B(new_n774), .C1(KEYINPUT112), .C2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n759), .B2(new_n675), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n391), .A2(new_n286), .A3(new_n648), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT113), .Z(new_n782));
  OAI21_X1  g581(.A(new_n782), .B1(new_n762), .B2(new_n763), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT114), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n780), .A2(new_n786), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1338gat));
  OR2_X1    g587(.A1(new_n762), .A2(new_n763), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n679), .A2(new_n287), .A3(new_n648), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT115), .Z(new_n791));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n695), .A2(new_n679), .A3(new_n696), .A4(new_n758), .ZN(new_n794));
  AOI22_X1  g593(.A1(new_n789), .A2(new_n793), .B1(new_n794), .B2(G106gat), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n794), .A2(G106gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n791), .B1(new_n762), .B2(new_n763), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n796), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n795), .A2(new_n796), .B1(new_n797), .B2(new_n799), .ZN(G1339gat));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801));
  INV_X1    g600(.A(new_n610), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n603), .B1(new_n615), .B2(new_n595), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n595), .A2(new_n596), .A3(new_n593), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n611), .B1(new_n600), .B2(KEYINPUT18), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n648), .B(new_n805), .C1(new_n806), .C2(new_n620), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT117), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n601), .A2(new_n606), .A3(new_n611), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n648), .A4(new_n805), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n630), .A2(new_n636), .A3(new_n631), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n634), .A2(KEYINPUT54), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n636), .B1(new_n630), .B2(new_n631), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n646), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n647), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n612), .B2(new_n622), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n307), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n805), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n307), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n243), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n308), .A2(new_n648), .A3(new_n724), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n801), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n656), .A2(new_n725), .A3(new_n623), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n307), .A2(new_n822), .A3(new_n825), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n808), .B(new_n811), .C1(new_n623), .C2(new_n822), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n307), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT118), .B(new_n830), .C1(new_n833), .C2(new_n243), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n679), .B1(new_n390), .B2(new_n389), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n698), .A2(new_n488), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n829), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT119), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(new_n724), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n829), .A2(new_n834), .A3(new_n549), .A4(new_n836), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT120), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n342), .A2(new_n343), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n724), .A2(new_n846), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n839), .A2(new_n345), .B1(new_n845), .B2(new_n847), .ZN(G1340gat));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n341), .B1(new_n838), .B2(new_n648), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n346), .A2(new_n348), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n648), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT121), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n844), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n849), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n837), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n837), .A2(new_n857), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n648), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G120gat), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT122), .A3(new_n854), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n856), .A2(new_n862), .ZN(G1341gat));
  NOR2_X1   g662(.A1(new_n840), .A2(new_n755), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n755), .A2(new_n354), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n866), .A2(new_n354), .B1(new_n838), .B2(new_n867), .ZN(G1342gat));
  NOR3_X1   g667(.A1(new_n840), .A2(G134gat), .A3(new_n307), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n838), .A2(new_n692), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n871), .B(new_n872), .C1(new_n873), .C2(new_n355), .ZN(G1343gat));
  AND2_X1   g673(.A1(new_n829), .A2(new_n834), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n836), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n623), .A2(G141gat), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(new_n679), .A3(new_n675), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n836), .A2(new_n586), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n829), .A2(new_n834), .A3(new_n679), .ZN(new_n880));
  XNOR2_X1  g679(.A(KEYINPUT124), .B(KEYINPUT57), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n807), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n307), .B1(new_n823), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n243), .B1(new_n826), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n679), .B1(new_n886), .B2(new_n828), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n623), .B(new_n879), .C1(new_n883), .C2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(G141gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n878), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT58), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n878), .B(new_n894), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(G1344gat));
  AND3_X1   g695(.A1(new_n876), .A2(new_n679), .A3(new_n675), .ZN(new_n897));
  INV_X1    g696(.A(G148gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n897), .A2(new_n898), .A3(new_n648), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n879), .B1(new_n883), .B2(new_n889), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT59), .B(new_n898), .C1(new_n900), .C2(new_n648), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n829), .A2(new_n834), .A3(new_n679), .A4(new_n881), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n905), .A2(new_n648), .A3(new_n586), .A4(new_n836), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n906), .B2(G148gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n899), .B1(new_n901), .B2(new_n907), .ZN(G1345gat));
  AOI21_X1  g707(.A(G155gat), .B1(new_n897), .B2(new_n243), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n755), .A2(new_n400), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n909), .B1(new_n900), .B2(new_n910), .ZN(G1346gat));
  AOI21_X1  g710(.A(G162gat), .B1(new_n897), .B2(new_n692), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n307), .A2(new_n401), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n900), .B2(new_n913), .ZN(G1347gat));
  AND2_X1   g713(.A1(new_n875), .A2(new_n698), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n915), .A2(new_n488), .A3(new_n549), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n315), .A3(new_n724), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n875), .A2(new_n698), .A3(new_n835), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n623), .A3(new_n703), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n917), .B1(new_n315), .B2(new_n919), .ZN(G1348gat));
  AOI21_X1  g719(.A(G176gat), .B1(new_n916), .B2(new_n648), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n918), .A2(new_n703), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n725), .A2(new_n335), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1349gat));
  AND2_X1   g723(.A1(new_n243), .A2(new_n309), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n915), .A2(new_n488), .A3(new_n549), .A4(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n918), .A2(new_n703), .A3(new_n755), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n927), .B2(new_n223), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n926), .B(new_n930), .C1(new_n927), .C2(new_n223), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1350gat));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n310), .A3(new_n692), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n915), .A2(new_n488), .A3(new_n835), .A4(new_n692), .ZN(new_n934));
  XNOR2_X1  g733(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n934), .A2(G190gat), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n934), .B2(G190gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  NOR3_X1   g737(.A1(new_n673), .A2(new_n703), .A3(new_n674), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(KEYINPUT126), .A3(new_n679), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n875), .A2(new_n940), .A3(new_n698), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT126), .B1(new_n939), .B2(new_n679), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n457), .A3(new_n724), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n698), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n945), .B1(new_n903), .B2(new_n904), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n623), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(new_n948), .ZN(G1352gat));
  NAND3_X1  g748(.A1(new_n943), .A2(new_n458), .A3(new_n648), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT62), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n953));
  NOR4_X1   g752(.A1(new_n941), .A2(G204gat), .A3(new_n725), .A4(new_n942), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n951), .A2(KEYINPUT62), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n905), .A2(new_n648), .ZN(new_n957));
  OAI21_X1  g756(.A(G204gat), .B1(new_n957), .B2(new_n945), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n952), .A2(new_n956), .A3(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n237), .A3(new_n243), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n946), .A2(new_n243), .ZN(new_n961));
  AND3_X1   g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  AOI21_X1  g761(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(G1354gat));
  NAND3_X1  g763(.A1(new_n943), .A2(new_n463), .A3(new_n692), .ZN(new_n965));
  OAI21_X1  g764(.A(G218gat), .B1(new_n947), .B2(new_n307), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(new_n966), .ZN(G1355gat));
endmodule


