

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U321 ( .A(KEYINPUT66), .B(n415), .Z(n289) );
  INV_X1 U322 ( .A(KEYINPUT113), .ZN(n409) );
  XNOR2_X1 U323 ( .A(n450), .B(KEYINPUT123), .ZN(n581) );
  XOR2_X1 U324 ( .A(n548), .B(KEYINPUT28), .Z(n524) );
  XNOR2_X1 U325 ( .A(n452), .B(G218GAT), .ZN(n453) );
  XNOR2_X1 U326 ( .A(n454), .B(n453), .ZN(G1355GAT) );
  XOR2_X1 U327 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n291) );
  XNOR2_X1 U328 ( .A(KEYINPUT78), .B(KEYINPUT9), .ZN(n290) );
  XNOR2_X1 U329 ( .A(n291), .B(n290), .ZN(n312) );
  INV_X1 U330 ( .A(KEYINPUT8), .ZN(n292) );
  NAND2_X1 U331 ( .A1(G36GAT), .A2(n292), .ZN(n295) );
  INV_X1 U332 ( .A(G36GAT), .ZN(n293) );
  NAND2_X1 U333 ( .A1(n293), .A2(KEYINPUT8), .ZN(n294) );
  NAND2_X1 U334 ( .A1(n295), .A2(n294), .ZN(n297) );
  XNOR2_X1 U335 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n296) );
  XNOR2_X1 U336 ( .A(n297), .B(n296), .ZN(n415) );
  NAND2_X1 U337 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U338 ( .A(n289), .B(n298), .ZN(n302) );
  XOR2_X1 U339 ( .A(G162GAT), .B(G50GAT), .Z(n321) );
  XOR2_X1 U340 ( .A(G134GAT), .B(G43GAT), .Z(n342) );
  XNOR2_X1 U341 ( .A(n321), .B(n342), .ZN(n300) );
  XNOR2_X1 U342 ( .A(G85GAT), .B(KEYINPUT73), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n299), .B(G92GAT), .ZN(n378) );
  XNOR2_X1 U344 ( .A(n300), .B(n378), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n310) );
  XOR2_X1 U346 ( .A(G106GAT), .B(G190GAT), .Z(n304) );
  XNOR2_X1 U347 ( .A(G218GAT), .B(KEYINPUT65), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U349 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n306) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(KEYINPUT11), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U352 ( .A(n308), .B(n307), .Z(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X2 U354 ( .A(n312), .B(n311), .Z(n567) );
  XNOR2_X1 U355 ( .A(n567), .B(KEYINPUT104), .ZN(n313) );
  XNOR2_X1 U356 ( .A(n313), .B(KEYINPUT36), .ZN(n486) );
  XNOR2_X1 U357 ( .A(KEYINPUT97), .B(KEYINPUT26), .ZN(n356) );
  XOR2_X1 U358 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n315) );
  XNOR2_X1 U359 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U361 ( .A(n316), .B(KEYINPUT88), .Z(n318) );
  XOR2_X1 U362 ( .A(G155GAT), .B(G22GAT), .Z(n392) );
  XNOR2_X1 U363 ( .A(n392), .B(KEYINPUT23), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n318), .B(n317), .ZN(n325) );
  XOR2_X1 U365 ( .A(G141GAT), .B(KEYINPUT2), .Z(n320) );
  XNOR2_X1 U366 ( .A(KEYINPUT3), .B(KEYINPUT91), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n370) );
  XOR2_X1 U368 ( .A(n321), .B(n370), .Z(n323) );
  NAND2_X1 U369 ( .A1(G228GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U371 ( .A(n325), .B(n324), .Z(n335) );
  XNOR2_X1 U372 ( .A(G197GAT), .B(KEYINPUT90), .ZN(n326) );
  XNOR2_X1 U373 ( .A(n326), .B(KEYINPUT21), .ZN(n327) );
  XOR2_X1 U374 ( .A(n327), .B(KEYINPUT89), .Z(n329) );
  XNOR2_X1 U375 ( .A(G218GAT), .B(G211GAT), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n329), .B(n328), .ZN(n445) );
  XNOR2_X1 U377 ( .A(G78GAT), .B(KEYINPUT72), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n330), .B(KEYINPUT71), .ZN(n331) );
  XOR2_X1 U379 ( .A(n331), .B(G204GAT), .Z(n333) );
  XNOR2_X1 U380 ( .A(G148GAT), .B(G106GAT), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n390) );
  XNOR2_X1 U382 ( .A(n445), .B(n390), .ZN(n334) );
  XNOR2_X1 U383 ( .A(n335), .B(n334), .ZN(n548) );
  XOR2_X1 U384 ( .A(KEYINPUT64), .B(KEYINPUT82), .Z(n341) );
  XOR2_X1 U385 ( .A(KEYINPUT85), .B(KEYINPUT81), .Z(n337) );
  XNOR2_X1 U386 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n336) );
  XNOR2_X1 U387 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U388 ( .A(G120GAT), .B(G99GAT), .ZN(n338) );
  XNOR2_X1 U389 ( .A(n338), .B(G71GAT), .ZN(n386) );
  XNOR2_X1 U390 ( .A(n339), .B(n386), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n346) );
  XOR2_X1 U392 ( .A(G113GAT), .B(G15GAT), .Z(n413) );
  XOR2_X1 U393 ( .A(n413), .B(n342), .Z(n344) );
  NAND2_X1 U394 ( .A1(G227GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U396 ( .A(n346), .B(n345), .Z(n354) );
  XOR2_X1 U397 ( .A(KEYINPUT0), .B(G127GAT), .Z(n371) );
  XOR2_X1 U398 ( .A(G169GAT), .B(G176GAT), .Z(n348) );
  XNOR2_X1 U399 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U401 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n350) );
  XNOR2_X1 U402 ( .A(G190GAT), .B(KEYINPUT84), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U404 ( .A(n352), .B(n351), .Z(n444) );
  XNOR2_X1 U405 ( .A(n371), .B(n444), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n553) );
  NOR2_X1 U407 ( .A1(n548), .A2(n553), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n356), .B(n355), .ZN(n460) );
  INV_X1 U409 ( .A(n460), .ZN(n538) );
  XOR2_X1 U410 ( .A(G148GAT), .B(G155GAT), .Z(n358) );
  XNOR2_X1 U411 ( .A(G134GAT), .B(G85GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U413 ( .A(G57GAT), .B(G1GAT), .Z(n360) );
  XNOR2_X1 U414 ( .A(G120GAT), .B(G113GAT), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U416 ( .A(n362), .B(n361), .Z(n367) );
  XOR2_X1 U417 ( .A(KEYINPUT6), .B(KEYINPUT94), .Z(n364) );
  NAND2_X1 U418 ( .A1(G225GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U420 ( .A(KEYINPUT95), .B(n365), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n377) );
  XOR2_X1 U422 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n369) );
  XNOR2_X1 U423 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n375) );
  XOR2_X1 U425 ( .A(n371), .B(n370), .Z(n373) );
  XNOR2_X1 U426 ( .A(G29GAT), .B(G162GAT), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U428 ( .A(n375), .B(n374), .Z(n376) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n512) );
  XOR2_X1 U430 ( .A(KEYINPUT31), .B(n378), .Z(n380) );
  NAND2_X1 U431 ( .A1(G230GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U433 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n382) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(KEYINPUT70), .ZN(n381) );
  XNOR2_X1 U435 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U436 ( .A(n384), .B(n383), .Z(n388) );
  XNOR2_X1 U437 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n385) );
  XNOR2_X1 U438 ( .A(n385), .B(G64GAT), .ZN(n391) );
  XNOR2_X1 U439 ( .A(n391), .B(n386), .ZN(n387) );
  XNOR2_X1 U440 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n390), .B(n389), .ZN(n577) );
  INV_X1 U442 ( .A(KEYINPUT45), .ZN(n407) );
  XOR2_X1 U443 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U444 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U445 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U446 ( .A(G1GAT), .B(G8GAT), .Z(n416) );
  XOR2_X1 U447 ( .A(n395), .B(n416), .Z(n397) );
  XNOR2_X1 U448 ( .A(G78GAT), .B(G211GAT), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n397), .B(n396), .ZN(n405) );
  XOR2_X1 U450 ( .A(G15GAT), .B(G71GAT), .Z(n399) );
  XNOR2_X1 U451 ( .A(G127GAT), .B(G183GAT), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n401) );
  XNOR2_X1 U454 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U456 ( .A(n403), .B(n402), .Z(n404) );
  XNOR2_X1 U457 ( .A(n405), .B(n404), .ZN(n564) );
  NOR2_X1 U458 ( .A1(n486), .A2(n564), .ZN(n406) );
  XNOR2_X1 U459 ( .A(n407), .B(n406), .ZN(n408) );
  NOR2_X1 U460 ( .A1(n577), .A2(n408), .ZN(n410) );
  XNOR2_X1 U461 ( .A(n410), .B(n409), .ZN(n428) );
  XOR2_X1 U462 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n412) );
  XNOR2_X1 U463 ( .A(G197GAT), .B(G169GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U465 ( .A(n414), .B(n413), .Z(n418) );
  XNOR2_X1 U466 ( .A(n415), .B(n416), .ZN(n417) );
  XNOR2_X1 U467 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U468 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n420) );
  NAND2_X1 U469 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U470 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U471 ( .A(n422), .B(n421), .Z(n427) );
  XOR2_X1 U472 ( .A(G22GAT), .B(G43GAT), .Z(n424) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(G50GAT), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U475 ( .A(n425), .B(KEYINPUT67), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n427), .B(n426), .ZN(n555) );
  NAND2_X1 U477 ( .A1(n428), .A2(n555), .ZN(n436) );
  XNOR2_X1 U478 ( .A(KEYINPUT112), .B(KEYINPUT47), .ZN(n434) );
  NAND2_X1 U479 ( .A1(n567), .A2(n564), .ZN(n432) );
  XNOR2_X1 U480 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n430) );
  XNOR2_X1 U481 ( .A(KEYINPUT41), .B(n577), .ZN(n559) );
  NOR2_X1 U482 ( .A1(n555), .A2(n559), .ZN(n429) );
  XOR2_X1 U483 ( .A(n430), .B(n429), .Z(n431) );
  NOR2_X1 U484 ( .A1(n432), .A2(n431), .ZN(n433) );
  XNOR2_X1 U485 ( .A(n434), .B(n433), .ZN(n435) );
  NAND2_X1 U486 ( .A1(n436), .A2(n435), .ZN(n437) );
  XNOR2_X1 U487 ( .A(n437), .B(KEYINPUT48), .ZN(n521) );
  XOR2_X1 U488 ( .A(KEYINPUT96), .B(G204GAT), .Z(n439) );
  XNOR2_X1 U489 ( .A(G8GAT), .B(G64GAT), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U491 ( .A(G92GAT), .B(G36GAT), .Z(n441) );
  NAND2_X1 U492 ( .A1(G226GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U494 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U495 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U496 ( .A(n447), .B(n446), .ZN(n514) );
  NAND2_X1 U497 ( .A1(n521), .A2(n514), .ZN(n448) );
  XNOR2_X1 U498 ( .A(n448), .B(KEYINPUT54), .ZN(n551) );
  NOR2_X1 U499 ( .A1(n512), .A2(n551), .ZN(n449) );
  NAND2_X1 U500 ( .A1(n538), .A2(n449), .ZN(n450) );
  INV_X1 U501 ( .A(n581), .ZN(n451) );
  NOR2_X1 U502 ( .A1(n486), .A2(n451), .ZN(n454) );
  XNOR2_X1 U503 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n452) );
  XOR2_X1 U504 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n476) );
  NOR2_X1 U505 ( .A1(n555), .A2(n577), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT74), .B(n455), .Z(n488) );
  NAND2_X1 U507 ( .A1(n514), .A2(n553), .ZN(n456) );
  XNOR2_X1 U508 ( .A(KEYINPUT98), .B(n456), .ZN(n457) );
  NAND2_X1 U509 ( .A1(n457), .A2(n548), .ZN(n459) );
  XOR2_X1 U510 ( .A(KEYINPUT25), .B(KEYINPUT99), .Z(n458) );
  XNOR2_X1 U511 ( .A(n459), .B(n458), .ZN(n462) );
  XOR2_X1 U512 ( .A(n514), .B(KEYINPUT27), .Z(n467) );
  NOR2_X1 U513 ( .A1(n467), .A2(n460), .ZN(n461) );
  NOR2_X1 U514 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n463), .B(KEYINPUT100), .ZN(n464) );
  NOR2_X1 U516 ( .A1(n512), .A2(n464), .ZN(n465) );
  XNOR2_X1 U517 ( .A(n465), .B(KEYINPUT101), .ZN(n470) );
  XNOR2_X1 U518 ( .A(KEYINPUT86), .B(n553), .ZN(n466) );
  NOR2_X1 U519 ( .A1(n524), .A2(n466), .ZN(n468) );
  INV_X1 U520 ( .A(n512), .ZN(n549) );
  NOR2_X1 U521 ( .A1(n549), .A2(n467), .ZN(n520) );
  NAND2_X1 U522 ( .A1(n468), .A2(n520), .ZN(n469) );
  NAND2_X1 U523 ( .A1(n470), .A2(n469), .ZN(n483) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n472) );
  INV_X1 U525 ( .A(n564), .ZN(n580) );
  NAND2_X1 U526 ( .A1(n580), .A2(n567), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U528 ( .A1(n483), .A2(n473), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT102), .ZN(n500) );
  NOR2_X1 U530 ( .A1(n488), .A2(n500), .ZN(n481) );
  NAND2_X1 U531 ( .A1(n481), .A2(n512), .ZN(n475) );
  XNOR2_X1 U532 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n481), .A2(n514), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U537 ( .A1(n481), .A2(n553), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U539 ( .A1(n481), .A2(n524), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U541 ( .A(G29GAT), .B(KEYINPUT39), .Z(n491) );
  NAND2_X1 U542 ( .A1(n564), .A2(n483), .ZN(n484) );
  XOR2_X1 U543 ( .A(KEYINPUT105), .B(n484), .Z(n485) );
  NOR2_X1 U544 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U545 ( .A(KEYINPUT37), .B(n487), .ZN(n510) );
  NOR2_X1 U546 ( .A1(n510), .A2(n488), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n489), .B(KEYINPUT38), .ZN(n496) );
  NAND2_X1 U548 ( .A1(n496), .A2(n512), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U550 ( .A1(n496), .A2(n514), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT106), .ZN(n493) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n496), .A2(n553), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT40), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  XOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT107), .Z(n498) );
  NAND2_X1 U557 ( .A1(n524), .A2(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  INV_X1 U559 ( .A(n555), .ZN(n574) );
  NOR2_X1 U560 ( .A1(n559), .A2(n574), .ZN(n499) );
  XOR2_X1 U561 ( .A(KEYINPUT108), .B(n499), .Z(n511) );
  NOR2_X1 U562 ( .A1(n511), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(KEYINPUT109), .B(n501), .Z(n506) );
  NAND2_X1 U564 ( .A1(n512), .A2(n506), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(KEYINPUT42), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NAND2_X1 U567 ( .A1(n506), .A2(n514), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n504), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U569 ( .A1(n506), .A2(n553), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n508) );
  NAND2_X1 U572 ( .A1(n506), .A2(n524), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U575 ( .A1(n511), .A2(n510), .ZN(n517) );
  NAND2_X1 U576 ( .A1(n512), .A2(n517), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U578 ( .A1(n517), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n553), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n524), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n518), .B(KEYINPUT44), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n522), .Z(n537) );
  NAND2_X1 U587 ( .A1(n553), .A2(n537), .ZN(n523) );
  NOR2_X1 U588 ( .A1(n524), .A2(n523), .ZN(n533) );
  NAND2_X1 U589 ( .A1(n533), .A2(n574), .ZN(n525) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n528) );
  INV_X1 U592 ( .A(n559), .ZN(n526) );
  NAND2_X1 U593 ( .A1(n533), .A2(n526), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(G120GAT), .B(n529), .Z(G1341GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n580), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n535) );
  INV_X1 U600 ( .A(n567), .ZN(n532) );
  NAND2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(n536), .ZN(G1343GAT) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n555), .A2(n545), .ZN(n539) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n539), .Z(G1344GAT) );
  NOR2_X1 U607 ( .A1(n559), .A2(n545), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n542), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n564), .A2(n545), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n567), .A2(n545), .ZN(n546) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(n546), .Z(n547) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n547), .ZN(G1347GAT) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT55), .B(n552), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n566) );
  NOR2_X1 U621 ( .A1(n555), .A2(n566), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n558), .ZN(G1348GAT) );
  NOR2_X1 U625 ( .A1(n566), .A2(n559), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NOR2_X1 U630 ( .A1(n564), .A2(n566), .ZN(n565) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n565), .Z(G1350GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(G190GAT), .B(n570), .Z(G1351GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(n573), .Z(n576) );
  NAND2_X1 U640 ( .A1(n581), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U643 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(KEYINPUT126), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n583), .ZN(G1354GAT) );
endmodule

