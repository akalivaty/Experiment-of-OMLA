//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n463), .A2(new_n465), .A3(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(KEYINPUT66), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n467), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n463), .A2(new_n465), .A3(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G101), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n469), .B1(new_n476), .B2(KEYINPUT66), .ZN(G160));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n463), .A2(new_n465), .A3(new_n461), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT67), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OR3_X1    g063(.A1(new_n486), .A2(KEYINPUT67), .A3(new_n487), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n482), .A2(new_n484), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n478), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n462), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n498), .B(new_n499), .C1(G102), .C2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(new_n461), .B2(G114), .ZN(new_n501));
  NOR2_X1   g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT70), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n485), .A2(KEYINPUT72), .A3(new_n506), .A4(G138), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n461), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n509), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n505), .B1(new_n511), .B2(new_n516), .ZN(G164));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT6), .A2(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G50), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n526), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n522), .A2(G62), .ZN(new_n532));
  NAND2_X1  g107(.A1(G75), .A2(G543), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT73), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n530), .A2(new_n535), .ZN(G166));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n523), .A2(new_n524), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n518), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n540), .A2(new_n522), .B1(new_n541), .B2(G51), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n526), .A2(new_n547), .B1(new_n528), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n531), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n549), .A2(new_n551), .ZN(G171));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  INV_X1    g128(.A(G43), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n526), .A2(new_n553), .B1(new_n528), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n556), .A2(new_n531), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT74), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n568));
  NOR2_X1   g143(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n566), .B1(new_n541), .B2(G53), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(KEYINPUT76), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n522), .A2(KEYINPUT77), .ZN(new_n576));
  INV_X1    g151(.A(G65), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n519), .A2(new_n521), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR3_X1   g155(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G78), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n518), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT76), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n585), .B1(new_n571), .B2(new_n573), .ZN(new_n586));
  INV_X1    g161(.A(new_n526), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G91), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n575), .A2(new_n584), .A3(new_n586), .A4(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  INV_X1    g165(.A(G166), .ZN(G303));
  NAND2_X1  g166(.A1(new_n541), .A2(G49), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT78), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n522), .A2(G74), .ZN(new_n594));
  AOI22_X1  g169(.A1(G87), .A2(new_n587), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(G288));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  INV_X1    g172(.A(G48), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n526), .A2(new_n597), .B1(new_n528), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n522), .A2(G61), .ZN(new_n600));
  NAND2_X1  g175(.A1(G73), .A2(G543), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT79), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n531), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n599), .A2(new_n603), .ZN(G305));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  INV_X1    g180(.A(G47), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n526), .A2(new_n605), .B1(new_n528), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n531), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(G290));
  NAND2_X1  g186(.A1(G301), .A2(G868), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n578), .B(new_n579), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT80), .B(G66), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G79), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(new_n518), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT81), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n619));
  OAI221_X1 g194(.A(new_n619), .B1(new_n616), .B2(new_n518), .C1(new_n613), .C2(new_n614), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n618), .A2(new_n620), .A3(G651), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n587), .A2(G92), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT10), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n541), .A2(G54), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n621), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n612), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n612), .B1(new_n626), .B2(G868), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  XNOR2_X1  g204(.A(G299), .B(KEYINPUT82), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G280));
  XOR2_X1   g206(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  AND2_X1   g209(.A1(new_n621), .A2(new_n624), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n635), .A2(new_n633), .A3(new_n623), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G868), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g213(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g214(.A1(new_n485), .A2(G135), .ZN(new_n640));
  OR2_X1    g215(.A1(G99), .A2(G2105), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n641), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n479), .B(KEYINPUT68), .ZN(new_n643));
  INV_X1    g218(.A(G123), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n640), .B(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT84), .ZN(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT12), .Z(new_n650));
  XOR2_X1   g225(.A(KEYINPUT13), .B(G2100), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  XOR2_X1   g230(.A(G2427), .B(G2430), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT16), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1341), .B(G1348), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT86), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2067), .B(G2678), .Z(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT87), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  NOR2_X1   g249(.A1(G2072), .A2(G2078), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n443), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT89), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n673), .B(new_n678), .C1(new_n677), .C2(new_n676), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n671), .B(new_n674), .C1(new_n443), .C2(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n672), .B(new_n674), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n676), .B(KEYINPUT17), .Z(new_n683));
  OAI211_X1 g258(.A(new_n679), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n647), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(G2100), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G227));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT20), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n691), .A2(new_n693), .A3(new_n695), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n698), .B(new_n699), .C1(new_n697), .C2(new_n696), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1991), .B(G1996), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1981), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n702), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT90), .B(G1986), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(G229));
  NAND2_X1  g282(.A1(new_n485), .A2(G131), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT92), .Z(new_n709));
  NAND2_X1  g284(.A1(new_n481), .A2(G119), .ZN(new_n710));
  OR2_X1    g285(.A1(G95), .A2(G2105), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n711), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G25), .ZN(new_n717));
  OAI21_X1  g292(.A(KEYINPUT91), .B1(new_n717), .B2(G29), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n717), .A2(KEYINPUT91), .A3(G29), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G24), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n610), .B2(new_n723), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT94), .B(G1986), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n725), .B(new_n726), .Z(new_n727));
  NOR2_X1   g302(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G16), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(G288), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT33), .B(G1976), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n723), .A2(G6), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n599), .A2(new_n603), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(new_n723), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT32), .B(G1981), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G22), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G166), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1971), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n733), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n728), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n745), .A2(KEYINPUT96), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n728), .A2(new_n746), .A3(new_n744), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n750), .C1(new_n746), .C2(new_n745), .ZN(new_n751));
  NAND2_X1  g326(.A1(G168), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G16), .B2(G21), .ZN(new_n753));
  INV_X1    g328(.A(G1966), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT106), .Z(new_n756));
  XOR2_X1   g331(.A(KEYINPUT31), .B(G11), .Z(new_n757));
  INV_X1    g332(.A(G29), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT30), .B(G28), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n646), .B2(new_n758), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n753), .A2(new_n754), .ZN(new_n763));
  NOR2_X1   g338(.A1(G5), .A2(G16), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G171), .B2(G16), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G1961), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n762), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(KEYINPUT107), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(KEYINPUT107), .ZN(new_n769));
  NOR2_X1   g344(.A1(G27), .A2(G29), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G164), .B2(G29), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n769), .C1(G2078), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n758), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n758), .ZN(new_n774));
  MUX2_X1   g349(.A(new_n773), .B(new_n774), .S(KEYINPUT108), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT29), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n758), .A2(G33), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n485), .A2(G139), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT102), .B(KEYINPUT25), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n478), .A2(G127), .ZN(new_n783));
  INV_X1    g358(.A(G115), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n462), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n779), .B(new_n782), .C1(G2105), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(new_n758), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT103), .Z(new_n788));
  AOI22_X1  g363(.A1(new_n788), .A2(G2072), .B1(G2078), .B2(new_n771), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT100), .B(KEYINPUT28), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT101), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n758), .A2(G26), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n791), .B(new_n792), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n485), .A2(G140), .ZN(new_n794));
  NOR2_X1   g369(.A1(G104), .A2(G2105), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n796));
  INV_X1    g371(.A(G128), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n794), .B1(new_n795), .B2(new_n796), .C1(new_n643), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT99), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n793), .B1(new_n799), .B2(G29), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G2067), .ZN(new_n801));
  NOR2_X1   g376(.A1(G4), .A2(G16), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n626), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT97), .B(G1348), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n803), .B(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n777), .A2(new_n789), .A3(new_n801), .A4(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(G29), .A2(G32), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n481), .A2(G129), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n485), .A2(G141), .ZN(new_n811));
  NAND3_X1  g386(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT26), .Z(new_n813));
  NAND4_X1  g388(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n758), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT27), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1996), .ZN(new_n817));
  INV_X1    g392(.A(G1961), .ZN(new_n818));
  INV_X1    g393(.A(new_n765), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n723), .A2(KEYINPUT23), .A3(G20), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT23), .ZN(new_n822));
  INV_X1    g397(.A(G20), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G16), .ZN(new_n824));
  INV_X1    g399(.A(G299), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n821), .B(new_n824), .C1(new_n825), .C2(new_n723), .ZN(new_n826));
  INV_X1    g401(.A(G1956), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n820), .B(new_n828), .C1(G2090), .C2(new_n776), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n772), .A2(new_n807), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(G16), .A2(G19), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n558), .B2(G16), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT98), .B(G1341), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT24), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n758), .B1(new_n835), .B2(G34), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT105), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n835), .A2(G34), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n837), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT66), .B1(new_n468), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT66), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n471), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n841), .B1(new_n846), .B2(new_n758), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G2084), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n751), .A2(new_n830), .A3(new_n834), .A4(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n788), .A2(G2072), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT104), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n849), .A2(new_n851), .ZN(G311));
  AND2_X1   g427(.A1(new_n751), .A2(new_n830), .ZN(new_n853));
  INV_X1    g428(.A(new_n851), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n853), .A2(new_n854), .A3(new_n834), .A4(new_n848), .ZN(G150));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n526), .A2(new_n856), .B1(new_n528), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(new_n531), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n558), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n861), .B1(new_n557), .B2(new_n555), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n625), .A2(new_n633), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n864), .B1(new_n871), .B2(G860), .ZN(G145));
  XNOR2_X1  g447(.A(new_n814), .B(new_n786), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n799), .Z(new_n874));
  AND3_X1   g449(.A1(new_n509), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT71), .B1(new_n509), .B2(KEYINPUT4), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n510), .B(new_n507), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n494), .A2(new_n495), .B1(new_n500), .B2(new_n503), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n873), .B(new_n799), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G164), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n481), .A2(G130), .B1(G142), .B2(new_n485), .ZN(new_n884));
  NOR2_X1   g459(.A1(G106), .A2(G2105), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n650), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n715), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n891));
  INV_X1    g466(.A(new_n889), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(new_n882), .A3(new_n880), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n883), .A2(KEYINPUT110), .A3(new_n889), .ZN(new_n895));
  XOR2_X1   g470(.A(new_n646), .B(KEYINPUT109), .Z(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n846), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G162), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n896), .B(G160), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n490), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n890), .A2(new_n898), .A3(new_n900), .A4(new_n893), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g481(.A(new_n636), .B(new_n867), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n635), .A2(new_n825), .A3(new_n623), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n625), .A2(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n915), .A3(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(KEYINPUT111), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n908), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n625), .B(new_n825), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n907), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(new_n913), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n907), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  INV_X1    g499(.A(new_n920), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G288), .B(new_n610), .ZN(new_n927));
  XNOR2_X1  g502(.A(G305), .B(G166), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n927), .B(new_n928), .Z(new_n929));
  AND3_X1   g504(.A1(new_n921), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n921), .B2(new_n926), .ZN(new_n931));
  OAI21_X1  g506(.A(G868), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n861), .A2(G868), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(G295));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n932), .A2(new_n936), .A3(new_n934), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n932), .B2(new_n934), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(G331));
  XNOR2_X1  g514(.A(G171), .B(G286), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n867), .B(new_n940), .Z(new_n941));
  XNOR2_X1  g516(.A(new_n914), .B(KEYINPUT115), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n916), .B(KEYINPUT114), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n867), .A2(new_n940), .A3(KEYINPUT113), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n945), .B1(new_n941), .B2(KEYINPUT113), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n911), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n929), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n917), .A2(new_n913), .A3(new_n946), .ZN(new_n949));
  INV_X1    g524(.A(new_n929), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n941), .A2(new_n919), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n903), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n948), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n956), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n948), .A2(new_n954), .A3(KEYINPUT43), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT44), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(G164), .B2(G1384), .ZN(new_n967));
  NAND2_X1  g542(.A1(G160), .A2(G40), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G2067), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n799), .B(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n814), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n715), .B(new_n721), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n969), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n969), .ZN(new_n977));
  NOR2_X1   g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT116), .ZN(new_n979));
  NAND2_X1  g554(.A1(G290), .A2(G1986), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n979), .B(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n843), .A2(G40), .A3(new_n845), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n877), .B2(new_n878), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n983), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n985));
  AOI211_X1 g560(.A(new_n966), .B(G1384), .C1(new_n877), .C2(new_n878), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G2078), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n983), .B1(new_n984), .B2(new_n991), .ZN(new_n992));
  AOI211_X1 g567(.A(KEYINPUT50), .B(G1384), .C1(new_n877), .C2(new_n878), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n989), .A2(new_n990), .B1(new_n994), .B2(new_n818), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n987), .A2(KEYINPUT53), .A3(new_n988), .ZN(new_n996));
  AOI211_X1 g571(.A(KEYINPUT62), .B(G301), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT117), .B(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(G286), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT123), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n754), .B1(new_n985), .B2(new_n986), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT121), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OR3_X1    g578(.A1(new_n992), .A2(G2084), .A3(new_n993), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT121), .B(new_n754), .C1(new_n985), .C2(new_n986), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1003), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI211_X1 g581(.A(KEYINPUT51), .B(new_n1000), .C1(new_n1006), .C2(new_n998), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT124), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1000), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT124), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(new_n1011), .A3(G8), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n1006), .B2(new_n1000), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n997), .B(new_n1007), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT58), .B(G1341), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n984), .A2(new_n983), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT122), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n984), .A2(KEYINPUT122), .A3(new_n983), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n985), .A2(G1996), .A3(new_n986), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n558), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT59), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n558), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n827), .B1(new_n992), .B2(new_n993), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n613), .A2(new_n577), .B1(new_n582), .B2(new_n518), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n1030), .A2(G651), .B1(G91), .B2(new_n587), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT57), .B1(new_n572), .B2(new_n574), .ZN(new_n1032));
  AOI22_X1  g607(.A1(G299), .A2(KEYINPUT57), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT56), .B(G2072), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n967), .A2(new_n1034), .A3(new_n983), .A4(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1029), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT61), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT61), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1029), .A2(new_n1033), .A3(new_n1036), .A4(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1020), .A2(new_n970), .A3(new_n1021), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n805), .B1(new_n992), .B2(new_n993), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT60), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1042), .A2(new_n626), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1042), .A2(new_n625), .A3(new_n1043), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n625), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT60), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1028), .A2(new_n1041), .A3(new_n1045), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1037), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n1029), .A2(new_n1036), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1051), .A2(new_n1033), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n471), .A2(new_n475), .A3(G40), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT125), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n967), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n990), .B1(new_n1058), .B2(KEYINPUT126), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n988), .C1(KEYINPUT126), .C2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n995), .B1(new_n1060), .B2(new_n986), .ZN(new_n1061));
  XNOR2_X1  g636(.A(G171), .B(KEYINPUT54), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n995), .A2(new_n996), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(new_n1064), .B2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1053), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1016), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n730), .A2(G1976), .ZN(new_n1068));
  INV_X1    g643(.A(new_n998), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n984), .B2(new_n983), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n730), .A2(G1976), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1073), .A2(KEYINPUT118), .A3(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n994), .A2(G2090), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n987), .A2(G1971), .ZN(new_n1081));
  OAI21_X1  g656(.A(G8), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G303), .A2(G8), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT55), .ZN(new_n1084));
  OR2_X1    g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n998), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1084), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G305), .A2(G1981), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1981), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n735), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(KEYINPUT49), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT49), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1095), .A3(new_n1070), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1096), .A2(KEYINPUT119), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(KEYINPUT119), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1079), .A2(new_n1085), .A3(new_n1087), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1007), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1006), .A2(new_n1011), .A3(G8), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1011), .B1(new_n1006), .B2(G8), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1102), .A2(new_n1103), .A3(new_n1000), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1015), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1064), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1100), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1067), .A2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G288), .A2(G1976), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1112));
  OR3_X1    g687(.A1(new_n1112), .A2(KEYINPUT120), .A3(new_n1088), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT120), .B1(new_n1112), .B2(new_n1088), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1070), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1087), .A2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1006), .A2(G168), .A3(new_n998), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1085), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(new_n1099), .A3(new_n1079), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1079), .A2(new_n1099), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT63), .B1(new_n1122), .B2(new_n1118), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1115), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n982), .B1(new_n1109), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n814), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n977), .B1(new_n971), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n969), .A2(new_n972), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT46), .Z(new_n1129));
  NOR2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  XOR2_X1   g705(.A(new_n1130), .B(KEYINPUT47), .Z(new_n1131));
  NOR3_X1   g706(.A1(new_n974), .A2(new_n721), .A3(new_n715), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n799), .A2(G2067), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n969), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n969), .A2(new_n978), .ZN(new_n1135));
  XNOR2_X1  g710(.A(new_n1135), .B(KEYINPUT48), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n976), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1131), .A2(new_n1134), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT127), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1138), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1115), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n1067), .B2(new_n1108), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1140), .B(new_n1141), .C1(new_n1143), .C2(new_n982), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1139), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g720(.A1(new_n905), .A2(G319), .ZN(new_n1147));
  NOR2_X1   g721(.A1(G401), .A2(G229), .ZN(new_n1148));
  NAND4_X1  g722(.A1(new_n1147), .A2(new_n959), .A3(new_n686), .A4(new_n1148), .ZN(G225));
  INV_X1    g723(.A(G225), .ZN(G308));
endmodule


