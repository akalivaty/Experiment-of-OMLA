//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989;
  OAI21_X1  g000(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT93), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(new_n204), .B2(new_n207), .ZN(new_n209));
  XOR2_X1   g008(.A(KEYINPUT95), .B(G36gat), .Z(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT94), .B(G29gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G43gat), .A2(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(G43gat), .A2(G50gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT15), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n220));
  XOR2_X1   g019(.A(KEYINPUT96), .B(G50gat), .Z(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(G43gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n202), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n222), .A2(new_n217), .A3(new_n212), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT97), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT17), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n219), .A2(new_n224), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT97), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n229), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n233), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n235), .B1(G1gat), .B2(new_n233), .ZN(new_n236));
  INV_X1    g035(.A(G8gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n225), .A2(new_n238), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(G229gat), .A2(G233gat), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n240), .A2(KEYINPUT18), .A3(new_n242), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n225), .B(new_n238), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT99), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n244), .A2(KEYINPUT99), .A3(new_n248), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n241), .B1(new_n231), .B2(new_n239), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT18), .B1(new_n253), .B2(new_n243), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT11), .B(G169gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT12), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n253), .A2(new_n243), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT18), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT100), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT100), .ZN(new_n265));
  AOI211_X1 g064(.A(new_n265), .B(KEYINPUT18), .C1(new_n253), .C2(new_n243), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n249), .A2(new_n261), .ZN(new_n268));
  AOI22_X1  g067(.A1(new_n256), .A2(new_n261), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G183gat), .B(G211gat), .Z(new_n270));
  OR2_X1    g069(.A1(G57gat), .A2(G64gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G57gat), .A2(G64gat), .ZN(new_n272));
  AND2_X1   g071(.A1(G71gat), .A2(G78gat), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n271), .B(new_n272), .C1(new_n273), .C2(KEYINPUT9), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(KEYINPUT101), .B2(new_n273), .ZN(new_n275));
  NOR2_X1   g074(.A1(G71gat), .A2(G78gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n277), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n279), .B(new_n274), .C1(KEYINPUT101), .C2(new_n273), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n278), .A2(KEYINPUT102), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT102), .B1(new_n278), .B2(new_n280), .ZN(new_n282));
  OR2_X1    g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT21), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n285), .B(KEYINPUT103), .Z(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n287));
  NAND2_X1  g086(.A1(G231gat), .A2(G233gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n285), .B(KEYINPUT103), .ZN(new_n291));
  INV_X1    g090(.A(new_n289), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G127gat), .B(G155gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n290), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n295), .B1(new_n290), .B2(new_n293), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n270), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(new_n270), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(new_n296), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n238), .B1(new_n283), .B2(new_n284), .ZN(new_n304));
  XOR2_X1   g103(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n302), .A3(new_n306), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G85gat), .ZN(new_n311));
  INV_X1    g110(.A(G92gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT107), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT107), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(G85gat), .A3(G92gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n315), .A3(KEYINPUT7), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n317));
  OAI211_X1 g116(.A(KEYINPUT107), .B(new_n317), .C1(new_n311), .C2(new_n312), .ZN(new_n318));
  NAND2_X1  g117(.A1(G99gat), .A2(G106gat), .ZN(new_n319));
  AOI22_X1  g118(.A1(KEYINPUT8), .A2(new_n319), .B1(new_n311), .B2(new_n312), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(G99gat), .B(G106gat), .Z(new_n322));
  OR3_X1    g121(.A1(new_n321), .A2(KEYINPUT108), .A3(new_n322), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n321), .A2(new_n322), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n322), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT108), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n231), .A2(new_n232), .A3(new_n323), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n323), .ZN(new_n328));
  AND2_X1   g127(.A1(G232gat), .A2(G233gat), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n328), .A2(new_n228), .B1(KEYINPUT41), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G190gat), .B(G218gat), .Z(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n329), .A2(KEYINPUT41), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT106), .ZN(new_n336));
  XNOR2_X1  g135(.A(G134gat), .B(G162gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n331), .A2(new_n332), .ZN(new_n340));
  OR3_X1    g139(.A1(new_n334), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n334), .B2(new_n340), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G230gat), .ZN(new_n345));
  INV_X1    g144(.A(G233gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n278), .A2(new_n280), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n324), .A3(new_n325), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT109), .B(KEYINPUT10), .Z(new_n350));
  NOR2_X1   g149(.A1(new_n281), .A2(new_n282), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n349), .B(new_n350), .C1(new_n328), .C2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n328), .A2(new_n351), .A3(KEYINPUT10), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n347), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n328), .B2(new_n351), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n347), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G120gat), .B(G148gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT110), .ZN(new_n360));
  XNOR2_X1  g159(.A(G176gat), .B(G204gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n357), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n310), .A2(new_n344), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369));
  INV_X1    g168(.A(G155gat), .ZN(new_n370));
  INV_X1    g169(.A(G162gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G141gat), .B(G148gat), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n369), .B(new_n372), .C1(new_n373), .C2(KEYINPUT2), .ZN(new_n374));
  INV_X1    g173(.A(G141gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G148gat), .ZN(new_n376));
  INV_X1    g175(.A(G148gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G141gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n378), .A3(KEYINPUT81), .ZN(new_n379));
  OR3_X1    g178(.A1(new_n377), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n372), .A2(new_n369), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n369), .A2(KEYINPUT82), .A3(KEYINPUT2), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT82), .B1(new_n369), .B2(KEYINPUT2), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n374), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n369), .A2(KEYINPUT2), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n369), .A2(KEYINPUT82), .A3(KEYINPUT2), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(new_n381), .A3(new_n379), .A4(new_n380), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT85), .A3(new_n374), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n388), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  XOR2_X1   g196(.A(G127gat), .B(G134gat), .Z(new_n398));
  INV_X1    g197(.A(G113gat), .ZN(new_n399));
  INV_X1    g198(.A(G120gat), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT1), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT70), .B(G113gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G120gat), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n401), .B1(new_n399), .B2(new_n400), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n403), .A2(new_n405), .B1(new_n406), .B2(new_n398), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n396), .A2(new_n397), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n374), .A3(new_n394), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n409), .B1(new_n410), .B2(KEYINPUT4), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n386), .A2(KEYINPUT83), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n394), .A2(new_n414), .A3(new_n374), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT3), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT84), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n413), .A2(new_n415), .A3(new_n418), .A4(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n405), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n406), .A2(new_n398), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT3), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n374), .B(new_n423), .C1(new_n382), .C2(new_n385), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n417), .A2(new_n419), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n396), .A2(new_n409), .A3(new_n397), .A4(new_n407), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n412), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  OR3_X1    g228(.A1(new_n427), .A2(KEYINPUT5), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n410), .B2(new_n397), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n388), .A2(new_n395), .A3(KEYINPUT4), .A4(new_n407), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n415), .A3(new_n422), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n410), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n429), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT5), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n428), .B1(new_n435), .B2(new_n410), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT86), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AOI221_X4 g241(.A(new_n431), .B1(new_n425), .B2(new_n434), .C1(new_n439), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n439), .A2(new_n442), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n434), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT87), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n430), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G1gat), .B(G29gat), .Z(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT88), .B(KEYINPUT0), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  INV_X1    g253(.A(new_n452), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n430), .B(new_n455), .C1(new_n443), .C2(new_n446), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(KEYINPUT6), .A3(new_n452), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT77), .ZN(new_n460));
  NAND2_X1  g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n464), .A2(KEYINPUT26), .ZN(new_n465));
  INV_X1    g264(.A(G169gat), .ZN(new_n466));
  INV_X1    g265(.A(G176gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G183gat), .ZN(new_n470));
  INV_X1    g269(.A(G190gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(KEYINPUT26), .B2(new_n464), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(KEYINPUT27), .B(G183gat), .Z(new_n476));
  INV_X1    g275(.A(KEYINPUT28), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n476), .A2(new_n477), .A3(G190gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT68), .B(G183gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT27), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT28), .B1(new_n484), .B2(new_n471), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n479), .B1(new_n485), .B2(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n470), .A2(KEYINPUT68), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G183gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n480), .B1(new_n490), .B2(KEYINPUT27), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n477), .B1(new_n491), .B2(G190gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT69), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n475), .B1(new_n486), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n496));
  OR3_X1    g295(.A1(new_n496), .A2(KEYINPUT67), .A3(new_n472), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT67), .B1(new_n496), .B2(new_n472), .ZN(new_n498));
  NAND3_X1  g297(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n471), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n464), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n502), .B1(new_n468), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n464), .A2(KEYINPUT23), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n504), .A2(KEYINPUT25), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n470), .A2(new_n471), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n499), .B(new_n508), .C1(new_n472), .C2(KEYINPUT24), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT65), .B(G176gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n466), .A2(KEYINPUT23), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n509), .B(new_n504), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n463), .B1(new_n495), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n478), .B1(new_n492), .B2(new_n493), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n485), .A2(KEYINPUT69), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n474), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n501), .A2(new_n506), .B1(new_n512), .B2(new_n513), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT75), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n495), .A2(new_n522), .A3(new_n515), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n461), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n516), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G211gat), .B(G218gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT74), .ZN(new_n528));
  INV_X1    g327(.A(G211gat), .ZN(new_n529));
  OR2_X1    g328(.A1(KEYINPUT73), .A2(G218gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(KEYINPUT73), .A2(G218gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n533));
  XNOR2_X1  g332(.A(G197gat), .B(G204gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n528), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  OAI221_X1 g335(.A(new_n534), .B1(new_n527), .B2(KEYINPUT74), .C1(new_n532), .C2(KEYINPUT22), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n460), .B1(new_n526), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n495), .A2(new_n525), .A3(new_n515), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT76), .B(KEYINPUT29), .Z(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n461), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n541), .B(new_n539), .C1(new_n524), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n461), .B1(new_n521), .B2(new_n523), .ZN(new_n545));
  OAI211_X1 g344(.A(KEYINPUT77), .B(new_n538), .C1(new_n545), .C2(new_n516), .ZN(new_n546));
  XNOR2_X1  g345(.A(G8gat), .B(G36gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(G64gat), .B(G92gat), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(new_n548), .Z(new_n549));
  NAND4_X1  g348(.A1(new_n540), .A2(new_n544), .A3(new_n546), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT80), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n546), .A2(new_n544), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT80), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(new_n553), .A3(new_n540), .A4(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n524), .A2(new_n525), .ZN(new_n558));
  INV_X1    g357(.A(new_n516), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT77), .B1(new_n560), .B2(new_n538), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n544), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT78), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n549), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT78), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n540), .A2(new_n565), .A3(new_n544), .A4(new_n546), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n564), .A2(new_n556), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n540), .A2(new_n544), .A3(new_n546), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT79), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT79), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n552), .A2(new_n571), .A3(new_n540), .A4(new_n568), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n459), .A2(new_n557), .A3(new_n567), .A4(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(G78gat), .B(G106gat), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT90), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT92), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n424), .A2(new_n542), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n580), .B2(new_n538), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n539), .A2(new_n579), .A3(KEYINPUT92), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n413), .A2(new_n415), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT29), .B1(new_n536), .B2(new_n537), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n584), .B(new_n585), .C1(KEYINPUT3), .C2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n413), .A3(new_n415), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(KEYINPUT91), .A3(new_n416), .ZN(new_n589));
  INV_X1    g388(.A(G228gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(new_n346), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n583), .A2(new_n587), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  OR3_X1    g391(.A1(new_n533), .A2(new_n527), .A3(new_n535), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n527), .B1(new_n533), .B2(new_n535), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n542), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n595), .A2(new_n423), .B1(new_n388), .B2(new_n395), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n538), .ZN(new_n597));
  OAI22_X1  g396(.A1(new_n596), .A2(new_n597), .B1(new_n590), .B2(new_n346), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G22gat), .ZN(new_n600));
  INV_X1    g399(.A(G22gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n592), .A2(new_n601), .A3(new_n598), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n577), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT31), .B(G50gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(new_n577), .A3(new_n602), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n605), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n600), .A2(new_n577), .A3(new_n602), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT72), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n407), .B1(new_n519), .B2(new_n520), .ZN(new_n613));
  INV_X1    g412(.A(G227gat), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n346), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n495), .A2(new_n422), .A3(new_n515), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT32), .ZN(new_n618));
  XOR2_X1   g417(.A(G15gat), .B(G43gat), .Z(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G99gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n622), .B1(new_n617), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT34), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n613), .A2(new_n616), .ZN(new_n626));
  INV_X1    g425(.A(new_n615), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI211_X1 g427(.A(KEYINPUT34), .B(new_n615), .C1(new_n613), .C2(new_n616), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n624), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n624), .A2(new_n628), .A3(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n618), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n628), .ZN(new_n634));
  INV_X1    g433(.A(new_n629), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n617), .A2(new_n623), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n622), .ZN(new_n637));
  INV_X1    g436(.A(new_n618), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n637), .A2(new_n638), .A3(new_n630), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n612), .B1(new_n633), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT71), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n633), .B2(new_n639), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n643));
  OAI22_X1  g442(.A1(KEYINPUT71), .A2(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n631), .A2(new_n632), .A3(new_n618), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n638), .B1(new_n637), .B2(new_n630), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT72), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n641), .A3(KEYINPUT36), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n574), .A2(new_n611), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n427), .A2(new_n429), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n435), .A2(new_n428), .A3(new_n410), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT39), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n427), .A2(new_n653), .A3(new_n429), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n652), .A2(new_n455), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n652), .A2(KEYINPUT40), .A3(new_n455), .A4(new_n654), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n453), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n573), .A2(new_n567), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT30), .B1(new_n551), .B2(new_n554), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n611), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n552), .A2(new_n540), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT37), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n549), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n563), .A2(KEYINPUT37), .A3(new_n566), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n541), .B(new_n538), .C1(new_n524), .C2(new_n543), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n670), .A2(KEYINPUT37), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n560), .A2(new_n539), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT38), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n673), .B(new_n564), .C1(new_n665), .C2(KEYINPUT37), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n457), .A2(new_n674), .A3(new_n555), .A4(new_n458), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n662), .B(new_n663), .C1(new_n669), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n649), .A2(new_n676), .ZN(new_n677));
  AND4_X1   g476(.A1(new_n607), .A2(new_n610), .A3(new_n639), .A4(new_n633), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT35), .B1(new_n574), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n660), .A2(new_n661), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT35), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n459), .A4(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  AOI211_X1 g483(.A(new_n269), .B(new_n368), .C1(new_n677), .C2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n459), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  INV_X1    g487(.A(new_n681), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AND3_X1   g489(.A1(new_n685), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n237), .B1(new_n685), .B2(new_n689), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT42), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT42), .B2(new_n691), .ZN(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n633), .A2(new_n639), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n685), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n644), .A2(new_n648), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n685), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n698), .B1(new_n701), .B2(new_n695), .ZN(G1326gat));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n611), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT43), .B(G22gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1327gat));
  AOI21_X1  g504(.A(new_n344), .B1(new_n677), .B2(new_n684), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n310), .A2(new_n269), .A3(new_n366), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(new_n459), .A3(new_n211), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT45), .Z(new_n710));
  INV_X1    g509(.A(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n677), .A2(new_n684), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n677), .A2(new_n684), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n344), .A2(KEYINPUT44), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n712), .A2(new_n343), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT44), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n711), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n686), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n211), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n721), .B1(new_n720), .B2(new_n686), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n710), .B1(new_n723), .B2(new_n724), .ZN(G1328gat));
  NOR3_X1   g524(.A1(new_n708), .A2(new_n681), .A3(new_n210), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT46), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n720), .A2(KEYINPUT113), .A3(new_n689), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n210), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT113), .B1(new_n720), .B2(new_n689), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(G1329gat));
  NOR2_X1   g530(.A1(new_n696), .A2(G43gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n706), .A2(new_n707), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n717), .A2(new_n719), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n700), .A3(new_n707), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  INV_X1    g537(.A(G43gat), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n720), .B2(new_n700), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n733), .A2(KEYINPUT47), .ZN(new_n741));
  OAI22_X1  g540(.A1(new_n738), .A2(KEYINPUT47), .B1(new_n740), .B2(new_n741), .ZN(G1330gat));
  AND2_X1   g541(.A1(new_n611), .A2(new_n221), .ZN(new_n743));
  AND3_X1   g542(.A1(new_n736), .A2(new_n707), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n708), .A2(new_n663), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(new_n221), .ZN(new_n746));
  OAI21_X1  g545(.A(KEYINPUT48), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n720), .A2(new_n743), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n748), .B(new_n749), .C1(new_n221), .C2(new_n745), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(G1331gat));
  AND2_X1   g550(.A1(new_n713), .A2(new_n715), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n308), .A2(new_n309), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n267), .A2(new_n268), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n244), .A2(KEYINPUT99), .A3(new_n248), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT99), .B1(new_n244), .B2(new_n248), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n755), .A2(new_n756), .A3(new_n254), .ZN(new_n757));
  INV_X1    g556(.A(new_n261), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n754), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n753), .A2(new_n759), .A3(new_n343), .A4(new_n367), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n686), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n689), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT49), .B(G64gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n689), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1333gat));
  NOR2_X1   g567(.A1(new_n696), .A2(G71gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n760), .A3(new_n769), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n713), .A2(new_n700), .A3(new_n715), .A4(new_n760), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G71gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n761), .A2(new_n611), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g576(.A1(new_n310), .A2(new_n759), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n366), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n717), .B2(new_n719), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n780), .A2(new_n686), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n706), .A2(KEYINPUT51), .A3(new_n778), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT51), .B1(new_n706), .B2(new_n778), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n686), .A2(new_n311), .A3(new_n366), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n781), .A2(new_n311), .B1(new_n785), .B2(new_n786), .ZN(G1336gat));
  AOI21_X1  g586(.A(new_n312), .B1(new_n780), .B2(new_n689), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n367), .A2(G92gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n689), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT52), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n689), .B(new_n789), .C1(new_n783), .C2(new_n784), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  AOI211_X1 g593(.A(new_n681), .B(new_n779), .C1(new_n717), .C2(new_n719), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n312), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1337gat));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798));
  INV_X1    g597(.A(G99gat), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n780), .B2(new_n700), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n367), .A2(G99gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n697), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n785), .A2(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n800), .B2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n697), .B(new_n801), .C1(new_n783), .C2(new_n784), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n699), .B(new_n779), .C1(new_n717), .C2(new_n719), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n805), .B(KEYINPUT115), .C1(new_n806), .C2(new_n799), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1338gat));
  NOR3_X1   g607(.A1(new_n663), .A2(G106gat), .A3(new_n367), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT116), .ZN(new_n810));
  INV_X1    g609(.A(new_n784), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(new_n782), .ZN(new_n812));
  INV_X1    g611(.A(new_n779), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n736), .A2(new_n611), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  INV_X1    g615(.A(new_n809), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n785), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(G106gat), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n780), .B2(new_n611), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n815), .A2(new_n816), .B1(new_n818), .B2(new_n820), .ZN(G1339gat));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n352), .A2(new_n353), .ZN(new_n823));
  INV_X1    g622(.A(new_n347), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n825), .A2(new_n826), .A3(new_n354), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n364), .B1(new_n354), .B2(new_n826), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n822), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n355), .A2(KEYINPUT54), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT55), .B(new_n828), .C1(new_n831), .C2(new_n825), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n832), .A3(new_n365), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n830), .A2(new_n832), .A3(KEYINPUT117), .A4(new_n365), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n759), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n253), .A2(new_n243), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n245), .A2(new_n247), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n260), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n754), .A2(new_n366), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n343), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n343), .A2(new_n754), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n835), .A2(new_n836), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n753), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n310), .A2(new_n269), .A3(new_n344), .A4(new_n367), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n679), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n689), .A2(new_n459), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n848), .A2(new_n759), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(G113gat), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n852), .B1(new_n404), .B2(new_n851), .ZN(G1340gat));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n366), .A3(new_n849), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(G120gat), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n848), .A2(new_n310), .A3(new_n849), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g656(.A1(new_n689), .A2(new_n344), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(KEYINPUT118), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n859), .A2(G134gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n848), .A2(new_n686), .ZN(new_n861));
  XOR2_X1   g660(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n860), .B2(new_n861), .ZN(new_n865));
  INV_X1    g664(.A(new_n858), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(G1343gat));
  OAI21_X1  g667(.A(new_n841), .B1(new_n269), .B2(new_n833), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT120), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n841), .B(KEYINPUT120), .C1(new_n269), .C2(new_n833), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n344), .ZN(new_n874));
  INV_X1    g673(.A(new_n845), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n310), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n847), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n611), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n663), .B1(new_n846), .B2(new_n847), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n700), .A2(new_n459), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n681), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n269), .A2(new_n375), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n879), .A2(new_n882), .A3(new_n885), .A4(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT121), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n880), .A3(new_n759), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n890), .A2(new_n375), .B1(KEYINPUT121), .B2(new_n888), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n887), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n889), .B1(new_n887), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(G1344gat));
  AND2_X1   g693(.A1(new_n885), .A2(new_n880), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n377), .A3(new_n366), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n879), .A2(new_n882), .A3(new_n366), .A4(new_n885), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n377), .A2(KEYINPUT59), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n880), .A2(new_n881), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n663), .A2(KEYINPUT57), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n343), .B1(new_n871), .B2(new_n872), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n843), .A2(new_n833), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n753), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n847), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n366), .A3(new_n885), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n900), .B1(new_n909), .B2(G148gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n896), .B1(new_n899), .B2(new_n910), .ZN(G1345gat));
  NAND3_X1  g710(.A1(new_n879), .A2(new_n885), .A3(new_n882), .ZN(new_n912));
  OAI21_X1  g711(.A(G155gat), .B1(new_n912), .B2(new_n753), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n370), .A3(new_n310), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n912), .B2(new_n344), .ZN(new_n916));
  INV_X1    g715(.A(new_n859), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n917), .A2(new_n371), .A3(new_n883), .A4(new_n880), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1347gat));
  AOI21_X1  g718(.A(new_n686), .B1(new_n846), .B2(new_n847), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(KEYINPUT122), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922));
  AOI211_X1 g721(.A(new_n922), .B(new_n686), .C1(new_n846), .C2(new_n847), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n679), .A2(new_n681), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n759), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n920), .A2(new_n925), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n269), .A2(new_n466), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n926), .A2(new_n466), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  OAI211_X1 g728(.A(new_n366), .B(new_n925), .C1(new_n921), .C2(new_n923), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n467), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n510), .A3(new_n366), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(KEYINPUT123), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1349gat));
  NAND2_X1  g736(.A1(new_n846), .A2(new_n847), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n938), .A2(new_n459), .A3(new_n310), .A4(new_n925), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n920), .A2(KEYINPUT124), .A3(new_n310), .A4(new_n925), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n490), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n753), .A2(new_n476), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n925), .B(new_n945), .C1(new_n921), .C2(new_n923), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g746(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(G1350gat));
  AOI21_X1  g748(.A(new_n471), .B1(new_n927), .B2(new_n343), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT61), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n344), .A2(G190gat), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n925), .B(new_n953), .C1(new_n921), .C2(new_n923), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n952), .A2(new_n956), .ZN(G1351gat));
  INV_X1    g756(.A(G197gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n699), .A2(new_n459), .A3(new_n689), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n901), .A2(new_n907), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n960), .B2(new_n759), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n700), .A2(new_n681), .A3(new_n663), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n269), .A2(G197gat), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n962), .B(new_n963), .C1(new_n921), .C2(new_n923), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT127), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  NOR4_X1   g766(.A1(new_n901), .A2(new_n907), .A3(new_n269), .A4(new_n959), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n967), .B(new_n964), .C1(new_n968), .C2(new_n958), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n966), .A2(new_n969), .ZN(G1352gat));
  NOR2_X1   g769(.A1(new_n367), .A2(G204gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n924), .A2(new_n962), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT62), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n960), .A2(new_n366), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G204gat), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n924), .A2(new_n976), .A3(new_n962), .A4(new_n971), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n973), .A2(new_n975), .A3(new_n977), .ZN(G1353gat));
  INV_X1    g777(.A(KEYINPUT63), .ZN(new_n979));
  AOI211_X1 g778(.A(new_n979), .B(new_n529), .C1(new_n960), .C2(new_n310), .ZN(new_n980));
  INV_X1    g779(.A(new_n959), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n908), .A2(new_n310), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(KEYINPUT63), .B1(new_n982), .B2(G211gat), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n924), .A2(new_n962), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n310), .A2(new_n529), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n980), .A2(new_n983), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  NAND3_X1  g785(.A1(new_n924), .A2(new_n343), .A3(new_n962), .ZN(new_n987));
  INV_X1    g786(.A(G218gat), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n344), .B1(new_n530), .B2(new_n531), .ZN(new_n989));
  AOI22_X1  g788(.A1(new_n987), .A2(new_n988), .B1(new_n960), .B2(new_n989), .ZN(G1355gat));
endmodule


