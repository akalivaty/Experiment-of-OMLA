//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT6), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT78), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT78), .A2(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G104), .A3(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n191), .A2(G104), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT3), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G104), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT3), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n197), .A2(G101), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G101), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT78), .A2(G107), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT78), .A2(G107), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n206), .B2(new_n198), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT79), .B1(new_n201), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT2), .A2(G113), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n209), .B(KEYINPUT67), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT2), .A2(G113), .ZN(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(KEYINPUT5), .ZN(new_n215));
  INV_X1    g029(.A(G113), .ZN(new_n216));
  INV_X1    g030(.A(G116), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G119), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT5), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n214), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n204), .A2(new_n205), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n195), .B1(new_n222), .B2(G104), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n202), .B(new_n199), .C1(new_n223), .C2(KEYINPUT3), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n225));
  INV_X1    g039(.A(new_n207), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n208), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G110), .B(G122), .ZN(new_n229));
  OAI21_X1  g043(.A(G101), .B1(new_n197), .B2(new_n200), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n224), .A3(KEYINPUT4), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n212), .B1(new_n210), .B2(new_n211), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n214), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n234), .B(G101), .C1(new_n197), .C2(new_n200), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n228), .A2(new_n229), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n229), .B1(new_n228), .B2(new_n236), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n189), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n236), .ZN(new_n240));
  INV_X1    g054(.A(new_n229), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n188), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT65), .B1(new_n246), .B2(G143), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(G143), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G143), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n245), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(G146), .ZN(new_n254));
  AND4_X1   g068(.A1(KEYINPUT0), .A2(new_n248), .A3(new_n254), .A4(G128), .ZN(new_n255));
  OAI21_X1  g069(.A(G125), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G125), .ZN(new_n257));
  INV_X1    g071(.A(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(KEYINPUT1), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n248), .A3(new_n254), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n246), .A2(KEYINPUT65), .A3(G143), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n248), .B2(new_n247), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n258), .B1(new_n248), .B2(KEYINPUT1), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n257), .B(new_n260), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n256), .A2(new_n264), .A3(KEYINPUT83), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT83), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(G125), .C1(new_n253), .C2(new_n255), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G224), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(G902), .B1(new_n244), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G210), .B1(G237), .B2(G902), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT86), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n268), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n224), .A2(new_n226), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n221), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n220), .A2(KEYINPUT84), .ZN(new_n280));
  INV_X1    g094(.A(G119), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G116), .ZN(new_n282));
  OAI21_X1  g096(.A(G113), .B1(new_n282), .B2(KEYINPUT5), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT84), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n215), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n213), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n226), .A3(new_n224), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n229), .B(KEYINPUT8), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n276), .B1(new_n256), .B2(new_n264), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT85), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n291), .A2(KEYINPUT85), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n277), .B(new_n290), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n274), .B1(new_n268), .B2(new_n276), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT87), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n294), .ZN(new_n298));
  INV_X1    g112(.A(new_n289), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n201), .A2(new_n207), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n287), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n298), .A2(new_n292), .B1(new_n301), .B2(new_n279), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n303));
  INV_X1    g117(.A(new_n296), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n277), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n228), .A2(new_n236), .A3(new_n229), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n272), .A2(new_n273), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT88), .ZN(new_n309));
  INV_X1    g123(.A(G902), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n188), .B1(new_n242), .B2(new_n306), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n238), .A2(new_n189), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n271), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AND4_X1   g127(.A1(new_n310), .A2(new_n307), .A3(new_n313), .A4(new_n273), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n273), .B1(new_n272), .B2(new_n307), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n309), .B1(new_n316), .B2(KEYINPUT88), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n257), .A2(G140), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(KEYINPUT72), .A3(G125), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(KEYINPUT16), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT16), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G146), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n324), .A2(new_n246), .A3(new_n326), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n281), .B2(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n258), .A2(KEYINPUT23), .A3(G119), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n281), .A2(G128), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT70), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT70), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n333), .A2(new_n334), .A3(new_n338), .A4(new_n335), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(G110), .A3(new_n339), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n340), .A2(KEYINPUT71), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n327), .A2(KEYINPUT73), .A3(G146), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n258), .A2(G119), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n335), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n346), .B1(new_n340), .B2(KEYINPUT71), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n331), .A2(new_n341), .A3(new_n342), .A4(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n319), .A2(new_n320), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(G146), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n345), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(G110), .B2(new_n336), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n328), .A2(new_n349), .A3(new_n352), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n352), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n246), .B1(new_n324), .B2(new_n326), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT74), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G137), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n348), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n348), .B2(new_n359), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n310), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT25), .B(new_n310), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G217), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n371), .B1(G234), .B2(new_n310), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n364), .A2(new_n365), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n372), .A2(G902), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT76), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n249), .A2(new_n252), .ZN(new_n380));
  INV_X1    g194(.A(new_n245), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n255), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G137), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n383), .A2(G134), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(G134), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G134), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n388), .A2(G137), .ZN(new_n389));
  INV_X1    g203(.A(new_n386), .ZN(new_n390));
  NOR2_X1   g204(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G131), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n387), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n387), .B2(new_n392), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n382), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n387), .A2(new_n392), .A3(new_n393), .ZN(new_n397));
  OAI21_X1  g211(.A(G131), .B1(new_n389), .B2(new_n384), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n263), .B1(new_n252), .B2(new_n249), .ZN(new_n399));
  INV_X1    g213(.A(new_n260), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT30), .B1(new_n402), .B2(KEYINPUT64), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT64), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n405));
  AOI211_X1 g219(.A(new_n404), .B(new_n405), .C1(new_n396), .C2(new_n401), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n233), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT26), .B(G101), .Z(new_n408));
  NOR2_X1   g222(.A1(G237), .A2(G953), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G210), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n408), .B(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n214), .A2(new_n232), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n396), .A2(new_n415), .A3(new_n401), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT69), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT28), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n402), .A2(new_n233), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n421), .B2(new_n416), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n419), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(KEYINPUT69), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n413), .B(new_n420), .C1(new_n422), .C2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT31), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G472), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n407), .A2(KEYINPUT31), .A3(new_n414), .A4(new_n416), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n427), .A2(new_n428), .A3(new_n310), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT32), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n310), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n428), .A4(new_n427), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n418), .B1(new_n416), .B2(new_n419), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n396), .A2(new_n415), .A3(new_n401), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n415), .B1(new_n396), .B2(new_n401), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n437), .B1(new_n440), .B2(new_n419), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n413), .B1(new_n441), .B2(new_n420), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n442), .B2(KEYINPUT29), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n414), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n402), .A2(KEYINPUT64), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n405), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n402), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n415), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n413), .B1(new_n449), .B2(new_n438), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G472), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n379), .B1(new_n436), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(G214), .B1(G237), .B2(G902), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n456), .B(KEYINPUT81), .Z(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  OAI21_X1  g272(.A(G221), .B1(new_n458), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G469), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n208), .A2(KEYINPUT10), .A3(new_n462), .A4(new_n227), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n394), .A2(new_n395), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n231), .A2(new_n382), .A3(new_n235), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n248), .A2(new_n254), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n260), .B1(new_n466), .B2(new_n263), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n224), .A2(new_n226), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT10), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n269), .A2(G227), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT77), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G140), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n462), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n278), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n468), .ZN(new_n478));
  INV_X1    g292(.A(new_n464), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT12), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n481), .B(new_n464), .C1(new_n477), .C2(new_n468), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n471), .B(new_n475), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n463), .A2(new_n465), .A3(new_n470), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n479), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n475), .B1(new_n486), .B2(new_n471), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n461), .B(new_n310), .C1(new_n484), .C2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n461), .A2(new_n310), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n486), .A2(new_n471), .A3(new_n475), .ZN(new_n493));
  INV_X1    g307(.A(new_n468), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n462), .B1(new_n224), .B2(new_n226), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n479), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n481), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n478), .A2(KEYINPUT12), .A3(new_n479), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n475), .B1(new_n499), .B2(new_n471), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n492), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n471), .B1(new_n480), .B2(new_n482), .ZN(new_n502));
  INV_X1    g316(.A(new_n475), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n486), .A2(new_n471), .A3(new_n475), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(KEYINPUT80), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(G469), .A3(new_n506), .ZN(new_n507));
  AOI211_X1 g321(.A(new_n457), .B(new_n460), .C1(new_n491), .C2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(G237), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n269), .A3(G214), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n250), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n409), .A2(G143), .A3(G214), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(KEYINPUT18), .A2(G131), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n322), .A2(new_n516), .A3(new_n323), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n322), .B2(new_n323), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n517), .A2(new_n518), .A3(new_n246), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n515), .B1(new_n519), .B2(new_n351), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n518), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n322), .A2(new_n516), .A3(new_n323), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(G146), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n352), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT90), .A3(new_n515), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n331), .A2(new_n342), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n513), .A2(G131), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n511), .A2(new_n393), .A3(new_n512), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n533), .B2(new_n530), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n522), .A2(new_n527), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G113), .B(G122), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(new_n203), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n330), .A2(new_n329), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(new_n357), .ZN(new_n540));
  INV_X1    g354(.A(new_n342), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n520), .A2(new_n521), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT90), .B1(new_n526), .B2(new_n515), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n537), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT91), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n535), .A2(new_n547), .A3(new_n537), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n538), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G475), .B1(new_n549), .B2(G902), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT20), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n522), .A2(new_n527), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n533), .A2(new_n357), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n350), .A2(KEYINPUT19), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n517), .A2(new_n518), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(KEYINPUT19), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n553), .B1(new_n557), .B2(G146), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n537), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n545), .A2(KEYINPUT91), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n547), .B1(new_n535), .B2(new_n537), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(G475), .A2(G902), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n551), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n559), .B1(new_n546), .B2(new_n548), .ZN(new_n566));
  INV_X1    g380(.A(new_n564), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n566), .A2(KEYINPUT20), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n550), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G128), .B(G143), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT13), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n258), .A2(KEYINPUT13), .A3(G143), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n388), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n571), .A2(new_n573), .B1(new_n388), .B2(new_n570), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n217), .A2(G122), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT92), .ZN(new_n576));
  INV_X1    g390(.A(G122), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(G116), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n217), .A2(KEYINPUT92), .A3(G122), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n580), .A2(new_n222), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n222), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n458), .A2(new_n371), .A3(G953), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n570), .A2(new_n388), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n570), .A2(new_n388), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n580), .A2(new_n222), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT14), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n578), .B2(new_n579), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n575), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n578), .A2(new_n590), .A3(new_n579), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n191), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n583), .B(new_n584), .C1(new_n589), .C2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n593), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n597), .A2(new_n575), .A3(new_n591), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n588), .B(new_n587), .C1(new_n598), .C2(new_n191), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n584), .B1(new_n599), .B2(new_n583), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n310), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G478), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(KEYINPUT15), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n583), .B1(new_n589), .B2(new_n594), .ZN(new_n606));
  INV_X1    g420(.A(new_n584), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n608), .B2(new_n595), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT93), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n603), .A2(new_n605), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(KEYINPUT15), .B2(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT94), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT94), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n612), .A3(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(G234), .A2(G237), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(G952), .A3(new_n269), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(G902), .A3(G953), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT21), .B(G898), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n569), .A2(new_n617), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n317), .A2(new_n455), .A3(new_n508), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  AND3_X1   g441(.A1(new_n417), .A2(new_n425), .A3(new_n426), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n628), .B2(new_n432), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n629), .A2(KEYINPUT95), .A3(new_n430), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n631), .B(G472), .C1(new_n628), .C2(new_n432), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n460), .B1(new_n491), .B2(new_n507), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n307), .A2(new_n313), .A3(new_n310), .ZN(new_n635));
  INV_X1    g449(.A(new_n273), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n457), .B1(new_n637), .B2(new_n308), .ZN(new_n638));
  INV_X1    g452(.A(new_n379), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n633), .A2(new_n634), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT33), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n608), .B2(KEYINPUT96), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n608), .A2(new_n595), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(G478), .A3(new_n310), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT97), .B(G478), .Z(new_n646));
  NAND3_X1  g460(.A1(new_n603), .A2(new_n610), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n569), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n640), .A2(new_n624), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n203), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(new_n617), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n624), .B(KEYINPUT99), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n654), .A2(new_n569), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n640), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT35), .B(G107), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G9));
  INV_X1    g475(.A(new_n372), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n368), .B2(new_n369), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n348), .A2(new_n359), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n376), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n630), .B2(new_n632), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n317), .A2(new_n625), .A3(new_n508), .A4(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  OR2_X1    g487(.A1(new_n663), .A2(new_n668), .ZN(new_n674));
  INV_X1    g488(.A(new_n457), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n674), .B(new_n675), .C1(new_n314), .C2(new_n315), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n563), .A2(new_n551), .A3(new_n564), .ZN(new_n677));
  OAI21_X1  g491(.A(KEYINPUT20), .B1(new_n566), .B2(new_n567), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n619), .B(KEYINPUT100), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(G900), .B2(new_n621), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n617), .A2(new_n679), .A3(new_n550), .A4(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n501), .A2(G469), .A3(new_n506), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n488), .A2(new_n490), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n459), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n431), .A2(new_n435), .B1(G472), .B2(new_n453), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XNOR2_X1  g504(.A(new_n681), .B(KEYINPUT39), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n634), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT40), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n317), .B(KEYINPUT38), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n413), .B1(new_n407), .B2(new_n416), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n440), .A2(new_n413), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n310), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n436), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n569), .A2(new_n617), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n457), .A3(new_n674), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n694), .A3(new_n699), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  AND2_X1   g517(.A1(new_n645), .A2(new_n647), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n679), .B2(new_n550), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n638), .A2(new_n705), .A3(new_n674), .A4(new_n681), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n436), .A2(new_n454), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n634), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT101), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n676), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n569), .A2(new_n648), .A3(new_n681), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n688), .A2(new_n710), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  OAI21_X1  g529(.A(new_n675), .B1(new_n314), .B2(new_n315), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n310), .B1(new_n484), .B2(new_n487), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G469), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n459), .A3(new_n488), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n624), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n569), .A2(new_n721), .A3(new_n648), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n455), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND3_X1  g539(.A1(new_n720), .A2(new_n657), .A3(new_n455), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  AOI21_X1  g541(.A(new_n669), .B1(new_n436), .B2(new_n454), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n720), .A2(new_n625), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NOR2_X1   g544(.A1(new_n700), .A2(new_n716), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n719), .A2(new_n656), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n373), .A2(new_n733), .A3(new_n378), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT102), .B1(new_n663), .B2(new_n377), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT103), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n629), .A2(new_n430), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n737), .B1(new_n736), .B2(new_n738), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n731), .B(new_n732), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT104), .B(G122), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G24));
  NAND3_X1  g557(.A1(new_n569), .A2(new_n648), .A3(new_n681), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n674), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT105), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n629), .A2(new_n430), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n747), .B2(new_n669), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n744), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n720), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  INV_X1    g565(.A(KEYINPUT42), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n734), .A2(new_n735), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT109), .B1(new_n753), .B2(new_n687), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n707), .A2(new_n755), .A3(new_n736), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n637), .A2(KEYINPUT88), .A3(new_n308), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT88), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n314), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n457), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n504), .A2(new_n505), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n762), .B1(new_n764), .B2(G469), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n763), .A2(KEYINPUT106), .A3(new_n461), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n460), .B1(new_n767), .B2(new_n491), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n761), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n761), .B2(new_n768), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n757), .B(new_n712), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n761), .A2(new_n768), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(KEYINPUT107), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n761), .A2(new_n768), .A3(new_n769), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(KEYINPUT110), .A3(new_n712), .A4(new_n757), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n774), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n455), .B(new_n712), .C1(new_n770), .C2(new_n771), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n752), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT108), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT108), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n784), .A3(new_n752), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n780), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  INV_X1    g601(.A(new_n682), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n455), .B(new_n788), .C1(new_n770), .C2(new_n771), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT111), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n778), .A2(new_n791), .A3(new_n455), .A4(new_n788), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  NAND3_X1  g608(.A1(new_n679), .A2(new_n550), .A3(new_n648), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(KEYINPUT112), .B2(new_n798), .ZN(new_n799));
  AOI211_X1 g613(.A(new_n633), .B(new_n669), .C1(new_n797), .C2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(KEYINPUT44), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n761), .B1(new_n800), .B2(KEYINPUT44), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT45), .B1(new_n501), .B2(new_n506), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  OAI21_X1  g618(.A(G469), .B1(new_n763), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n490), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT46), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n488), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n806), .B2(new_n807), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n460), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n691), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n801), .A2(new_n802), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(new_n383), .ZN(G39));
  NAND4_X1  g628(.A1(new_n761), .A2(new_n712), .A3(new_n379), .A4(new_n687), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n811), .A2(KEYINPUT47), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n811), .A2(KEYINPUT47), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n318), .ZN(G42));
  NAND3_X1  g633(.A1(new_n736), .A2(new_n675), .A3(new_n459), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT113), .Z(new_n821));
  NAND2_X1  g635(.A1(new_n718), .A2(new_n488), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(KEYINPUT49), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n823), .A2(new_n795), .A3(new_n699), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n821), .A2(new_n694), .A3(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT51), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n758), .A2(new_n760), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n675), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n719), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n680), .B1(new_n797), .B2(new_n799), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n745), .A2(new_n748), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n699), .A2(new_n379), .A3(new_n619), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n679), .A2(new_n550), .A3(new_n704), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n694), .A2(new_n675), .A3(new_n719), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n830), .B1(new_n739), .B2(new_n740), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n839), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n836), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n816), .B(new_n817), .C1(new_n459), .C2(new_n822), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n761), .A3(new_n839), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT115), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n826), .B1(new_n847), .B2(KEYINPUT116), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n269), .A2(G952), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n839), .B2(new_n720), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n649), .B2(new_n834), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n754), .A2(new_n756), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n829), .A2(new_n830), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT48), .Z(new_n857));
  NOR3_X1   g671(.A1(new_n853), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n844), .B2(new_n846), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n844), .A2(new_n846), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n863), .B2(new_n859), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n848), .B(new_n858), .C1(new_n864), .C2(new_n826), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n780), .A2(new_n783), .A3(new_n785), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n749), .A2(new_n720), .B1(new_n683), .B2(new_n688), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n669), .A2(new_n681), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n731), .A2(new_n699), .A3(new_n768), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n714), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT52), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n714), .A2(new_n868), .A3(KEYINPUT52), .A4(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n656), .B(new_n379), .C1(new_n630), .C2(new_n632), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n679), .A2(new_n550), .A3(new_n613), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n649), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n317), .A3(new_n878), .A4(new_n508), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n741), .A2(new_n726), .A3(new_n879), .ZN(new_n880));
  AND4_X1   g694(.A1(new_n626), .A2(new_n671), .A3(new_n723), .A4(new_n729), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n712), .B(new_n831), .C1(new_n770), .C2(new_n771), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n611), .A2(new_n612), .A3(new_n681), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n569), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n669), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n883), .B1(new_n569), .B2(new_n884), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n688), .A3(new_n761), .A4(new_n887), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n875), .A2(new_n889), .A3(new_n793), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n866), .B1(new_n867), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n888), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n790), .B2(new_n792), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n786), .A3(KEYINPUT53), .A4(new_n875), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n891), .A2(KEYINPUT54), .A3(new_n894), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n865), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(G952), .A2(G953), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n825), .B1(new_n899), .B2(new_n900), .ZN(G75));
  XNOR2_X1  g715(.A(new_n244), .B(new_n271), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n310), .B1(new_n891), .B2(new_n894), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n904), .A2(G210), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n269), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n905), .A2(KEYINPUT56), .A3(new_n903), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(G51));
  XNOR2_X1  g725(.A(new_n489), .B(KEYINPUT57), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n897), .A2(new_n898), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(new_n487), .B2(new_n484), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n803), .A2(new_n805), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n904), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n907), .B1(new_n914), .B2(new_n916), .ZN(G54));
  AND2_X1   g731(.A1(KEYINPUT58), .A2(G475), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n904), .A2(new_n563), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n563), .B1(new_n904), .B2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n907), .ZN(G60));
  NAND2_X1  g735(.A1(G478), .A2(G902), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT59), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n897), .A2(new_n898), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n644), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n907), .ZN(G63));
  XNOR2_X1  g742(.A(KEYINPUT118), .B(KEYINPUT60), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n371), .A2(new_n310), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n891), .B2(new_n894), .ZN(new_n933));
  INV_X1    g747(.A(new_n374), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n908), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT119), .B(new_n908), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n933), .A2(new_n666), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n939), .A2(KEYINPUT61), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n935), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n895), .A2(new_n931), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n907), .B1(new_n946), .B2(new_n374), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n947), .A2(KEYINPUT120), .A3(KEYINPUT61), .A4(new_n939), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n942), .A2(new_n949), .ZN(G66));
  NAND2_X1  g764(.A1(new_n880), .A2(new_n881), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n269), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT121), .Z(new_n953));
  INV_X1    g767(.A(G224), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n623), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n239), .B(new_n243), .C1(G898), .C2(new_n269), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  NOR2_X1   g772(.A1(new_n403), .A2(new_n406), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n556), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n714), .A2(new_n868), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n702), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n878), .A2(new_n455), .ZN(new_n964));
  OR3_X1    g778(.A1(new_n964), .A2(new_n828), .A3(new_n692), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n813), .A2(new_n818), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n960), .B1(new_n967), .B2(G953), .ZN(new_n968));
  AND4_X1   g782(.A1(new_n691), .A2(new_n811), .A3(new_n731), .A4(new_n855), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  AND4_X1   g784(.A1(new_n793), .A2(new_n966), .A3(new_n961), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n971), .B2(new_n786), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n269), .A2(G900), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n968), .B1(new_n975), .B2(new_n960), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT122), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n976), .B(new_n978), .ZN(G72));
  NOR3_X1   g793(.A1(new_n449), .A2(new_n414), .A3(new_n438), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n951), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n971), .A2(new_n786), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n428), .A2(new_n310), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n695), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n895), .A2(new_n988), .A3(new_n981), .A4(new_n986), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n908), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n963), .A2(new_n982), .A3(new_n965), .A4(new_n966), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n991), .A2(KEYINPUT126), .A3(new_n986), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n986), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n988), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n987), .B(new_n990), .C1(new_n992), .C2(new_n995), .ZN(G57));
endmodule


