//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980;
  NAND2_X1  g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT99), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g005(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT99), .ZN(new_n208));
  XNOR2_X1  g007(.A(G71gat), .B(G78gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G57gat), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n211), .A2(KEYINPUT98), .A3(G64gat), .ZN(new_n212));
  INV_X1    g011(.A(G64gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G57gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT98), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(new_n213), .B2(G57gat), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G71gat), .A2(G78gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G71gat), .A2(G78gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT97), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT97), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n211), .A2(G64gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n207), .B1(new_n214), .B2(new_n224), .ZN(new_n225));
  OAI22_X1  g024(.A1(new_n210), .A2(new_n217), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G127gat), .B(G155gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G183gat), .B(G211gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G231gat), .A2(G233gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT101), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n233), .B(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G22gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G15gat), .ZN(new_n240));
  INV_X1    g039(.A(G15gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G22gat), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT16), .B1(KEYINPUT92), .B2(G1gat), .ZN(new_n243));
  AND2_X1   g042(.A1(KEYINPUT92), .A2(G1gat), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n240), .B(new_n242), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(G1gat), .B1(new_n240), .B2(new_n242), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G15gat), .B(G22gat), .ZN(new_n249));
  NOR3_X1   g048(.A1(new_n249), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n250));
  OAI21_X1  g049(.A(G8gat), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT94), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n247), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT93), .B1(new_n249), .B2(G1gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n245), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT94), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(G8gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n246), .ZN(new_n259));
  INV_X1    g058(.A(G8gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n260), .A3(new_n245), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT95), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n227), .A2(KEYINPUT21), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n238), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n238), .A2(new_n264), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n268), .A3(new_n266), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G85gat), .A2(G92gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT7), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT7), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(G85gat), .A3(G92gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G99gat), .A2(G106gat), .ZN(new_n278));
  INV_X1    g077(.A(G85gat), .ZN(new_n279));
  INV_X1    g078(.A(G92gat), .ZN(new_n280));
  AOI22_X1  g079(.A1(KEYINPUT8), .A2(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G99gat), .B(G106gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(new_n281), .A3(new_n283), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(KEYINPUT91), .A2(G29gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(KEYINPUT91), .A2(G29gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G36gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT14), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(G29gat), .B2(G36gat), .ZN(new_n293));
  INV_X1    g092(.A(G29gat), .ZN(new_n294));
  INV_X1    g093(.A(G36gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT14), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n291), .A2(KEYINPUT15), .A3(new_n293), .A4(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT15), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n295), .B1(new_n288), .B2(new_n289), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n293), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G43gat), .B(G50gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n297), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT17), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n299), .A2(new_n300), .ZN(new_n305));
  INV_X1    g104(.A(new_n302), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT15), .A3(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n304), .B1(new_n303), .B2(new_n307), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n287), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n303), .A2(new_n307), .ZN(new_n311));
  INV_X1    g110(.A(new_n287), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G190gat), .B(G218gat), .Z(new_n316));
  XOR2_X1   g115(.A(new_n315), .B(new_n316), .Z(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G134gat), .B(G162gat), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n319), .B(new_n320), .Z(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n318), .B1(KEYINPUT104), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n321), .B(KEYINPUT104), .Z(new_n324));
  NAND2_X1  g123(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n272), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G230gat), .A2(G233gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n287), .A2(new_n226), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT105), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n215), .A2(new_n213), .A3(G57gat), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT98), .B1(new_n211), .B2(G64gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n211), .A2(G64gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n334), .A2(new_n206), .A3(new_n208), .A4(new_n209), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n214), .A2(new_n224), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n220), .B(new_n222), .C1(new_n336), .C2(new_n207), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n335), .A2(new_n337), .A3(new_n285), .A4(new_n286), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n329), .A2(new_n330), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n312), .A2(new_n227), .A3(KEYINPUT105), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT10), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n328), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n328), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n339), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G120gat), .B(G148gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G176gat), .B(G204gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n346), .A3(new_n350), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n327), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n257), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n256), .B1(new_n255), .B2(G8gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n262), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n311), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n258), .B(new_n262), .C1(new_n308), .C2(new_n309), .ZN(new_n360));
  NAND2_X1  g159(.A1(G229gat), .A2(G233gat), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT18), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G113gat), .B(G141gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(G197gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT11), .B(G169gat), .ZN(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT12), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n258), .A2(new_n262), .A3(new_n303), .A4(new_n307), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n359), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n361), .B(KEYINPUT13), .Z(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT18), .A4(new_n361), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n364), .A2(new_n369), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT96), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n362), .A2(new_n363), .B1(new_n371), .B2(new_n372), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT96), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n369), .A4(new_n374), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n374), .ZN(new_n380));
  INV_X1    g179(.A(new_n369), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n376), .A2(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n355), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(G71gat), .B(G99gat), .Z(new_n384));
  XNOR2_X1  g183(.A(G15gat), .B(G43gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n386), .A2(KEYINPUT68), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(KEYINPUT68), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT33), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(KEYINPUT64), .B(G176gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(G169gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G169gat), .ZN(new_n394));
  INV_X1    g193(.A(G176gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n398), .B2(new_n391), .ZN(new_n399));
  NAND2_X1  g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT24), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G183gat), .ZN(new_n403));
  INV_X1    g202(.A(G190gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n393), .A2(new_n399), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT25), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT65), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT24), .B1(new_n400), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n413), .A2(new_n405), .A3(new_n406), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT25), .B1(new_n396), .B2(new_n391), .ZN(new_n415));
  NOR2_X1   g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(KEYINPUT23), .B2(new_n397), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n408), .A2(new_n409), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT26), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n396), .A2(new_n420), .A3(new_n397), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(KEYINPUT26), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n400), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT27), .B1(new_n403), .B2(KEYINPUT66), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT66), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(G183gat), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n427), .A3(new_n404), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT28), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT27), .B(G183gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT28), .A3(new_n404), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n423), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n419), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G127gat), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT67), .B1(new_n435), .B2(G134gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G113gat), .B(G120gat), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(KEYINPUT1), .ZN(new_n438));
  XNOR2_X1  g237(.A(G127gat), .B(G134gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n439), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n441), .B(new_n436), .C1(KEYINPUT1), .C2(new_n437), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n434), .B(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI211_X1 g245(.A(KEYINPUT32), .B(new_n389), .C1(new_n444), .C2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n444), .A2(new_n446), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n386), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(KEYINPUT33), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n444), .A2(new_n446), .ZN(new_n453));
  XNOR2_X1  g252(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT69), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n444), .A2(new_n456), .A3(KEYINPUT34), .A4(new_n446), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n458), .B(new_n447), .C1(new_n450), .C2(new_n451), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n460), .A2(KEYINPUT36), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT36), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT86), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466));
  NAND2_X1  g265(.A1(G228gat), .A2(G233gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT82), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT3), .ZN(new_n469));
  XNOR2_X1  g268(.A(G155gat), .B(G162gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G141gat), .ZN(new_n472));
  INV_X1    g271(.A(G148gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT2), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(KEYINPUT77), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT77), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT2), .ZN(new_n478));
  NAND2_X1  g277(.A1(G141gat), .A2(G148gat), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n474), .A2(new_n476), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT78), .B(G155gat), .Z(new_n482));
  AOI21_X1  g281(.A(new_n475), .B1(new_n482), .B2(G162gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n470), .A2(new_n474), .A3(new_n479), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n469), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT22), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n488), .A2(KEYINPUT70), .B1(G211gat), .B2(G218gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT22), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G211gat), .B(G218gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(G197gat), .B(G204gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n487), .A2(new_n498), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n470), .A2(new_n474), .A3(new_n479), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT78), .B(G155gat), .ZN(new_n501));
  INV_X1    g300(.A(G162gat), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT2), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n500), .A2(new_n503), .B1(new_n471), .B2(new_n480), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n486), .B1(new_n496), .B2(new_n497), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n469), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT83), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n510));
  INV_X1    g309(.A(new_n493), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT29), .B1(new_n512), .B2(new_n495), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n509), .B1(new_n513), .B2(KEYINPUT3), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n468), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n499), .A2(new_n514), .A3(G228gat), .A4(G233gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n466), .B1(new_n518), .B2(G22gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n516), .A2(new_n239), .A3(new_n517), .ZN(new_n520));
  XNOR2_X1  g319(.A(G78gat), .B(G106gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G50gat), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n521), .B(new_n522), .Z(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n239), .B1(new_n516), .B2(new_n517), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n466), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n516), .A2(new_n239), .A3(new_n517), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n529), .B2(new_n527), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT84), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n526), .A2(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(KEYINPUT84), .B(new_n523), .C1(new_n529), .C2(new_n527), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n465), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n530), .A2(new_n531), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n518), .A2(G22gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT85), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n520), .A2(new_n524), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n537), .A2(new_n538), .A3(new_n528), .ZN(new_n539));
  AND4_X1   g338(.A1(new_n465), .A2(new_n535), .A3(new_n539), .A4(new_n533), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT73), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n430), .A2(new_n432), .ZN(new_n543));
  INV_X1    g342(.A(new_n423), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n417), .B1(new_n390), .B2(new_n392), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT25), .B1(new_n546), .B2(new_n407), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n406), .B1(G183gat), .B2(G190gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n412), .B2(new_n411), .ZN(new_n549));
  NOR3_X1   g348(.A1(new_n549), .A2(new_n417), .A3(new_n415), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n545), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G226gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT71), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n419), .B2(new_n433), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n545), .B(KEYINPUT72), .C1(new_n547), .C2(new_n550), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n553), .A2(new_n486), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n554), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n542), .B1(new_n561), .B2(new_n498), .ZN(new_n562));
  INV_X1    g361(.A(new_n553), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n557), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n551), .A2(new_n560), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n564), .A2(new_n498), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n498), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n559), .B1(new_n556), .B2(new_n557), .ZN(new_n568));
  OAI211_X1 g367(.A(KEYINPUT73), .B(new_n567), .C1(new_n568), .C2(new_n554), .ZN(new_n569));
  XOR2_X1   g368(.A(G8gat), .B(G36gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT75), .ZN(new_n571));
  XNOR2_X1  g370(.A(G64gat), .B(G92gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND4_X1  g372(.A1(new_n562), .A2(new_n566), .A3(new_n569), .A4(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT30), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n560), .ZN(new_n577));
  INV_X1    g376(.A(new_n554), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT73), .B1(new_n579), .B2(new_n567), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n569), .A2(new_n566), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT74), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT74), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n562), .A2(new_n583), .A3(new_n566), .A4(new_n569), .ZN(new_n584));
  INV_X1    g383(.A(new_n573), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n582), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  XNOR2_X1  g387(.A(G1gat), .B(G29gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT0), .ZN(new_n590));
  XNOR2_X1  g389(.A(G57gat), .B(G85gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n590), .B(new_n591), .Z(new_n592));
  XOR2_X1   g391(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n443), .A2(new_n509), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n500), .A2(new_n503), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n595), .A2(new_n440), .A3(new_n481), .A4(new_n442), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G225gat), .A2(G233gat), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n593), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(KEYINPUT4), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT4), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n504), .A2(new_n602), .A3(new_n440), .A4(new_n442), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n485), .A2(new_n443), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n504), .A2(new_n469), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n600), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n485), .A2(new_n443), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n509), .A2(KEYINPUT3), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n599), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(KEYINPUT80), .A3(new_n603), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT80), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n613), .A3(KEYINPUT4), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n611), .A2(new_n612), .A3(new_n593), .A4(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n592), .B1(new_n608), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT6), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT6), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n608), .A2(new_n615), .A3(new_n592), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT81), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n620), .B(new_n621), .C1(new_n616), .C2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n574), .A2(new_n575), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT76), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n576), .A2(new_n586), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n588), .A2(new_n624), .A3(new_n625), .A4(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n464), .B1(new_n541), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n582), .A2(KEYINPUT37), .A3(new_n584), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT87), .B(KEYINPUT37), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n562), .A2(new_n566), .A3(new_n569), .A4(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n632), .A2(new_n585), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT38), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n636), .A2(KEYINPUT37), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n579), .A2(new_n498), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT38), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n639), .A2(new_n632), .A3(KEYINPUT88), .A4(new_n585), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n620), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n574), .B(new_n617), .C1(new_n616), .C2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT88), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n639), .A2(new_n632), .A3(new_n585), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n635), .A2(new_n640), .A3(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n612), .B(new_n614), .C1(new_n606), .C2(new_n605), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n599), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n597), .A2(new_n599), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n650), .A3(new_n599), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n592), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n652), .A2(KEYINPUT40), .A3(new_n592), .A4(new_n653), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n656), .A2(new_n618), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n576), .A2(new_n586), .A3(new_n625), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n658), .A2(new_n659), .B1(new_n532), .B2(new_n533), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n646), .A2(new_n660), .A3(KEYINPUT89), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT89), .B1(new_n646), .B2(new_n660), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n629), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n532), .A2(new_n533), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n460), .A2(new_n461), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT35), .B1(new_n628), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n659), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT35), .B1(new_n670), .B2(new_n617), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n669), .A2(new_n664), .A3(new_n666), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT90), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n665), .B1(new_n533), .B2(new_n532), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT90), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n674), .A2(new_n675), .A3(new_n669), .A4(new_n671), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n668), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n663), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n383), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n624), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g482(.A(new_n260), .B1(new_n680), .B2(new_n659), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT16), .B(G8gat), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n679), .A2(new_n669), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT42), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(KEYINPUT42), .B2(new_n686), .ZN(G1325gat));
  AOI21_X1  g487(.A(G15gat), .B1(new_n680), .B2(new_n666), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n464), .A2(G15gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT106), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n689), .B1(new_n680), .B2(new_n691), .ZN(G1326gat));
  INV_X1    g491(.A(new_n541), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n679), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT43), .B(G22gat), .Z(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n678), .B2(new_n326), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n629), .B(KEYINPUT107), .C1(new_n661), .C2(new_n662), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n658), .A2(new_n659), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(new_n664), .ZN(new_n704));
  INV_X1    g503(.A(new_n642), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n644), .A2(new_n643), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n640), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT38), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n708), .B1(new_n630), .B2(new_n633), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n702), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n646), .A2(new_n660), .A3(KEYINPUT89), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT107), .B1(new_n713), .B2(new_n629), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n677), .B1(new_n701), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n326), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n699), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n272), .ZN(new_n720));
  INV_X1    g519(.A(new_n354), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n382), .A3(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n697), .B1(new_n719), .B2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n718), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n663), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n700), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n728), .B2(new_n677), .ZN(new_n729));
  OAI211_X1 g528(.A(KEYINPUT109), .B(new_n722), .C1(new_n729), .C2(new_n699), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n290), .B1(new_n731), .B2(new_n624), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n678), .A2(new_n326), .A3(new_n722), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n733), .A2(new_n624), .A3(new_n290), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT45), .Z(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(G1328gat));
  OAI21_X1  g535(.A(G36gat), .B1(new_n731), .B2(new_n669), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n733), .A2(G36gat), .A3(new_n669), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT46), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(new_n719), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n722), .ZN(new_n742));
  INV_X1    g541(.A(new_n464), .ZN(new_n743));
  OAI21_X1  g542(.A(G43gat), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n665), .A2(G43gat), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n733), .A2(KEYINPUT110), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT110), .B1(new_n733), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n744), .A2(KEYINPUT47), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n464), .A3(new_n730), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G43gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n749), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT111), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI22_X1  g554(.A1(new_n751), .A2(G43gat), .B1(new_n748), .B2(new_n747), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n756), .A2(new_n757), .A3(KEYINPUT47), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n750), .B1(new_n755), .B2(new_n758), .ZN(G1330gat));
  OAI21_X1  g558(.A(G50gat), .B1(new_n742), .B2(new_n664), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n733), .A2(G50gat), .A3(new_n693), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(KEYINPUT48), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n724), .A2(new_n541), .A3(new_n730), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n764), .A2(KEYINPUT112), .A3(G50gat), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT112), .B1(new_n764), .B2(G50gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n761), .B(KEYINPUT113), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n768), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g568(.A1(new_n715), .A2(new_n382), .A3(new_n327), .A4(new_n721), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n624), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(new_n211), .ZN(G1332gat));
  NOR2_X1   g571(.A1(new_n770), .A2(new_n669), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  AND2_X1   g573(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n773), .B2(new_n774), .ZN(G1333gat));
  OAI21_X1  g576(.A(G71gat), .B1(new_n770), .B2(new_n743), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n665), .A2(G71gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n770), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1334gat));
  NOR2_X1   g581(.A1(new_n770), .A2(new_n693), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(G78gat), .Z(G1335gat));
  INV_X1    g583(.A(new_n382), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n720), .A2(new_n785), .A3(new_n354), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n741), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT115), .B1(new_n787), .B2(new_n624), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G85gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n787), .A2(KEYINPUT115), .A3(new_n624), .ZN(new_n790));
  INV_X1    g589(.A(new_n715), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n272), .A2(new_n382), .A3(new_n326), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(KEYINPUT51), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(KEYINPUT51), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n721), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n681), .A2(new_n279), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n789), .A2(new_n790), .B1(new_n796), .B2(new_n797), .ZN(G1336gat));
  OAI21_X1  g597(.A(G92gat), .B1(new_n787), .B2(new_n669), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n669), .A2(G92gat), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT116), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n796), .B2(new_n801), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT52), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  OAI221_X1 g605(.A(new_n799), .B1(new_n803), .B2(new_n806), .C1(new_n796), .C2(new_n801), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1337gat));
  OAI21_X1  g607(.A(G99gat), .B1(new_n787), .B2(new_n743), .ZN(new_n809));
  OR2_X1    g608(.A1(new_n665), .A2(G99gat), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n796), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(G1338gat));
  NOR2_X1   g612(.A1(new_n664), .A2(G106gat), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n721), .B(new_n814), .C1(new_n794), .C2(new_n795), .ZN(new_n815));
  OAI21_X1  g614(.A(G106gat), .B1(new_n787), .B2(new_n664), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G106gat), .B1(new_n787), .B2(new_n693), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n817), .ZN(G1339gat));
  NAND3_X1  g620(.A1(new_n327), .A2(new_n382), .A3(new_n354), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n339), .A2(new_n340), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n342), .ZN(new_n825));
  INV_X1    g624(.A(new_n343), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n825), .A2(new_n345), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n344), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n328), .C1(new_n341), .C2(new_n343), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n830), .A2(KEYINPUT118), .A3(new_n351), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT118), .B1(new_n830), .B2(new_n351), .ZN(new_n832));
  OAI211_X1 g631(.A(KEYINPUT55), .B(new_n828), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n827), .A2(KEYINPUT54), .A3(new_n344), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n351), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n830), .A2(KEYINPUT118), .A3(new_n351), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n834), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n353), .B(new_n833), .C1(new_n839), .C2(KEYINPUT55), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n382), .ZN(new_n841));
  INV_X1    g640(.A(new_n368), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n361), .B1(new_n359), .B2(new_n360), .ZN(new_n843));
  INV_X1    g642(.A(new_n372), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n359), .A2(new_n370), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n843), .B1(KEYINPUT119), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n845), .A2(KEYINPUT119), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n354), .B(new_n848), .C1(new_n376), .C2(new_n379), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n716), .B1(new_n841), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n840), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n376), .B2(new_n379), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n326), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n720), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n823), .A2(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n855), .A2(new_n681), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n856), .A2(new_n669), .A3(new_n674), .ZN(new_n857));
  AOI21_X1  g656(.A(G113gat), .B1(new_n857), .B2(new_n785), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n855), .A2(new_n693), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n859), .A2(new_n681), .A3(new_n669), .A4(new_n666), .ZN(new_n860));
  INV_X1    g659(.A(G113gat), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n860), .A2(new_n861), .A3(new_n382), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n858), .A2(new_n862), .ZN(G1340gat));
  AOI21_X1  g662(.A(G120gat), .B1(new_n857), .B2(new_n721), .ZN(new_n864));
  INV_X1    g663(.A(G120gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n860), .A2(new_n865), .A3(new_n354), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(G1341gat));
  NAND3_X1  g666(.A1(new_n857), .A2(new_n435), .A3(new_n720), .ZN(new_n868));
  OAI21_X1  g667(.A(G127gat), .B1(new_n860), .B2(new_n272), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(G1342gat));
  INV_X1    g669(.A(G134gat), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n857), .A2(new_n871), .A3(new_n326), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  OAI21_X1  g672(.A(G134gat), .B1(new_n860), .B2(new_n716), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n464), .A2(new_n624), .A3(new_n659), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n664), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n855), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g679(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n382), .B1(new_n840), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n837), .A2(new_n838), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n834), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n833), .A2(new_n353), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT121), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n849), .B1(new_n884), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n716), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT122), .B(new_n849), .C1(new_n884), .C2(new_n890), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n853), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(new_n272), .ZN(new_n896));
  OAI211_X1 g695(.A(KEYINPUT57), .B(new_n541), .C1(new_n896), .C2(new_n823), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n878), .B1(new_n882), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n472), .B1(new_n898), .B2(new_n785), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n464), .A2(new_n664), .A3(new_n659), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n856), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n472), .A3(new_n785), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n904), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT58), .B1(new_n906), .B2(new_n899), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1344gat));
  NAND3_X1  g707(.A1(new_n903), .A2(new_n473), .A3(new_n721), .ZN(new_n909));
  AOI211_X1 g708(.A(KEYINPUT59), .B(new_n473), .C1(new_n898), .C2(new_n721), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  INV_X1    g710(.A(new_n881), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n879), .B(new_n912), .C1(new_n823), .C2(new_n854), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n895), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(KEYINPUT123), .B(new_n853), .C1(new_n893), .C2(new_n894), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n272), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n693), .B1(new_n917), .B2(new_n822), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n913), .B1(new_n918), .B2(KEYINPUT57), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n721), .A3(new_n877), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n911), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n909), .B1(new_n910), .B2(new_n921), .ZN(G1345gat));
  INV_X1    g721(.A(new_n898), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n482), .B1(new_n923), .B2(new_n272), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n903), .A2(new_n501), .A3(new_n720), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1346gat));
  AOI21_X1  g725(.A(G162gat), .B1(new_n903), .B2(new_n326), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n716), .A2(new_n502), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n898), .B2(new_n928), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n669), .A2(new_n681), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n855), .A2(new_n674), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n394), .A3(new_n785), .ZN(new_n932));
  INV_X1    g731(.A(new_n930), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n665), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n859), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G169gat), .B1(new_n935), .B2(new_n382), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n932), .B1(new_n938), .B2(new_n939), .ZN(G1348gat));
  NOR3_X1   g739(.A1(new_n935), .A2(new_n390), .A3(new_n354), .ZN(new_n941));
  AOI21_X1  g740(.A(G176gat), .B1(new_n931), .B2(new_n721), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(G1349gat));
  OAI21_X1  g742(.A(G183gat), .B1(new_n935), .B2(new_n272), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n931), .A2(new_n431), .A3(new_n720), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n404), .A3(new_n326), .ZN(new_n948));
  OAI21_X1  g747(.A(G190gat), .B1(new_n935), .B2(new_n716), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NOR2_X1   g751(.A1(new_n933), .A2(new_n464), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n880), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(G197gat), .B1(new_n955), .B2(new_n785), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n953), .B(KEYINPUT125), .Z(new_n957));
  AND2_X1   g756(.A1(new_n919), .A2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n785), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  INV_X1    g759(.A(G204gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n955), .A2(new_n961), .A3(new_n721), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT62), .Z(new_n963));
  AND2_X1   g762(.A1(new_n958), .A2(new_n721), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n964), .B2(new_n961), .ZN(G1353gat));
  INV_X1    g764(.A(G211gat), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n954), .A2(new_n272), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n855), .A2(new_n966), .A3(new_n879), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n919), .A2(new_n967), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT63), .ZN(new_n971));
  AOI211_X1 g770(.A(new_n971), .B(new_n966), .C1(new_n919), .C2(new_n967), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g774(.A(KEYINPUT126), .B(new_n968), .C1(new_n970), .C2(new_n972), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1354gat));
  INV_X1    g776(.A(G218gat), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n955), .A2(new_n978), .A3(new_n326), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n958), .A2(new_n326), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n978), .ZN(G1355gat));
endmodule


