//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  AND2_X1   g000(.A1(KEYINPUT68), .A2(G953), .ZN(new_n187));
  NOR2_X1   g001(.A1(KEYINPUT68), .A2(G953), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G210), .A3(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G116), .B(G119), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT2), .B(G113), .Z(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n195), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  OR2_X1    g017(.A1(KEYINPUT64), .A2(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT64), .A2(G134), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G137), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n203), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n204), .A2(G137), .A3(new_n205), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n209), .A2(G137), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT11), .B1(new_n206), .B2(new_n207), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n211), .B1(new_n218), .B2(new_n203), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n220), .A2(new_n221), .A3(G128), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G143), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n224), .B(G146), .C1(new_n226), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n230));
  INV_X1    g044(.A(G128), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n224), .A2(G146), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n231), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n229), .A2(new_n230), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n230), .B1(new_n229), .B2(new_n235), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n223), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n219), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n240));
  AND2_X1   g054(.A1(KEYINPUT64), .A2(G134), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT64), .A2(G134), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n212), .B1(new_n243), .B2(G137), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n214), .B1(new_n243), .B2(G137), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n203), .B(new_n244), .C1(new_n245), .C2(new_n212), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n220), .ZN(new_n248));
  NAND2_X1  g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n220), .A2(KEYINPUT0), .A3(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n202), .B1(new_n239), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n208), .A2(new_n210), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G131), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n246), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n260), .A2(new_n261), .B1(G143), .B2(new_n233), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT66), .B(new_n248), .C1(new_n262), .C2(new_n231), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n229), .A2(new_n230), .A3(new_n235), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n222), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n201), .B(KEYINPUT67), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n253), .B1(new_n240), .B2(new_n246), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n256), .B1(new_n269), .B2(KEYINPUT28), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n201), .B(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n239), .A2(new_n255), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n194), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n266), .A2(KEYINPUT30), .A3(new_n268), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT30), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n239), .B2(new_n255), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n201), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(new_n194), .A3(new_n273), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT30), .B1(new_n266), .B2(new_n268), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n239), .A2(new_n255), .A3(new_n278), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n269), .B1(new_n286), .B2(new_n201), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT31), .A3(new_n194), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n276), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT32), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  XOR2_X1   g107(.A(KEYINPUT69), .B(KEYINPUT32), .Z(new_n294));
  INV_X1    g108(.A(new_n276), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT31), .B1(new_n287), .B2(new_n194), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n202), .B1(new_n284), .B2(new_n285), .ZN(new_n297));
  INV_X1    g111(.A(new_n194), .ZN(new_n298));
  NOR4_X1   g112(.A1(new_n297), .A2(new_n282), .A3(new_n298), .A4(new_n269), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n295), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n294), .B1(new_n300), .B2(new_n291), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n270), .A2(new_n194), .A3(new_n275), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n298), .B1(new_n297), .B2(new_n269), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n272), .B1(new_n239), .B2(new_n255), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT28), .B1(new_n269), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT70), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n273), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT70), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT28), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n275), .A2(KEYINPUT71), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT71), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n273), .A2(new_n316), .A3(new_n274), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n298), .A2(new_n305), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(G902), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n306), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n312), .B1(new_n311), .B2(KEYINPUT28), .ZN(new_n324));
  AOI211_X1 g138(.A(KEYINPUT70), .B(new_n274), .C1(new_n310), .C2(new_n273), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT72), .ZN(new_n329));
  OAI21_X1  g143(.A(G472), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n302), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G110), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n231), .A2(G119), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT74), .ZN(new_n334));
  INV_X1    g148(.A(G119), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n334), .A2(KEYINPUT23), .B1(new_n335), .B2(G128), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(KEYINPUT74), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n332), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n335), .A2(G128), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n343), .A2(KEYINPUT73), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(KEYINPUT73), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G140), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(KEYINPUT75), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT75), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(G125), .A3(G140), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(KEYINPUT16), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT16), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(new_n348), .B2(G140), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n352), .A2(new_n233), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n233), .B1(new_n352), .B2(new_n354), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(new_n338), .A3(new_n332), .A4(new_n340), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n341), .A2(new_n342), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n336), .A2(KEYINPUT76), .A3(new_n332), .A4(new_n338), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G125), .B(G140), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n356), .B1(new_n233), .B2(new_n366), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n346), .A2(new_n358), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G137), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(KEYINPUT77), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n346), .A2(new_n358), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n365), .A2(new_n367), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n372), .ZN(new_n377));
  INV_X1    g191(.A(G217), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n378), .B1(G234), .B2(new_n323), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G902), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n374), .A2(KEYINPUT25), .A3(new_n323), .A4(new_n377), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n372), .B(KEYINPUT77), .Z(new_n384));
  OAI211_X1 g198(.A(new_n323), .B(new_n377), .C1(new_n384), .C2(new_n368), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n382), .B1(new_n388), .B2(new_n379), .ZN(new_n389));
  XOR2_X1   g203(.A(new_n389), .B(KEYINPUT78), .Z(new_n390));
  NAND2_X1  g204(.A1(new_n331), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT20), .ZN(new_n392));
  NOR2_X1   g206(.A1(G475), .A2(G902), .ZN(new_n393));
  OR2_X1    g207(.A1(KEYINPUT68), .A2(G953), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT68), .A2(G953), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n394), .A2(G214), .A3(new_n190), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n224), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n189), .A2(G143), .A3(G214), .A4(new_n190), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT18), .A3(G131), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n366), .A2(new_n233), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n349), .A2(G146), .A3(new_n351), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT18), .A2(G131), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n397), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT87), .B(G104), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n407), .B(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n399), .A2(G131), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n397), .A2(new_n398), .A3(new_n203), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n357), .B1(new_n410), .B2(new_n411), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n406), .B(new_n409), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n410), .A2(new_n412), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n366), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n349), .A2(KEYINPUT19), .A3(new_n351), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n233), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT86), .B1(new_n422), .B2(new_n356), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n352), .A2(new_n354), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n424), .B(new_n421), .C1(new_n425), .C2(new_n233), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n417), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n409), .B1(new_n427), .B2(new_n406), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n392), .B(new_n393), .C1(new_n416), .C2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n393), .ZN(new_n430));
  OAI21_X1  g244(.A(KEYINPUT88), .B1(new_n416), .B2(new_n428), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n427), .A2(new_n406), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n432), .B(new_n415), .C1(new_n433), .C2(new_n409), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n430), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n429), .B1(new_n435), .B2(new_n392), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n406), .B1(new_n413), .B2(new_n414), .ZN(new_n437));
  INV_X1    g251(.A(new_n409), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n439), .A2(new_n415), .ZN(new_n440));
  OAI21_X1  g254(.A(G475), .B1(new_n440), .B2(G902), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT9), .B(G234), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n443), .A2(new_n378), .A3(G953), .ZN(new_n444));
  XNOR2_X1  g258(.A(G116), .B(G122), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G122), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G116), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n448), .A2(KEYINPUT14), .ZN(new_n449));
  INV_X1    g263(.A(G107), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(KEYINPUT14), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n452), .A3(G107), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n224), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n231), .A2(G143), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n455), .B2(new_n456), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n459), .A2(new_n206), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n455), .A2(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT90), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n243), .B1(new_n463), .B2(new_n458), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n454), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n206), .B1(new_n459), .B2(new_n460), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n458), .A3(new_n243), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(KEYINPUT91), .A3(new_n454), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(G128), .A3(new_n224), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(G134), .C1(new_n462), .C2(new_n473), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n445), .B(new_n450), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(new_n469), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n444), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n444), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n480), .B(new_n477), .C1(new_n467), .C2(new_n471), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n323), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G478), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(KEYINPUT15), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n470), .A2(KEYINPUT91), .A3(new_n454), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT91), .B1(new_n470), .B2(new_n454), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n478), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n480), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n472), .A2(new_n478), .A3(new_n444), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n484), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI211_X1 g307(.A(new_n323), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT21), .B(G898), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT92), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G953), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G952), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(G234), .B2(G237), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n485), .A2(new_n493), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT93), .B1(new_n442), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n504), .A2(new_n436), .A3(new_n507), .A4(new_n441), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G210), .B1(G237), .B2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n265), .A2(new_n348), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n253), .A2(G125), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G224), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(G953), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n516), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n512), .B2(new_n513), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n195), .A2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT5), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n522), .A2(new_n335), .A3(G116), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT83), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n522), .A2(new_n335), .A3(KEYINPUT83), .A4(G116), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n521), .A2(G113), .A3(new_n525), .A4(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT80), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n450), .A3(G104), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT3), .ZN(new_n530));
  INV_X1    g344(.A(G101), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT3), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n528), .A2(new_n532), .A3(new_n450), .A4(G104), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n450), .A2(G104), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n530), .A2(new_n531), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(G104), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G107), .ZN(new_n538));
  OAI21_X1  g352(.A(G101), .B1(new_n538), .B2(new_n534), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n527), .A2(new_n200), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G110), .B(G122), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n530), .A2(new_n533), .A3(new_n535), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT81), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT4), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT81), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n530), .A2(new_n545), .A3(new_n533), .A4(new_n535), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n543), .A2(new_n544), .A3(G101), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n201), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n536), .A2(KEYINPUT4), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n531), .B1(new_n542), .B2(KEYINPUT81), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(new_n546), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n540), .B(new_n541), .C1(new_n548), .C2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n540), .B1(new_n548), .B2(new_n551), .ZN(new_n555));
  INV_X1    g369(.A(new_n541), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n556), .A3(new_n553), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n520), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n541), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n540), .A2(KEYINPUT85), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n527), .A2(new_n200), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n536), .A2(new_n539), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n540), .A2(KEYINPUT85), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n561), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n514), .B1(new_n569), .B2(new_n516), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n512), .A2(KEYINPUT7), .A3(new_n518), .A4(new_n513), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n568), .A2(new_n570), .A3(new_n552), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n323), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n511), .B1(new_n560), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n560), .A2(new_n573), .A3(new_n511), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G214), .B1(G237), .B2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G221), .B1(new_n443), .B2(G902), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n581), .B(KEYINPUT79), .Z(new_n582));
  INV_X1    g396(.A(G469), .ZN(new_n583));
  OAI21_X1  g397(.A(KEYINPUT10), .B1(new_n265), .B2(new_n564), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n234), .A2(KEYINPUT1), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n220), .B2(G128), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n536), .B(new_n539), .C1(new_n222), .C2(new_n586), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n587), .A2(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n247), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n543), .A2(G101), .A3(new_n546), .ZN(new_n591));
  INV_X1    g405(.A(new_n549), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n254), .A3(new_n547), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n189), .A2(G227), .ZN(new_n596));
  XOR2_X1   g410(.A(G110), .B(G140), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n223), .B(new_n564), .C1(new_n236), .C2(new_n237), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n587), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n602), .A2(new_n247), .A3(KEYINPUT12), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT12), .B1(new_n602), .B2(new_n247), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g421(.A(new_n564), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n238), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n587), .A2(KEYINPUT10), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n594), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n247), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n599), .B1(new_n612), .B2(new_n595), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n583), .B(new_n323), .C1(new_n606), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT82), .ZN(new_n615));
  INV_X1    g429(.A(new_n595), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n590), .B1(new_n589), .B2(new_n594), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n598), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n595), .B(new_n599), .C1(new_n603), .C2(new_n604), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT82), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n620), .A2(new_n621), .A3(new_n583), .A4(new_n323), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n595), .B1(new_n603), .B2(new_n604), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n598), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n612), .A2(new_n595), .A3(new_n599), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n583), .B1(new_n627), .B2(new_n323), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n582), .B1(new_n623), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n509), .A2(new_n580), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n391), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n531), .ZN(G3));
  INV_X1    g447(.A(G472), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n300), .B2(new_n323), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n289), .A2(new_n292), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n390), .A2(new_n630), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT96), .B(G478), .Z(new_n640));
  OAI21_X1  g454(.A(KEYINPUT97), .B1(new_n491), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT97), .ZN(new_n642));
  INV_X1    g456(.A(new_n640), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n482), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT95), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT33), .B1(new_n479), .B2(new_n481), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n489), .A2(new_n648), .A3(new_n490), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n483), .A2(G902), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n651), .ZN(new_n653));
  AOI211_X1 g467(.A(KEYINPUT95), .B(new_n653), .C1(new_n647), .C2(new_n649), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n645), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g469(.A1(new_n655), .A2(new_n442), .A3(new_n502), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n579), .B1(new_n576), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n558), .A2(new_n559), .ZN(new_n659));
  INV_X1    g473(.A(new_n520), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(new_n323), .A3(new_n572), .A4(new_n510), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(KEYINPUT94), .A3(new_n574), .ZN(new_n663));
  AND2_X1   g477(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT98), .B1(new_n656), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n655), .A2(new_n442), .A3(new_n502), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n658), .A2(new_n663), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n639), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT99), .Z(new_n671));
  XOR2_X1   g485(.A(KEYINPUT34), .B(G104), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G6));
  XNOR2_X1  g487(.A(new_n435), .B(new_n392), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n675), .B(G475), .C1(new_n440), .C2(G902), .ZN(new_n676));
  AOI21_X1  g490(.A(G902), .B1(new_n439), .B2(new_n415), .ZN(new_n677));
  INV_X1    g491(.A(G475), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT100), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n485), .A2(new_n493), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n502), .B(KEYINPUT101), .Z(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n667), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n639), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT35), .B(G107), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G9));
  NAND2_X1  g503(.A1(new_n388), .A2(new_n379), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n373), .A2(KEYINPUT36), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n369), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n380), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n635), .A2(new_n636), .A3(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n509), .A2(new_n696), .A3(new_n580), .A4(new_n630), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT37), .B(G110), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G12));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n701), .B1(new_n328), .B2(KEYINPUT72), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n320), .A2(new_n321), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n634), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n294), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n289), .B2(new_n292), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n300), .A2(KEYINPUT32), .A3(new_n291), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n630), .B(new_n694), .C1(new_n704), .C2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(G900), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n494), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT102), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT102), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n712), .A2(new_n501), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n674), .A2(new_n682), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n664), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n700), .B1(new_n709), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n695), .B1(new_n302), .B2(new_n330), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n716), .A2(new_n667), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(KEYINPUT103), .A3(new_n630), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G128), .ZN(G30));
  XNOR2_X1  g538(.A(new_n577), .B(KEYINPUT38), .ZN(new_n725));
  INV_X1    g539(.A(new_n681), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n442), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n725), .A2(new_n579), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n311), .A2(new_n298), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n281), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(G472), .B1(new_n730), .B2(G902), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n706), .A2(new_n707), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(new_n695), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(new_n714), .B(KEYINPUT39), .Z(new_n734));
  NAND2_X1  g548(.A1(new_n630), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n735), .A2(KEYINPUT40), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(KEYINPUT40), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n224), .ZN(G45));
  NAND3_X1  g553(.A1(new_n655), .A2(new_n442), .A3(new_n715), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n667), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n331), .A2(new_n630), .A3(new_n694), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G146), .ZN(G48));
  XNOR2_X1  g557(.A(new_n389), .B(KEYINPUT78), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n302), .B2(new_n330), .ZN(new_n745));
  INV_X1    g559(.A(new_n582), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n620), .A2(new_n323), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n623), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n745), .B(new_n750), .C1(new_n665), .C2(new_n669), .ZN(new_n751));
  XNOR2_X1  g565(.A(KEYINPUT41), .B(G113), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT104), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n751), .B(new_n753), .ZN(G15));
  NAND3_X1  g568(.A1(new_n745), .A2(new_n686), .A3(new_n750), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT105), .B(G116), .Z(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G18));
  NOR2_X1   g571(.A1(new_n749), .A2(new_n667), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n720), .A2(new_n509), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  NAND2_X1  g574(.A1(new_n283), .A2(new_n288), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n315), .A2(new_n317), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n313), .B2(new_n309), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n298), .B1(new_n763), .B2(KEYINPUT106), .ZN(new_n764));
  INV_X1    g578(.A(new_n762), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n314), .A2(new_n765), .A3(KEYINPUT106), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n761), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n635), .B1(new_n768), .B2(new_n291), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n727), .A2(new_n685), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n758), .A2(new_n769), .A3(new_n389), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G122), .ZN(G24));
  NAND4_X1  g586(.A1(new_n741), .A2(new_n769), .A3(new_n750), .A4(new_n694), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  AOI21_X1  g588(.A(new_n628), .B1(new_n615), .B2(new_n622), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n662), .A2(new_n578), .A3(new_n574), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n582), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n740), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n331), .A2(new_n390), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n389), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT32), .B1(new_n300), .B2(new_n291), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n293), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n782), .B1(new_n784), .B2(new_n330), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(KEYINPUT42), .A3(new_n778), .A4(new_n777), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT108), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n781), .A2(new_n789), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT109), .B(G131), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(G33));
  NAND3_X1  g607(.A1(new_n745), .A2(new_n717), .A3(new_n777), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G134), .ZN(G36));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n436), .A2(new_n441), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n655), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n798), .B2(KEYINPUT110), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n798), .B2(new_n796), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(KEYINPUT43), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n637), .A2(new_n695), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT44), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n625), .A2(new_n626), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(KEYINPUT45), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(KEYINPUT45), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(G469), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(G469), .A2(G902), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT46), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n623), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n810), .A2(KEYINPUT46), .A3(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n746), .A3(new_n734), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n806), .A2(new_n776), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n804), .A2(KEYINPUT44), .A3(new_n805), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G137), .ZN(G39));
  OR4_X1    g635(.A1(new_n331), .A2(new_n390), .A3(new_n740), .A4(new_n776), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n816), .A2(new_n746), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT47), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n816), .A2(KEYINPUT47), .A3(new_n746), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(new_n347), .ZN(G42));
  INV_X1    g642(.A(new_n776), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n750), .A2(new_n829), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n501), .B(new_n830), .C1(new_n802), .C2(new_n803), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n785), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT48), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n834), .A3(new_n785), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n390), .A2(new_n500), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n830), .A2(new_n837), .A3(new_n732), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n655), .A2(new_n442), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n501), .B1(new_n802), .B2(new_n803), .ZN(new_n842));
  INV_X1    g656(.A(new_n769), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n782), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n499), .B(new_n841), .C1(new_n845), .C2(new_n758), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n623), .A2(new_n582), .A3(new_n748), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n825), .A2(new_n826), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n829), .A3(new_n845), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n843), .A2(new_n695), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n655), .A2(new_n442), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n838), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT115), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n838), .A2(new_n854), .A3(new_n851), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n831), .A2(new_n850), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n849), .A2(KEYINPUT51), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n725), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n858), .A2(new_n578), .A3(new_n749), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n842), .A2(new_n844), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT50), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n836), .B(new_n846), .C1(new_n857), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n845), .A2(KEYINPUT50), .A3(new_n859), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n860), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n849), .A2(new_n856), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n864), .A2(KEYINPUT114), .A3(new_n866), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n862), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n726), .A2(new_n680), .A3(new_n714), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n874), .A2(new_n674), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n720), .A2(new_n777), .A3(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n777), .A2(new_n769), .A3(new_n694), .A4(new_n778), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n794), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n578), .B(new_n684), .C1(new_n575), .C2(new_n576), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n726), .A2(new_n436), .A3(new_n441), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n879), .B1(new_n839), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n390), .A3(new_n630), .A4(new_n637), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n697), .C1(new_n391), .C2(new_n631), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n751), .A2(new_n755), .A3(new_n759), .A4(new_n771), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n788), .A2(new_n884), .A3(new_n885), .A4(new_n790), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n775), .A2(new_n582), .A3(new_n714), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n667), .A2(new_n727), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n887), .A2(new_n888), .A3(new_n695), .A4(new_n732), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n742), .A2(new_n773), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n723), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT52), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n723), .A3(KEYINPUT52), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n886), .A2(KEYINPUT53), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n890), .A2(KEYINPUT52), .A3(new_n723), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT52), .B1(new_n890), .B2(new_n723), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n788), .A2(new_n884), .A3(new_n885), .A4(new_n790), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n896), .A2(new_n902), .A3(KEYINPUT113), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT113), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n904), .B(new_n897), .C1(new_n900), .C2(new_n901), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(KEYINPUT54), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n897), .B1(new_n781), .B2(new_n786), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n884), .A2(new_n885), .A3(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n895), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n902), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n873), .A2(new_n906), .A3(new_n912), .ZN(new_n913));
  OR2_X1    g727(.A1(G952), .A2(G953), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n623), .A2(new_n748), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n916), .A2(KEYINPUT49), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT112), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n389), .A2(new_n578), .A3(new_n746), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n732), .A2(new_n798), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n858), .B1(KEYINPUT49), .B2(new_n916), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n915), .A2(new_n922), .ZN(G75));
  NOR2_X1   g737(.A1(new_n189), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT53), .B1(new_n886), .B2(new_n895), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n900), .A2(new_n909), .ZN(new_n927));
  OAI211_X1 g741(.A(G210), .B(G902), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n659), .A2(new_n660), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n560), .ZN(new_n932));
  XNOR2_X1  g746(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n925), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT118), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n929), .A2(KEYINPUT117), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n929), .A2(KEYINPUT117), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n928), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n936), .B1(new_n928), .B2(new_n939), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n935), .A2(new_n942), .ZN(G51));
  OAI21_X1  g757(.A(new_n907), .B1(new_n900), .B2(new_n909), .ZN(new_n944));
  OAI21_X1  g758(.A(KEYINPUT119), .B1(new_n926), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT54), .B1(new_n926), .B2(new_n927), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT119), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n902), .A2(new_n947), .A3(new_n907), .A4(new_n911), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n811), .B(KEYINPUT57), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n620), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n902), .A2(new_n911), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(G902), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(new_n810), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n924), .B1(new_n952), .B2(new_n955), .ZN(G54));
  NAND2_X1  g770(.A1(new_n431), .A2(new_n434), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(KEYINPUT58), .A2(G475), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n925), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n650), .B(KEYINPUT120), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n949), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n925), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n906), .A2(new_n912), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n969), .B2(new_n965), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n926), .B2(new_n927), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n374), .A2(new_n377), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n924), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND4_X1   g791(.A1(KEYINPUT121), .A2(new_n953), .A3(new_n692), .A4(new_n974), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n973), .B1(new_n902), .B2(new_n911), .ZN(new_n979));
  AOI21_X1  g793(.A(KEYINPUT121), .B1(new_n979), .B2(new_n692), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(KEYINPUT61), .B(new_n977), .C1(new_n978), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G66));
  OAI21_X1  g799(.A(G953), .B1(new_n496), .B2(new_n515), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n751), .A2(new_n755), .A3(new_n759), .A4(new_n771), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n883), .ZN(new_n988));
  INV_X1    g802(.A(new_n189), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n558), .B(new_n559), .C1(G898), .C2(new_n189), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT122), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(G69));
  NAND2_X1  g807(.A1(new_n419), .A2(new_n420), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n286), .B(new_n994), .Z(new_n995));
  AND2_X1   g809(.A1(new_n995), .A2(KEYINPUT124), .ZN(new_n996));
  OAI21_X1  g810(.A(G900), .B1(new_n996), .B2(G227), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n989), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n995), .B1(G227), .B2(new_n189), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n827), .B1(new_n818), .B2(new_n819), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n723), .A2(new_n742), .A3(new_n773), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT123), .Z(new_n1002));
  NAND2_X1  g816(.A1(new_n785), .A2(new_n888), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n794), .B1(new_n817), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n791), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1000), .A2(new_n1002), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n999), .B1(new_n1006), .B2(new_n189), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n839), .A2(new_n880), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n745), .A2(new_n829), .A3(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1000), .B1(new_n735), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n738), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1002), .A2(KEYINPUT62), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT62), .B1(new_n1002), .B2(new_n1012), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n995), .A2(new_n989), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT124), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n998), .B1(new_n1017), .B2(new_n1018), .ZN(G72));
  XNOR2_X1  g833(.A(new_n287), .B(KEYINPUT125), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n194), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n1011), .B(new_n988), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  AOI21_X1  g838(.A(new_n1021), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n988), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1024), .B1(new_n1006), .B2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1020), .A2(new_n194), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT126), .Z(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n281), .A2(new_n304), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n903), .A2(new_n905), .A3(new_n1024), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1030), .A2(new_n925), .A3(new_n1032), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1025), .A2(new_n1033), .ZN(G57));
endmodule


