//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n194), .A2(new_n197), .A3(new_n201), .A4(new_n198), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(KEYINPUT4), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n204), .A3(G101), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT0), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT64), .B1(new_n213), .B2(G143), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n211), .A3(G146), .ZN(new_n216));
  AOI211_X1 g030(.A(new_n209), .B(new_n212), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT0), .B1(new_n208), .B2(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n210), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n196), .A2(G104), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n193), .A2(G107), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n202), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n202), .B2(new_n222), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT10), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n214), .A2(new_n216), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n213), .A2(G143), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n228), .A2(new_n229), .A3(G128), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n211), .B2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n211), .A2(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n227), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n206), .A2(new_n219), .B1(new_n226), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n239));
  OAI211_X1 g053(.A(KEYINPUT79), .B(KEYINPUT1), .C1(new_n211), .C2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G128), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT79), .B1(new_n230), .B2(KEYINPUT1), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n231), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n202), .A2(new_n222), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n239), .B1(new_n248), .B2(new_n227), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n214), .A2(new_n216), .ZN(new_n250));
  OAI22_X1  g064(.A1(new_n250), .A2(new_n212), .B1(new_n241), .B2(new_n242), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n246), .B1(new_n251), .B2(new_n231), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n252), .A2(KEYINPUT80), .A3(KEYINPUT10), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n238), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT11), .A3(G134), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(G137), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n259), .A3(new_n263), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n254), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT83), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n219), .A2(new_n205), .A3(new_n203), .ZN(new_n273));
  INV_X1    g087(.A(new_n225), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n202), .A2(new_n222), .A3(new_n223), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n237), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT80), .B1(new_n252), .B2(KEYINPUT10), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT79), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n232), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(G128), .A3(new_n240), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n228), .A2(new_n230), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n217), .A2(new_n229), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n239), .B(new_n227), .C1(new_n283), .C2(new_n246), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n277), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT82), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n270), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n284), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n288), .A2(new_n286), .A3(new_n238), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n272), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n269), .B1(new_n254), .B2(KEYINPUT82), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n285), .A2(new_n286), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(KEYINPUT83), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n271), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g108(.A(G110), .B(G140), .ZN(new_n295));
  INV_X1    g109(.A(G953), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n296), .A2(G227), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n295), .B(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n192), .B1(new_n294), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n271), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n286), .B1(new_n288), .B2(new_n238), .ZN(new_n302));
  NOR4_X1   g116(.A1(new_n289), .A2(new_n302), .A3(new_n272), .A4(new_n269), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT83), .B1(new_n291), .B2(new_n292), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(KEYINPUT84), .A3(new_n298), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n271), .A2(new_n298), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n231), .A2(new_n236), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n248), .B1(new_n308), .B2(new_n247), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT12), .A3(new_n265), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n309), .A2(new_n270), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(KEYINPUT12), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n300), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G469), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT74), .B(G902), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n315), .A2(new_n190), .ZN(new_n318));
  INV_X1    g132(.A(new_n307), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n290), .B2(new_n293), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n299), .B1(new_n301), .B2(new_n312), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(G469), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n191), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n219), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G125), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n308), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT86), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT86), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n331), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G224), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n274), .A2(new_n275), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT66), .B(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G116), .ZN(new_n340));
  INV_X1    g154(.A(G116), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(KEYINPUT5), .A3(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n343), .B(G113), .C1(KEYINPUT5), .C2(new_n340), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT2), .B(G113), .Z(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n345), .A3(new_n342), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n345), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n340), .A2(new_n342), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g165(.A(KEYINPUT65), .B(new_n345), .C1(new_n340), .C2(new_n342), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n203), .A2(new_n205), .ZN(new_n354));
  OAI22_X1  g168(.A1(new_n338), .A2(new_n347), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n337), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n206), .B1(new_n352), .B2(new_n351), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n358), .B(KEYINPUT85), .C1(new_n338), .C2(new_n347), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n358), .B(new_n337), .C1(new_n338), .C2(new_n347), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n357), .A2(new_n359), .B1(new_n361), .B2(KEYINPUT6), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n336), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G210), .B1(G237), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT87), .ZN(new_n366));
  INV_X1    g180(.A(new_n335), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT7), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n326), .A2(new_n328), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n329), .A2(KEYINPUT7), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n347), .A2(new_n247), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n344), .A2(new_n246), .A3(new_n346), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n337), .B(KEYINPUT8), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n361), .A2(new_n369), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n190), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n363), .A2(new_n366), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n366), .B1(new_n363), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n325), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G125), .B(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT16), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT16), .ZN(new_n384));
  INV_X1    g198(.A(G140), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G125), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(G146), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(G146), .B1(new_n383), .B2(new_n386), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(G237), .A2(G953), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT88), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(new_n211), .ZN(new_n393));
  NOR2_X1   g207(.A1(KEYINPUT88), .A2(G143), .ZN(new_n394));
  OAI211_X1 g208(.A(G214), .B(new_n391), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(G214), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n392), .B2(new_n211), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n263), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n397), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(G131), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n390), .B(new_n399), .C1(new_n401), .C2(KEYINPUT17), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT91), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n193), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n382), .A2(new_n213), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n382), .B(KEYINPUT89), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(new_n213), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(KEYINPUT18), .ZN(new_n409));
  NAND2_X1  g223(.A1(KEYINPUT18), .A2(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n395), .A2(new_n397), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n402), .A2(new_n403), .A3(new_n405), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n390), .A2(new_n399), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n400), .A2(G131), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n398), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n405), .B(new_n412), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT91), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n382), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n213), .B(new_n420), .C1(new_n407), .C2(new_n419), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT90), .A3(new_n387), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n401), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT90), .B1(new_n421), .B2(new_n387), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n412), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n405), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n413), .A2(new_n418), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT92), .Z(new_n429));
  OAI21_X1  g243(.A(KEYINPUT20), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n425), .A2(new_n426), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n418), .A2(new_n413), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  INV_X1    g248(.A(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n402), .A2(new_n412), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n405), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n190), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n430), .A2(new_n436), .B1(new_n439), .B2(G475), .ZN(new_n440));
  INV_X1    g254(.A(G122), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G116), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n341), .A2(G122), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(KEYINPUT95), .A3(KEYINPUT14), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT95), .B1(new_n443), .B2(KEYINPUT14), .ZN(new_n446));
  OAI221_X1 g260(.A(new_n442), .B1(KEYINPUT14), .B2(new_n443), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G107), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n443), .A2(new_n442), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT93), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n196), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n211), .A2(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n209), .A2(G143), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT94), .ZN(new_n455));
  XNOR2_X1  g269(.A(G128), .B(G143), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT94), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n256), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n458), .A3(G134), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n448), .A2(new_n451), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT96), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n449), .A2(KEYINPUT93), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n449), .A2(KEYINPUT93), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(G107), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n451), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n452), .A2(KEYINPUT13), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(new_n256), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n456), .A2(KEYINPUT13), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n460), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT96), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n448), .A2(new_n451), .A3(new_n462), .A4(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n464), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT97), .ZN(new_n477));
  INV_X1    g291(.A(G217), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n188), .A2(new_n478), .A3(G953), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT97), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n464), .A2(new_n473), .A3(new_n481), .A4(new_n475), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n476), .A2(KEYINPUT97), .A3(new_n479), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n316), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(G478), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(G478), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n483), .A2(new_n316), .A3(new_n484), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n440), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n296), .A2(G952), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(G234), .B2(G237), .ZN(new_n492));
  AOI211_X1 g306(.A(new_n296), .B(new_n316), .C1(G234), .C2(G237), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n381), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n324), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n478), .B1(new_n316), .B2(G234), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n385), .A2(G125), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n327), .A2(G140), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n386), .B1(new_n501), .B2(new_n384), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n213), .ZN(new_n503));
  XNOR2_X1  g317(.A(KEYINPUT24), .B(G110), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT75), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G119), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(G128), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n508), .B1(new_n339), .B2(G128), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n503), .A2(new_n387), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(KEYINPUT66), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT66), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G119), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT23), .B1(new_n514), .B2(new_n209), .ZN(new_n515));
  OAI21_X1  g329(.A(KEYINPUT76), .B1(new_n339), .B2(G128), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT76), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n517), .A3(new_n209), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n508), .A2(KEYINPUT23), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G110), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n510), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g337(.A1(new_n506), .A2(new_n509), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n522), .A3(new_n520), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n387), .A2(new_n406), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n523), .B(KEYINPUT77), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT77), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n504), .A2(KEYINPUT75), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n509), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n388), .B2(new_n389), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n522), .B1(new_n519), .B2(new_n520), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n527), .B1(new_n524), .B2(new_n525), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT22), .B(G137), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n296), .A2(G221), .A3(G234), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n538), .B(new_n539), .Z(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n528), .A2(new_n537), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n529), .A3(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT25), .B1(new_n545), .B2(new_n316), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n547));
  INV_X1    g361(.A(new_n316), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n547), .B(new_n548), .C1(new_n542), .C2(new_n544), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n498), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n498), .A2(G902), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(KEYINPUT78), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n267), .A2(new_n219), .A3(new_n268), .ZN(new_n556));
  INV_X1    g370(.A(new_n260), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n256), .A2(G137), .ZN(new_n558));
  OAI21_X1  g372(.A(G131), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n264), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n236), .B2(new_n231), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n556), .A2(KEYINPUT30), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT30), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n207), .B1(new_n235), .B2(new_n209), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n282), .B2(new_n209), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n566), .A2(new_n210), .B1(new_n264), .B2(new_n262), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n564), .B1(new_n567), .B2(new_n561), .ZN(new_n568));
  INV_X1    g382(.A(new_n353), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n563), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n556), .A2(new_n353), .A3(new_n562), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT69), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT26), .B(G101), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n391), .A2(G210), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n571), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n572), .B1(new_n571), .B2(new_n578), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n555), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(KEYINPUT31), .A3(new_n570), .A4(new_n579), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n571), .A2(KEYINPUT28), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT28), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n556), .A2(new_n353), .A3(new_n562), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n569), .B1(new_n561), .B2(new_n567), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n577), .B(KEYINPUT70), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n582), .A2(new_n584), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(G472), .A2(G902), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n593), .B(KEYINPUT71), .Z(new_n594));
  OAI21_X1  g408(.A(KEYINPUT72), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT32), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n582), .A2(new_n584), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n590), .A2(new_n591), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n594), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n592), .A2(KEYINPUT32), .A3(new_n594), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(KEYINPUT72), .A3(new_n596), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n556), .A2(new_n562), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n569), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n588), .A2(KEYINPUT29), .A3(new_n608), .A4(new_n578), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT73), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n570), .A2(new_n571), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n577), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT29), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n612), .B(new_n613), .C1(new_n590), .C2(new_n591), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n316), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n554), .B1(new_n606), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n497), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  OAI21_X1  g433(.A(G472), .B1(new_n592), .B2(new_n548), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n604), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n554), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n324), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n363), .A2(new_n377), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n364), .ZN(new_n625));
  INV_X1    g439(.A(new_n325), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n365), .B1(new_n363), .B2(new_n377), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n430), .A2(new_n436), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n439), .A2(G475), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n495), .ZN(new_n632));
  INV_X1    g446(.A(G478), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n548), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n483), .A2(new_n484), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n476), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n479), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n476), .A2(new_n639), .A3(new_n480), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT33), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n635), .B1(new_n638), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n485), .A2(new_n633), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n631), .B(new_n632), .C1(new_n645), .C2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n623), .A2(new_n628), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  NAND2_X1  g466(.A1(new_n487), .A2(new_n489), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n440), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n495), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n623), .A2(new_n628), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  OR2_X1    g472(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n543), .B(new_n659), .Z(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n552), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n550), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n621), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n497), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT99), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT37), .B(G110), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  AOI21_X1  g481(.A(new_n662), .B1(new_n606), .B2(new_n616), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n492), .B1(new_n493), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n653), .A2(new_n440), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n653), .A2(new_n440), .A3(KEYINPUT100), .A4(new_n671), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n668), .A2(new_n324), .A3(new_n628), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  XOR2_X1   g492(.A(new_n670), .B(KEYINPUT39), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n324), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n681));
  INV_X1    g495(.A(G472), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n608), .A2(new_n571), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n591), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n580), .B2(new_n581), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n682), .B1(new_n685), .B2(new_n190), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n606), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n379), .A2(new_n380), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n440), .B1(new_n487), .B2(new_n489), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n325), .A3(new_n662), .ZN(new_n694));
  OR3_X1    g508(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n680), .A2(KEYINPUT40), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n681), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n211), .ZN(G45));
  AOI21_X1  g512(.A(KEYINPUT33), .B1(new_n483), .B2(new_n484), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n637), .B1(new_n641), .B2(new_n642), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n634), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n701), .A2(new_n646), .B1(new_n629), .B2(new_n630), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n671), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n668), .A2(new_n324), .A3(new_n628), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  AND3_X1   g520(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n708), .A3(new_n191), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n617), .A3(new_n628), .A4(new_n649), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n617), .A3(new_n628), .A4(new_n655), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NOR2_X1   g528(.A1(new_n490), .A2(new_n495), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n709), .A2(new_n715), .A3(new_n628), .A4(new_n668), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G119), .ZN(G21));
  AND2_X1   g531(.A1(new_n628), .A2(new_n693), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n632), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n588), .A2(new_n608), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n591), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n597), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n600), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n620), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n554), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n720), .A2(new_n709), .A3(KEYINPUT102), .A4(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT102), .ZN(new_n728));
  INV_X1    g542(.A(new_n708), .ZN(new_n729));
  INV_X1    g543(.A(new_n191), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n317), .A4(new_n726), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n728), .B1(new_n731), .B2(new_n719), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NOR2_X1   g548(.A1(new_n707), .A2(new_n708), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n736), .B1(new_n662), .B2(new_n725), .ZN(new_n737));
  INV_X1    g551(.A(new_n552), .ZN(new_n738));
  INV_X1    g552(.A(new_n660), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n550), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n620), .A3(KEYINPUT103), .A4(new_n724), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n703), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n735), .A2(new_n730), .A3(new_n628), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  NAND2_X1  g558(.A1(new_n317), .A2(new_n323), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n191), .A2(new_n626), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n690), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT104), .B1(new_n601), .B2(new_n602), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n599), .A2(new_n596), .A3(new_n600), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT32), .B1(new_n592), .B2(new_n594), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n616), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n554), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n704), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT42), .B1(new_n749), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n747), .B1(new_n317), .B2(new_n323), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n617), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n758), .B2(new_n762), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G131), .ZN(G33));
  NAND2_X1  g580(.A1(new_n674), .A2(new_n675), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n617), .A2(new_n760), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G134), .ZN(G36));
  AND2_X1   g586(.A1(new_n314), .A2(new_n316), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n307), .B1(new_n303), .B2(new_n304), .ZN(new_n774));
  INV_X1    g588(.A(new_n321), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(KEYINPUT45), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT107), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n778), .A3(KEYINPUT45), .A4(new_n775), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n780), .B1(new_n320), .B2(new_n321), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n777), .A2(G469), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT46), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n318), .A2(new_n783), .ZN(new_n784));
  AOI22_X1  g598(.A1(new_n773), .A2(new_n315), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n318), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n730), .A3(new_n679), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n792));
  AND2_X1   g606(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n793));
  OAI221_X1 g607(.A(new_n440), .B1(new_n792), .B2(new_n793), .C1(new_n645), .C2(new_n647), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n631), .B1(new_n646), .B2(new_n701), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n794), .B1(new_n795), .B2(new_n793), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n740), .A2(new_n621), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n796), .A2(KEYINPUT44), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n690), .A2(new_n325), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT44), .B1(new_n796), .B2(new_n797), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n791), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NAND2_X1  g618(.A1(new_n782), .A2(new_n784), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n317), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT46), .B1(new_n782), .B2(new_n786), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n730), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT47), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI211_X1 g624(.A(KEYINPUT47), .B(new_n730), .C1(new_n806), .C2(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n606), .A2(new_n616), .ZN(new_n813));
  NOR4_X1   g627(.A1(new_n813), .A2(new_n756), .A3(new_n800), .A4(new_n703), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n692), .A2(new_n796), .A3(new_n626), .A4(new_n492), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n818), .A2(new_n731), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n818), .B2(new_n731), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n800), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n709), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n796), .A2(new_n492), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n737), .A2(new_n741), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n689), .A2(new_n756), .A3(new_n492), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n631), .A2(new_n645), .A3(new_n647), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n822), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT47), .B1(new_n789), .B2(new_n730), .ZN(new_n834));
  INV_X1    g648(.A(new_n811), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT112), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n810), .A2(new_n837), .A3(new_n811), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT109), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n707), .B2(new_n708), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n839), .A2(new_n841), .A3(new_n191), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n796), .A2(new_n492), .A3(new_n726), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n800), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n833), .B1(new_n847), .B2(KEYINPUT113), .ZN(new_n848));
  INV_X1    g662(.A(new_n846), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n842), .B1(new_n812), .B2(KEYINPUT112), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n850), .B2(new_n838), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT51), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT114), .B1(new_n828), .B2(new_n832), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n822), .A2(KEYINPUT51), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n843), .A2(new_n810), .A3(new_n811), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n846), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n828), .A2(new_n832), .A3(KEYINPUT114), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n856), .A2(new_n858), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n709), .A2(new_n628), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT115), .B1(new_n863), .B2(new_n845), .ZN(new_n864));
  INV_X1    g678(.A(new_n845), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n628), .A4(new_n709), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n491), .B1(new_n830), .B2(new_n702), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT48), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n755), .A2(new_n756), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n870), .B1(new_n826), .B2(new_n872), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n824), .A2(KEYINPUT48), .A3(new_n871), .A4(new_n825), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n868), .B(new_n869), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n875), .A2(new_n876), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n862), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n817), .B1(new_n854), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  INV_X1    g696(.A(new_n833), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n851), .B2(new_n852), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n847), .A2(KEYINPUT113), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n875), .A2(new_n876), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n857), .B1(new_n846), .B2(new_n859), .ZN(new_n888));
  INV_X1    g702(.A(new_n861), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n855), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n887), .A2(new_n877), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n891), .A3(KEYINPUT117), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n743), .A2(new_n677), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT52), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n740), .A2(new_n191), .A3(new_n670), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n688), .A2(new_n745), .A3(new_n718), .A4(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n894), .A2(new_n895), .A3(new_n705), .A4(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n743), .A2(new_n677), .A3(new_n705), .A4(new_n897), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT52), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n490), .A2(new_n670), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n668), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n742), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n760), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n905), .A2(new_n771), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n765), .A2(new_n898), .A3(new_n900), .A4(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n710), .A2(new_n713), .A3(new_n716), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n496), .B(new_n324), .C1(new_n617), .C2(new_n663), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT110), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n648), .B2(new_n381), .ZN(new_n911));
  INV_X1    g725(.A(new_n366), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n624), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n626), .B1(new_n913), .B2(new_n378), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n632), .A3(new_n653), .A4(new_n440), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(KEYINPUT110), .A3(new_n702), .A4(new_n632), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n911), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(new_n324), .A3(new_n622), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT111), .B1(new_n909), .B2(new_n918), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n909), .A2(new_n918), .A3(KEYINPUT111), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n908), .B(new_n733), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n893), .B1(new_n907), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT54), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n733), .A2(new_n710), .A3(new_n713), .A4(new_n716), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n920), .A2(new_n919), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n899), .B(new_n895), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n894), .A2(new_n895), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n905), .A2(new_n771), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n758), .A2(KEYINPUT53), .A3(new_n762), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n922), .A2(new_n923), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n928), .A2(new_n893), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n929), .A2(new_n763), .A3(new_n764), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n926), .A2(new_n934), .A3(new_n927), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n923), .B1(new_n922), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n881), .A2(new_n892), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g753(.A1(G952), .A2(G953), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n839), .A2(new_n841), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n943), .A2(KEYINPUT49), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(KEYINPUT49), .ZN(new_n945));
  AND4_X1   g759(.A1(new_n756), .A2(new_n692), .A3(new_n746), .A4(new_n795), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n689), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n947), .ZN(G75));
  NAND2_X1  g762(.A1(new_n922), .A2(new_n932), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n548), .A3(new_n365), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n360), .A2(new_n362), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(new_n336), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT55), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n955), .B1(new_n950), .B2(new_n951), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n296), .A2(G952), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(G51));
  INV_X1    g773(.A(new_n782), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n949), .A2(new_n548), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT118), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n923), .B1(new_n922), .B2(new_n932), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n933), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n318), .B(KEYINPUT57), .Z(new_n966));
  OAI21_X1  g780(.A(new_n314), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n958), .B1(new_n963), .B2(new_n967), .ZN(G54));
  NAND2_X1  g782(.A1(new_n949), .A2(new_n548), .ZN(new_n969));
  NAND2_X1  g783(.A1(KEYINPUT58), .A2(G475), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n427), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n958), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n969), .A2(new_n427), .A3(new_n970), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(G60));
  NAND2_X1  g789(.A1(new_n638), .A2(new_n644), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n933), .A2(new_n937), .ZN(new_n977));
  NAND2_X1  g791(.A1(G478), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT59), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n976), .A2(new_n979), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n972), .B1(new_n965), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n980), .A2(new_n982), .ZN(G63));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT120), .ZN(new_n985));
  XNOR2_X1  g799(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n949), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n545), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(KEYINPUT121), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n949), .A2(new_n660), .A3(new_n987), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n992), .A2(new_n972), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n545), .B1(new_n949), .B2(new_n987), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT121), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n991), .A2(new_n993), .A3(KEYINPUT61), .A4(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT61), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n992), .A2(new_n972), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n994), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(G66));
  OAI21_X1  g815(.A(G953), .B1(new_n494), .B2(new_n334), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1002), .B1(new_n926), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n952), .B1(G898), .B2(new_n296), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G69));
  INV_X1    g819(.A(KEYINPUT124), .ZN(new_n1006));
  INV_X1    g820(.A(new_n702), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n800), .B1(new_n1007), .B2(new_n654), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n617), .A2(new_n324), .A3(new_n1008), .A4(new_n679), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n815), .A2(new_n803), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n743), .A2(new_n677), .A3(new_n705), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT123), .ZN(new_n1012));
  INV_X1    g826(.A(new_n697), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1010), .B1(new_n1014), .B2(KEYINPUT62), .ZN(new_n1015));
  OR2_X1    g829(.A1(new_n1011), .A2(KEYINPUT123), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1011), .A2(KEYINPUT123), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n697), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT62), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(G953), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n563), .A2(new_n568), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT122), .Z(new_n1023));
  OAI21_X1  g837(.A(new_n420), .B1(new_n407), .B2(new_n419), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1006), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1025), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n815), .A2(new_n803), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1028), .B(new_n1009), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g845(.A(KEYINPUT124), .B(new_n1027), .C1(new_n1031), .C2(G953), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1027), .B1(G900), .B2(G953), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n872), .A2(new_n718), .ZN(new_n1034));
  AOI22_X1  g848(.A1(new_n791), .A2(new_n1034), .B1(new_n770), .B2(new_n769), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1028), .A2(new_n1035), .A3(new_n765), .A4(new_n1012), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1033), .B1(new_n1036), .B2(G953), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1026), .A2(new_n1032), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n296), .B1(G227), .B2(G900), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1039), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1026), .A2(new_n1032), .A3(new_n1041), .A4(new_n1037), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1040), .A2(new_n1042), .ZN(G72));
  XNOR2_X1  g857(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n682), .A2(new_n190), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1044), .B(new_n1045), .Z(new_n1046));
  INV_X1    g860(.A(new_n1046), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1047), .B1(new_n1036), .B2(new_n921), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n611), .A2(new_n578), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n958), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AND2_X1   g864(.A1(new_n922), .A2(new_n936), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT127), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n612), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1053), .B1(new_n581), .B2(new_n580), .ZN(new_n1054));
  NOR2_X1   g868(.A1(new_n612), .A2(new_n1052), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1047), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1050), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g871(.A1(new_n1029), .A2(new_n1030), .A3(new_n921), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1058), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n1059), .A2(KEYINPUT126), .A3(new_n1047), .ZN(new_n1060));
  INV_X1    g874(.A(KEYINPUT126), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1061), .B1(new_n1058), .B2(new_n1046), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n577), .B1(new_n570), .B2(new_n571), .ZN(new_n1064));
  AOI21_X1  g878(.A(new_n1057), .B1(new_n1063), .B2(new_n1064), .ZN(G57));
endmodule


