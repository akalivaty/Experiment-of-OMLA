

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778;

  INV_X1 U377 ( .A(G953), .ZN(n769) );
  AND2_X2 U378 ( .A1(n409), .A2(n368), .ZN(n641) );
  OR2_X2 U379 ( .A1(n659), .A2(G902), .ZN(n537) );
  NOR2_X1 U380 ( .A1(n697), .A2(n575), .ZN(n597) );
  XNOR2_X2 U381 ( .A(n408), .B(n462), .ZN(n652) );
  INV_X1 U382 ( .A(KEYINPUT81), .ZN(n449) );
  XNOR2_X1 U383 ( .A(n372), .B(KEYINPUT84), .ZN(n644) );
  NOR2_X1 U384 ( .A1(n609), .A2(n370), .ZN(n369) );
  XNOR2_X1 U385 ( .A(n618), .B(KEYINPUT35), .ZN(n776) );
  XNOR2_X1 U386 ( .A(n631), .B(n395), .ZN(n680) );
  NAND2_X1 U387 ( .A1(n406), .A2(n405), .ZN(n512) );
  XNOR2_X1 U388 ( .A(n478), .B(KEYINPUT0), .ZN(n611) );
  NAND2_X1 U389 ( .A1(n417), .A2(n413), .ZN(n478) );
  AND2_X1 U390 ( .A1(n686), .A2(n699), .ZN(n405) );
  XNOR2_X1 U391 ( .A(n535), .B(n357), .ZN(n751) );
  XNOR2_X1 U392 ( .A(n489), .B(n424), .ZN(n766) );
  XNOR2_X1 U393 ( .A(n450), .B(n449), .ZN(n479) );
  XNOR2_X1 U394 ( .A(n425), .B(G125), .ZN(n489) );
  XNOR2_X1 U395 ( .A(G143), .B(G128), .ZN(n450) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n530) );
  OR2_X1 U397 ( .A1(n386), .A2(n382), .ZN(n381) );
  XNOR2_X1 U398 ( .A(n446), .B(KEYINPUT85), .ZN(n639) );
  NAND2_X1 U399 ( .A1(n448), .A2(n447), .ZN(n446) );
  INV_X1 U400 ( .A(n619), .ZN(n447) );
  XNOR2_X1 U401 ( .A(n393), .B(G101), .ZN(n529) );
  XNOR2_X1 U402 ( .A(n528), .B(n527), .ZN(n539) );
  XNOR2_X1 U403 ( .A(G131), .B(G134), .ZN(n527) );
  XNOR2_X1 U404 ( .A(n392), .B(n451), .ZN(n535) );
  XNOR2_X1 U405 ( .A(G119), .B(G116), .ZN(n451) );
  XNOR2_X1 U406 ( .A(n452), .B(KEYINPUT3), .ZN(n392) );
  XNOR2_X1 U407 ( .A(G113), .B(KEYINPUT69), .ZN(n452) );
  INV_X1 U408 ( .A(G146), .ZN(n425) );
  XNOR2_X1 U409 ( .A(n479), .B(KEYINPUT4), .ZN(n528) );
  NOR2_X1 U410 ( .A1(n697), .A2(n696), .ZN(n625) );
  NOR2_X1 U411 ( .A1(n627), .A2(n439), .ZN(n430) );
  XNOR2_X1 U412 ( .A(n621), .B(KEYINPUT1), .ZN(n696) );
  XNOR2_X1 U413 ( .A(G110), .B(KEYINPUT88), .ZN(n454) );
  INV_X1 U414 ( .A(KEYINPUT73), .ZN(n382) );
  NOR2_X1 U415 ( .A1(n593), .A2(KEYINPUT47), .ZN(n387) );
  NOR2_X1 U416 ( .A1(n776), .A2(n411), .ZN(n410) );
  INV_X1 U417 ( .A(KEYINPUT44), .ZN(n411) );
  AND2_X1 U418 ( .A1(n639), .A2(n421), .ZN(n420) );
  NAND2_X1 U419 ( .A1(KEYINPUT64), .A2(KEYINPUT44), .ZN(n421) );
  NAND2_X1 U420 ( .A1(n680), .A2(n669), .ZN(n632) );
  NAND2_X1 U421 ( .A1(n645), .A2(n469), .ZN(n444) );
  XNOR2_X1 U422 ( .A(n489), .B(n458), .ZN(n459) );
  XNOR2_X1 U423 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n458) );
  INV_X1 U424 ( .A(n684), .ZN(n608) );
  XNOR2_X1 U425 ( .A(n396), .B(n604), .ZN(n371) );
  AND2_X1 U426 ( .A1(n603), .A2(n602), .ZN(n427) );
  XNOR2_X1 U427 ( .A(n577), .B(n576), .ZN(n691) );
  NOR2_X1 U428 ( .A1(n627), .A2(n626), .ZN(n708) );
  NAND2_X1 U429 ( .A1(n362), .A2(n441), .ZN(n577) );
  NAND2_X1 U430 ( .A1(n652), .A2(n469), .ZN(n445) );
  INV_X1 U431 ( .A(n652), .ZN(n443) );
  NAND2_X1 U432 ( .A1(n443), .A2(n442), .ZN(n441) );
  XNOR2_X1 U433 ( .A(n501), .B(n500), .ZN(n594) );
  OR2_X1 U434 ( .A1(n736), .A2(G902), .ZN(n501) );
  AND2_X1 U435 ( .A1(n414), .A2(n415), .ZN(n413) );
  INV_X1 U436 ( .A(n431), .ZN(n415) );
  XNOR2_X1 U437 ( .A(n389), .B(n391), .ZN(n403) );
  XNOR2_X1 U438 ( .A(n390), .B(n534), .ZN(n389) );
  XNOR2_X1 U439 ( .A(KEYINPUT16), .B(G122), .ZN(n453) );
  XNOR2_X1 U440 ( .A(n518), .B(n517), .ZN(n520) );
  XNOR2_X1 U441 ( .A(n538), .B(G110), .ZN(n518) );
  XNOR2_X1 U442 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n516) );
  XNOR2_X1 U443 ( .A(G107), .B(G122), .ZN(n480) );
  INV_X1 U444 ( .A(KEYINPUT11), .ZN(n400) );
  XNOR2_X1 U445 ( .A(G113), .B(G104), .ZN(n490) );
  XOR2_X1 U446 ( .A(KEYINPUT101), .B(G122), .Z(n491) );
  XOR2_X1 U447 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n494) );
  XNOR2_X1 U448 ( .A(G140), .B(KEYINPUT10), .ZN(n424) );
  XNOR2_X1 U449 ( .A(n765), .B(n544), .ZN(n731) );
  NAND2_X1 U450 ( .A1(n722), .A2(n645), .ZN(n649) );
  XNOR2_X1 U451 ( .A(n610), .B(KEYINPUT33), .ZN(n725) );
  NAND2_X1 U452 ( .A1(n429), .A2(n404), .ZN(n575) );
  NOR2_X1 U453 ( .A1(n621), .A2(n574), .ZN(n404) );
  XNOR2_X1 U454 ( .A(n430), .B(n366), .ZN(n429) );
  XNOR2_X1 U455 ( .A(n524), .B(n358), .ZN(n422) );
  BUF_X1 U456 ( .A(n735), .Z(n744) );
  AND2_X1 U457 ( .A1(n655), .A2(G953), .ZN(n748) );
  NAND2_X1 U458 ( .A1(n364), .A2(n378), .ZN(n603) );
  INV_X1 U459 ( .A(G237), .ZN(n465) );
  XNOR2_X1 U460 ( .A(n394), .B(n529), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n531), .B(G146), .ZN(n394) );
  XNOR2_X1 U462 ( .A(KEYINPUT74), .B(KEYINPUT97), .ZN(n532) );
  XOR2_X1 U463 ( .A(G137), .B(KEYINPUT5), .Z(n533) );
  XOR2_X1 U464 ( .A(G137), .B(KEYINPUT67), .Z(n538) );
  XOR2_X1 U465 ( .A(G146), .B(G140), .Z(n541) );
  XNOR2_X1 U466 ( .A(n539), .B(n538), .ZN(n765) );
  NAND2_X1 U467 ( .A1(n435), .A2(n434), .ZN(n433) );
  INV_X1 U468 ( .A(n444), .ZN(n435) );
  NAND2_X1 U469 ( .A1(n706), .A2(n373), .ZN(n376) );
  XNOR2_X1 U470 ( .A(n528), .B(n751), .ZN(n408) );
  AND2_X2 U471 ( .A1(n371), .A2(n426), .ZN(n767) );
  NOR2_X1 U472 ( .A1(n694), .A2(n581), .ZN(n583) );
  XNOR2_X1 U473 ( .A(n679), .B(n397), .ZN(n606) );
  INV_X1 U474 ( .A(KEYINPUT105), .ZN(n397) );
  NOR2_X1 U475 ( .A1(n445), .A2(n440), .ZN(n437) );
  NAND2_X1 U476 ( .A1(n436), .A2(n432), .ZN(n431) );
  AND2_X1 U477 ( .A1(n433), .A2(n438), .ZN(n432) );
  NAND2_X1 U478 ( .A1(n443), .A2(n360), .ZN(n436) );
  NAND2_X1 U479 ( .A1(n439), .A2(n471), .ZN(n438) );
  NAND2_X1 U480 ( .A1(n354), .A2(n362), .ZN(n417) );
  AND2_X1 U481 ( .A1(n375), .A2(n374), .ZN(n589) );
  INV_X1 U482 ( .A(n621), .ZN(n374) );
  XNOR2_X1 U483 ( .A(n376), .B(n585), .ZN(n375) );
  XOR2_X1 U484 ( .A(KEYINPUT112), .B(KEYINPUT28), .Z(n585) );
  XNOR2_X1 U485 ( .A(n594), .B(n398), .ZN(n591) );
  INV_X1 U486 ( .A(KEYINPUT103), .ZN(n398) );
  XNOR2_X1 U487 ( .A(n572), .B(n571), .ZN(n697) );
  AND2_X1 U488 ( .A1(n700), .A2(n699), .ZN(n572) );
  BUF_X1 U489 ( .A(n696), .Z(n402) );
  XNOR2_X1 U490 ( .A(G128), .B(G119), .ZN(n519) );
  XNOR2_X1 U491 ( .A(n483), .B(n407), .ZN(n487) );
  XNOR2_X1 U492 ( .A(n484), .B(n363), .ZN(n407) );
  XNOR2_X1 U493 ( .A(n495), .B(n399), .ZN(n497) );
  XNOR2_X1 U494 ( .A(n496), .B(n400), .ZN(n399) );
  NAND2_X1 U495 ( .A1(n636), .A2(n568), .ZN(n570) );
  INV_X1 U496 ( .A(KEYINPUT98), .ZN(n395) );
  XNOR2_X1 U497 ( .A(n630), .B(n629), .ZN(n631) );
  XOR2_X1 U498 ( .A(n592), .B(KEYINPUT107), .Z(n677) );
  XNOR2_X1 U499 ( .A(n401), .B(n367), .ZN(n734) );
  NAND2_X1 U500 ( .A1(n744), .A2(G469), .ZN(n401) );
  AND2_X1 U501 ( .A1(n441), .A2(n471), .ZN(n354) );
  AND2_X1 U502 ( .A1(n383), .A2(n365), .ZN(n355) );
  OR2_X1 U503 ( .A1(n716), .A2(n477), .ZN(n356) );
  XOR2_X1 U504 ( .A(n453), .B(KEYINPUT72), .Z(n357) );
  XOR2_X1 U505 ( .A(n526), .B(n525), .Z(n358) );
  XOR2_X1 U506 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n359) );
  NAND2_X1 U507 ( .A1(n687), .A2(KEYINPUT19), .ZN(n440) );
  INV_X1 U508 ( .A(n440), .ZN(n434) );
  XNOR2_X1 U509 ( .A(n579), .B(n578), .ZN(n605) );
  AND2_X1 U510 ( .A1(n442), .A2(n434), .ZN(n360) );
  INV_X1 U511 ( .A(n505), .ZN(n645) );
  AND2_X1 U512 ( .A1(n416), .A2(n417), .ZN(n361) );
  AND2_X1 U513 ( .A1(n445), .A2(n444), .ZN(n362) );
  INV_X1 U514 ( .A(n609), .ZN(n426) );
  NAND2_X1 U515 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U516 ( .A(G134), .B(G116), .Z(n363) );
  AND2_X1 U517 ( .A1(n381), .A2(n379), .ZN(n364) );
  AND2_X1 U518 ( .A1(n384), .A2(n382), .ZN(n365) );
  XOR2_X1 U519 ( .A(n573), .B(KEYINPUT110), .Z(n366) );
  XOR2_X1 U520 ( .A(n733), .B(n732), .Z(n367) );
  OR2_X1 U521 ( .A1(n640), .A2(KEYINPUT44), .ZN(n368) );
  INV_X1 U522 ( .A(KEYINPUT2), .ZN(n370) );
  NAND2_X1 U523 ( .A1(n371), .A2(n369), .ZN(n372) );
  NOR2_X1 U524 ( .A1(n700), .A2(n377), .ZN(n373) );
  INV_X1 U525 ( .A(n584), .ZN(n377) );
  NAND2_X1 U526 ( .A1(n386), .A2(n355), .ZN(n378) );
  NAND2_X1 U527 ( .A1(n380), .A2(KEYINPUT73), .ZN(n379) );
  NAND2_X1 U528 ( .A1(n383), .A2(n384), .ZN(n380) );
  NAND2_X1 U529 ( .A1(n675), .A2(KEYINPUT47), .ZN(n383) );
  AND2_X1 U530 ( .A1(n385), .A2(n674), .ZN(n384) );
  NAND2_X1 U531 ( .A1(n593), .A2(KEYINPUT47), .ZN(n385) );
  NAND2_X1 U532 ( .A1(n388), .A2(n387), .ZN(n386) );
  INV_X1 U533 ( .A(n675), .ZN(n388) );
  INV_X1 U534 ( .A(n535), .ZN(n391) );
  INV_X1 U535 ( .A(KEYINPUT65), .ZN(n393) );
  OR2_X1 U536 ( .A1(n639), .A2(n640), .ZN(n412) );
  OR2_X2 U537 ( .A1(n746), .A2(G902), .ZN(n423) );
  AND2_X1 U538 ( .A1(n513), .A2(G221), .ZN(n514) );
  NOR2_X1 U539 ( .A1(n605), .A2(n592), .ZN(n580) );
  NAND2_X1 U540 ( .A1(n427), .A2(n428), .ZN(n396) );
  NAND2_X1 U541 ( .A1(n606), .A2(n592), .ZN(n688) );
  XNOR2_X2 U542 ( .A(n570), .B(n569), .ZN(n620) );
  NOR2_X1 U543 ( .A1(n437), .A2(n356), .ZN(n414) );
  NAND2_X1 U544 ( .A1(n725), .A2(n628), .ZN(n614) );
  NOR2_X1 U545 ( .A1(n662), .A2(n748), .ZN(n663) );
  XNOR2_X1 U546 ( .A(n403), .B(n539), .ZN(n659) );
  INV_X1 U547 ( .A(n611), .ZN(n406) );
  NAND2_X1 U548 ( .A1(n412), .A2(n410), .ZN(n409) );
  NOR2_X1 U549 ( .A1(n437), .A2(n431), .ZN(n416) );
  NAND2_X1 U550 ( .A1(n638), .A2(n418), .ZN(n642) );
  NAND2_X1 U551 ( .A1(n419), .A2(n420), .ZN(n418) );
  NAND2_X1 U552 ( .A1(n776), .A2(KEYINPUT64), .ZN(n419) );
  XNOR2_X2 U553 ( .A(n423), .B(n422), .ZN(n700) );
  XNOR2_X1 U554 ( .A(n588), .B(KEYINPUT46), .ZN(n428) );
  INV_X1 U555 ( .A(n627), .ZN(n706) );
  INV_X1 U556 ( .A(n687), .ZN(n439) );
  NOR2_X1 U557 ( .A1(n645), .A2(n469), .ZN(n442) );
  INV_X1 U558 ( .A(n620), .ZN(n448) );
  XNOR2_X2 U559 ( .A(n590), .B(KEYINPUT80), .ZN(n675) );
  XNOR2_X1 U560 ( .A(n522), .B(n521), .ZN(n746) );
  XNOR2_X1 U561 ( .A(n515), .B(n514), .ZN(n522) );
  XNOR2_X1 U562 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U563 ( .A(KEYINPUT48), .ZN(n604) );
  INV_X1 U564 ( .A(KEYINPUT78), .ZN(n612) );
  XNOR2_X1 U565 ( .A(n612), .B(KEYINPUT34), .ZN(n613) );
  XNOR2_X1 U566 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U567 ( .A(n614), .B(n613), .ZN(n617) );
  XOR2_X1 U568 ( .A(G104), .B(G107), .Z(n455) );
  XNOR2_X1 U569 ( .A(n455), .B(n454), .ZN(n753) );
  INV_X1 U570 ( .A(n529), .ZN(n456) );
  XNOR2_X1 U571 ( .A(n753), .B(n456), .ZN(n543) );
  NAND2_X1 U572 ( .A1(n769), .A2(G224), .ZN(n457) );
  XNOR2_X1 U573 ( .A(n457), .B(KEYINPUT89), .ZN(n460) );
  XNOR2_X1 U574 ( .A(n543), .B(n461), .ZN(n462) );
  XNOR2_X1 U575 ( .A(G902), .B(KEYINPUT87), .ZN(n464) );
  INV_X1 U576 ( .A(KEYINPUT15), .ZN(n463) );
  XNOR2_X1 U577 ( .A(n464), .B(n463), .ZN(n505) );
  INV_X1 U578 ( .A(G902), .ZN(n466) );
  NAND2_X1 U579 ( .A1(n466), .A2(n465), .ZN(n470) );
  NAND2_X1 U580 ( .A1(n470), .A2(G210), .ZN(n468) );
  INV_X1 U581 ( .A(KEYINPUT82), .ZN(n467) );
  XNOR2_X1 U582 ( .A(n468), .B(n467), .ZN(n469) );
  NAND2_X1 U583 ( .A1(n470), .A2(G214), .ZN(n687) );
  INV_X1 U584 ( .A(KEYINPUT19), .ZN(n471) );
  NAND2_X1 U585 ( .A1(G237), .A2(G234), .ZN(n473) );
  INV_X1 U586 ( .A(KEYINPUT14), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n473), .B(n472), .ZN(n716) );
  NAND2_X1 U588 ( .A1(n769), .A2(G952), .ZN(n553) );
  INV_X1 U589 ( .A(G898), .ZN(n475) );
  NAND2_X1 U590 ( .A1(G953), .A2(G902), .ZN(n550) );
  INV_X1 U591 ( .A(n550), .ZN(n474) );
  NAND2_X1 U592 ( .A1(n475), .A2(n474), .ZN(n476) );
  AND2_X1 U593 ( .A1(n553), .A2(n476), .ZN(n477) );
  INV_X1 U594 ( .A(n479), .ZN(n484) );
  XOR2_X1 U595 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n481) );
  XNOR2_X1 U596 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U597 ( .A(n482), .B(KEYINPUT104), .Z(n483) );
  NAND2_X1 U598 ( .A1(G234), .A2(n769), .ZN(n485) );
  XOR2_X1 U599 ( .A(KEYINPUT8), .B(n485), .Z(n513) );
  NAND2_X1 U600 ( .A1(G217), .A2(n513), .ZN(n486) );
  XNOR2_X1 U601 ( .A(n487), .B(n486), .ZN(n741) );
  NOR2_X1 U602 ( .A1(n741), .A2(G902), .ZN(n488) );
  XNOR2_X1 U603 ( .A(n488), .B(G478), .ZN(n549) );
  XNOR2_X1 U604 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n766), .B(n492), .ZN(n498) );
  NAND2_X1 U606 ( .A1(G214), .A2(n530), .ZN(n493) );
  XNOR2_X1 U607 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U608 ( .A(G143), .B(G131), .ZN(n496) );
  XNOR2_X1 U609 ( .A(n498), .B(n497), .ZN(n736) );
  XOR2_X1 U610 ( .A(G475), .B(KEYINPUT102), .Z(n499) );
  XNOR2_X1 U611 ( .A(KEYINPUT13), .B(n499), .ZN(n500) );
  INV_X1 U612 ( .A(n594), .ZN(n502) );
  NAND2_X1 U613 ( .A1(n549), .A2(n502), .ZN(n504) );
  INV_X1 U614 ( .A(KEYINPUT106), .ZN(n503) );
  XNOR2_X1 U615 ( .A(n504), .B(n503), .ZN(n686) );
  NAND2_X1 U616 ( .A1(n505), .A2(G234), .ZN(n507) );
  XNOR2_X1 U617 ( .A(KEYINPUT20), .B(KEYINPUT94), .ZN(n506) );
  XNOR2_X1 U618 ( .A(n507), .B(n506), .ZN(n523) );
  AND2_X1 U619 ( .A1(n523), .A2(G221), .ZN(n510) );
  INV_X1 U620 ( .A(KEYINPUT95), .ZN(n508) );
  XNOR2_X1 U621 ( .A(n508), .B(KEYINPUT21), .ZN(n509) );
  XNOR2_X1 U622 ( .A(n510), .B(n509), .ZN(n699) );
  XNOR2_X1 U623 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n511) );
  XNOR2_X2 U624 ( .A(n512), .B(n511), .ZN(n636) );
  XNOR2_X1 U625 ( .A(KEYINPUT23), .B(n766), .ZN(n515) );
  XNOR2_X1 U626 ( .A(n359), .B(n516), .ZN(n517) );
  NAND2_X1 U627 ( .A1(G217), .A2(n523), .ZN(n524) );
  XNOR2_X1 U628 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n526) );
  INV_X1 U629 ( .A(KEYINPUT76), .ZN(n525) );
  NAND2_X1 U630 ( .A1(n530), .A2(G210), .ZN(n531) );
  XNOR2_X1 U631 ( .A(n533), .B(n532), .ZN(n534) );
  INV_X1 U632 ( .A(G472), .ZN(n536) );
  XNOR2_X2 U633 ( .A(n537), .B(n536), .ZN(n627) );
  NOR2_X1 U634 ( .A1(n700), .A2(n706), .ZN(n547) );
  NAND2_X1 U635 ( .A1(G227), .A2(n769), .ZN(n540) );
  XNOR2_X1 U636 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n543), .B(n542), .ZN(n544) );
  NOR2_X1 U638 ( .A1(G902), .A2(n731), .ZN(n546) );
  XNOR2_X1 U639 ( .A(KEYINPUT68), .B(G469), .ZN(n545) );
  XNOR2_X2 U640 ( .A(n546), .B(n545), .ZN(n621) );
  AND2_X1 U641 ( .A1(n547), .A2(n402), .ZN(n548) );
  AND2_X1 U642 ( .A1(n636), .A2(n548), .ZN(n619) );
  XOR2_X1 U643 ( .A(G110), .B(n619), .Z(G12) );
  INV_X1 U644 ( .A(n402), .ZN(n562) );
  NAND2_X1 U645 ( .A1(n549), .A2(n591), .ZN(n592) );
  INV_X1 U646 ( .A(n699), .ZN(n557) );
  NOR2_X1 U647 ( .A1(n550), .A2(n716), .ZN(n551) );
  XOR2_X1 U648 ( .A(KEYINPUT108), .B(n551), .Z(n552) );
  NOR2_X1 U649 ( .A1(G900), .A2(n552), .ZN(n555) );
  NOR2_X1 U650 ( .A1(n716), .A2(n553), .ZN(n554) );
  NOR2_X1 U651 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U652 ( .A(KEYINPUT83), .B(n556), .Z(n574) );
  NOR2_X1 U653 ( .A1(n557), .A2(n574), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n584), .A2(n687), .ZN(n558) );
  NOR2_X1 U655 ( .A1(n677), .A2(n558), .ZN(n561) );
  XNOR2_X1 U656 ( .A(n627), .B(KEYINPUT6), .ZN(n633) );
  INV_X1 U657 ( .A(n633), .ZN(n559) );
  NOR2_X1 U658 ( .A1(n700), .A2(n559), .ZN(n560) );
  NAND2_X1 U659 ( .A1(n561), .A2(n560), .ZN(n599) );
  NOR2_X1 U660 ( .A1(n562), .A2(n599), .ZN(n564) );
  XNOR2_X1 U661 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n563) );
  XNOR2_X1 U662 ( .A(n564), .B(n563), .ZN(n565) );
  INV_X1 U663 ( .A(n577), .ZN(n598) );
  NAND2_X1 U664 ( .A1(n565), .A2(n598), .ZN(n607) );
  XNOR2_X1 U665 ( .A(n607), .B(G140), .ZN(G42) );
  NOR2_X1 U666 ( .A1(n696), .A2(n700), .ZN(n567) );
  XNOR2_X1 U667 ( .A(n633), .B(KEYINPUT79), .ZN(n566) );
  AND2_X1 U668 ( .A1(n567), .A2(n566), .ZN(n568) );
  INV_X1 U669 ( .A(KEYINPUT32), .ZN(n569) );
  XOR2_X1 U670 ( .A(n620), .B(G119), .Z(G21) );
  INV_X1 U671 ( .A(KEYINPUT66), .ZN(n571) );
  XNOR2_X1 U672 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n573) );
  INV_X1 U673 ( .A(KEYINPUT38), .ZN(n576) );
  NAND2_X1 U674 ( .A1(n597), .A2(n691), .ZN(n579) );
  XOR2_X1 U675 ( .A(KEYINPUT70), .B(KEYINPUT39), .Z(n578) );
  XNOR2_X1 U676 ( .A(n580), .B(KEYINPUT40), .ZN(n778) );
  XOR2_X1 U677 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n587) );
  NAND2_X1 U678 ( .A1(n686), .A2(n687), .ZN(n694) );
  INV_X1 U679 ( .A(n691), .ZN(n581) );
  XNOR2_X1 U680 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n582) );
  XNOR2_X1 U681 ( .A(n583), .B(n582), .ZN(n724) );
  NAND2_X1 U682 ( .A1(n724), .A2(n589), .ZN(n586) );
  XNOR2_X1 U683 ( .A(n587), .B(n586), .ZN(n777) );
  NOR2_X1 U684 ( .A1(n778), .A2(n777), .ZN(n588) );
  NAND2_X1 U685 ( .A1(n589), .A2(n361), .ZN(n590) );
  OR2_X1 U686 ( .A1(n549), .A2(n591), .ZN(n679) );
  INV_X1 U687 ( .A(n688), .ZN(n593) );
  INV_X1 U688 ( .A(n549), .ZN(n595) );
  NAND2_X1 U689 ( .A1(n595), .A2(n594), .ZN(n615) );
  NOR2_X1 U690 ( .A1(n598), .A2(n615), .ZN(n596) );
  NAND2_X1 U691 ( .A1(n597), .A2(n596), .ZN(n674) );
  NOR2_X1 U692 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U693 ( .A(KEYINPUT36), .B(n600), .Z(n601) );
  NOR2_X1 U694 ( .A1(n402), .A2(n601), .ZN(n682) );
  INV_X1 U695 ( .A(n682), .ZN(n602) );
  NOR2_X1 U696 ( .A1(n605), .A2(n606), .ZN(n684) );
  NAND2_X1 U697 ( .A1(n625), .A2(n633), .ZN(n610) );
  INV_X1 U698 ( .A(n611), .ZN(n628) );
  XNOR2_X1 U699 ( .A(KEYINPUT77), .B(n615), .ZN(n616) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U701 ( .A1(n697), .A2(n621), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n622), .A2(n628), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT96), .B(n623), .Z(n624) );
  NAND2_X1 U704 ( .A1(n624), .A2(n627), .ZN(n669) );
  INV_X1 U705 ( .A(n625), .ZN(n626) );
  NAND2_X1 U706 ( .A1(n628), .A2(n708), .ZN(n630) );
  XOR2_X1 U707 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n629) );
  NAND2_X1 U708 ( .A1(n632), .A2(n688), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n402), .A2(n700), .ZN(n634) );
  NOR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n665) );
  AND2_X1 U712 ( .A1(n637), .A2(n665), .ZN(n638) );
  INV_X1 U713 ( .A(KEYINPUT64), .ZN(n640) );
  NOR2_X2 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X2 U715 ( .A(n643), .B(KEYINPUT45), .ZN(n719) );
  OR2_X2 U716 ( .A1(n644), .A2(n719), .ZN(n722) );
  XNOR2_X1 U717 ( .A(n767), .B(KEYINPUT75), .ZN(n646) );
  NOR2_X1 U718 ( .A1(n646), .A2(n719), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n647), .A2(KEYINPUT2), .ZN(n648) );
  NOR2_X4 U720 ( .A1(n649), .A2(n648), .ZN(n735) );
  NAND2_X1 U721 ( .A1(n735), .A2(G210), .ZN(n654) );
  XOR2_X1 U722 ( .A(KEYINPUT86), .B(KEYINPUT54), .Z(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(KEYINPUT55), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n656) );
  INV_X1 U726 ( .A(G952), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n748), .ZN(n658) );
  XOR2_X1 U728 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n657) );
  XNOR2_X1 U729 ( .A(n658), .B(n657), .ZN(G51) );
  XNOR2_X1 U730 ( .A(KEYINPUT63), .B(KEYINPUT115), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n735), .A2(G472), .ZN(n661) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT62), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(G57) );
  XNOR2_X1 U735 ( .A(G101), .B(n665), .ZN(G3) );
  NOR2_X1 U736 ( .A1(n669), .A2(n677), .ZN(n666) );
  XOR2_X1 U737 ( .A(G104), .B(n666), .Z(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n668) );
  XNOR2_X1 U739 ( .A(G107), .B(KEYINPUT116), .ZN(n667) );
  XNOR2_X1 U740 ( .A(n668), .B(n667), .ZN(n671) );
  NOR2_X1 U741 ( .A1(n679), .A2(n669), .ZN(n670) );
  XOR2_X1 U742 ( .A(n671), .B(n670), .Z(G9) );
  NOR2_X1 U743 ( .A1(n675), .A2(n679), .ZN(n673) );
  XNOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .ZN(n672) );
  XNOR2_X1 U745 ( .A(n673), .B(n672), .ZN(G30) );
  XNOR2_X1 U746 ( .A(G143), .B(n674), .ZN(G45) );
  NOR2_X1 U747 ( .A1(n675), .A2(n677), .ZN(n676) );
  XOR2_X1 U748 ( .A(G146), .B(n676), .Z(G48) );
  NOR2_X1 U749 ( .A1(n680), .A2(n677), .ZN(n678) );
  XOR2_X1 U750 ( .A(G113), .B(n678), .Z(G15) );
  NOR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U752 ( .A(G116), .B(n681), .Z(G18) );
  XNOR2_X1 U753 ( .A(G125), .B(n682), .ZN(n683) );
  XNOR2_X1 U754 ( .A(n683), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U755 ( .A(G134), .B(n684), .ZN(n685) );
  XNOR2_X1 U756 ( .A(n685), .B(KEYINPUT117), .ZN(G36) );
  INV_X1 U757 ( .A(n686), .ZN(n690) );
  NAND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U762 ( .A1(n695), .A2(n725), .ZN(n712) );
  NAND2_X1 U763 ( .A1(n697), .A2(n402), .ZN(n698) );
  XNOR2_X1 U764 ( .A(KEYINPUT50), .B(n698), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U766 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n702), .B(n701), .ZN(n703) );
  NAND2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U770 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U771 ( .A(KEYINPUT51), .B(n709), .ZN(n710) );
  NAND2_X1 U772 ( .A1(n710), .A2(n724), .ZN(n711) );
  NAND2_X1 U773 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U774 ( .A(n713), .B(KEYINPUT52), .ZN(n714) );
  XNOR2_X1 U775 ( .A(n714), .B(KEYINPUT119), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U777 ( .A1(n717), .A2(G952), .ZN(n718) );
  XNOR2_X1 U778 ( .A(n718), .B(KEYINPUT120), .ZN(n729) );
  INV_X1 U779 ( .A(n719), .ZN(n757) );
  NAND2_X1 U780 ( .A1(n757), .A2(n767), .ZN(n720) );
  NAND2_X1 U781 ( .A1(n720), .A2(n370), .ZN(n721) );
  NAND2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U783 ( .A1(n723), .A2(n769), .ZN(n727) );
  AND2_X1 U784 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U785 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U786 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U787 ( .A(KEYINPUT53), .B(n730), .Z(G75) );
  XNOR2_X1 U788 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n731), .B(KEYINPUT57), .ZN(n732) );
  NOR2_X1 U790 ( .A1(n748), .A2(n734), .ZN(G54) );
  NAND2_X1 U791 ( .A1(n735), .A2(G475), .ZN(n738) );
  XOR2_X1 U792 ( .A(n736), .B(KEYINPUT59), .Z(n737) );
  XNOR2_X1 U793 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U794 ( .A1(n739), .A2(n748), .ZN(n740) );
  XNOR2_X1 U795 ( .A(n740), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U796 ( .A1(n744), .A2(G478), .ZN(n742) );
  XNOR2_X1 U797 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U798 ( .A1(n748), .A2(n743), .ZN(G63) );
  NAND2_X1 U799 ( .A1(n744), .A2(G217), .ZN(n745) );
  XNOR2_X1 U800 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(G66) );
  XOR2_X1 U802 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n749) );
  XNOR2_X1 U803 ( .A(n749), .B(G101), .ZN(n750) );
  XNOR2_X1 U804 ( .A(n751), .B(n750), .ZN(n752) );
  XOR2_X1 U805 ( .A(n753), .B(n752), .Z(n755) );
  NOR2_X1 U806 ( .A1(G898), .A2(n769), .ZN(n754) );
  NOR2_X1 U807 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U808 ( .A(KEYINPUT124), .B(n756), .ZN(n764) );
  NAND2_X1 U809 ( .A1(n757), .A2(n769), .ZN(n762) );
  XOR2_X1 U810 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n759) );
  NAND2_X1 U811 ( .A1(G224), .A2(G953), .ZN(n758) );
  XNOR2_X1 U812 ( .A(n759), .B(n758), .ZN(n760) );
  NAND2_X1 U813 ( .A1(n760), .A2(G898), .ZN(n761) );
  NAND2_X1 U814 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n764), .B(n763), .ZN(G69) );
  XNOR2_X1 U816 ( .A(n765), .B(n766), .ZN(n771) );
  INV_X1 U817 ( .A(n771), .ZN(n768) );
  XNOR2_X1 U818 ( .A(n768), .B(n767), .ZN(n770) );
  NAND2_X1 U819 ( .A1(n770), .A2(n769), .ZN(n775) );
  XNOR2_X1 U820 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U822 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U823 ( .A1(n775), .A2(n774), .ZN(G72) );
  XOR2_X1 U824 ( .A(n776), .B(G122), .Z(G24) );
  XOR2_X1 U825 ( .A(G137), .B(n777), .Z(G39) );
  XOR2_X1 U826 ( .A(n778), .B(G131), .Z(G33) );
endmodule

