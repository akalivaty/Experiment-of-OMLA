//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1115, new_n1116;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT66), .B(KEYINPUT67), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  OR2_X1    g033(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n465), .B2(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n464), .A2(new_n467), .A3(G125), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n461), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n459), .B(new_n460), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n477), .ZN(G160));
  INV_X1    g053(.A(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n464), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n461), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n464), .A2(new_n470), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n464), .A2(KEYINPUT70), .A3(new_n470), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n485), .B1(G136), .B2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(KEYINPUT71), .B(KEYINPUT72), .Z(new_n493));
  XNOR2_X1  g068(.A(new_n492), .B(new_n493), .ZN(G162));
  OAI21_X1  g069(.A(KEYINPUT73), .B1(new_n470), .B2(G114), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT73), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n464), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT4), .B1(new_n475), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n510));
  NAND4_X1  g085(.A1(new_n461), .A2(new_n510), .A3(new_n464), .A4(new_n507), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(G164));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n513), .A2(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT75), .ZN(new_n516));
  OAI21_X1  g091(.A(G651), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n519), .A2(new_n513), .ZN(new_n522));
  AOI22_X1  g097(.A1(G50), .A2(new_n521), .B1(new_n522), .B2(G88), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n517), .A2(KEYINPUT76), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  XNOR2_X1  g102(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n528));
  AND3_X1   g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n519), .A2(new_n513), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  INV_X1    g109(.A(G51), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n533), .A2(new_n534), .B1(new_n520), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n532), .A2(new_n536), .ZN(G168));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n533), .A2(new_n538), .B1(new_n520), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  XOR2_X1   g119(.A(KEYINPUT79), .B(G43), .Z(new_n545));
  AOI22_X1  g120(.A1(new_n521), .A2(new_n545), .B1(new_n522), .B2(G81), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n513), .A2(G56), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n542), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n546), .B1(new_n547), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n550), .A2(new_n547), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(new_n513), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n522), .B2(G91), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT80), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n564), .B(new_n565), .C1(new_n520), .C2(new_n566), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n566), .B1(KEYINPUT80), .B2(KEYINPUT9), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n521), .B(new_n568), .C1(KEYINPUT80), .C2(KEYINPUT9), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n563), .A2(new_n567), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  XOR2_X1   g146(.A(G168), .B(KEYINPUT81), .Z(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G286));
  OAI21_X1  g148(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI221_X1 g151(.A(new_n574), .B1(new_n533), .B2(new_n575), .C1(new_n576), .C2(new_n520), .ZN(G288));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n533), .A2(new_n578), .B1(new_n520), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n542), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(G47), .A2(new_n521), .B1(new_n522), .B2(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n542), .B2(new_n586), .ZN(G290));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NOR2_X1   g163(.A1(G301), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n522), .A2(G92), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n560), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n521), .B2(G54), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT82), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n589), .B1(new_n597), .B2(new_n588), .ZN(G284));
  AOI21_X1  g173(.A(new_n589), .B1(new_n597), .B2(new_n588), .ZN(G321));
  NOR2_X1   g174(.A1(G299), .A2(G868), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(new_n572), .B2(G868), .ZN(G297));
  XNOR2_X1  g176(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n597), .B1(new_n603), .B2(G860), .ZN(G148));
  NAND2_X1  g179(.A1(new_n597), .A2(new_n603), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OR3_X1    g181(.A1(new_n606), .A2(KEYINPUT84), .A3(new_n588), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT84), .B1(new_n606), .B2(new_n588), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(new_n608), .C1(G868), .C2(new_n553), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n464), .A2(new_n471), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n481), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n461), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n490), .C2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n614), .A2(G2100), .B1(new_n619), .B2(G2096), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(G2096), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n620), .B(new_n621), .C1(G2100), .C2(new_n614), .ZN(G156));
  XOR2_X1   g197(.A(KEYINPUT15), .B(G2435), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2438), .ZN(new_n624));
  XOR2_X1   g199(.A(G2427), .B(G2430), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT85), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n636), .A2(G14), .A3(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT17), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT86), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n640), .A2(new_n641), .ZN(new_n646));
  INV_X1    g221(.A(new_n639), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n646), .B(new_n643), .C1(new_n647), .C2(new_n641), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n641), .A3(new_n642), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2096), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  AOI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n656), .C2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G229));
  INV_X1    g245(.A(G16), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G6), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n583), .B2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT89), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT32), .B(G1981), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(G22), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT91), .Z(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(G166), .B2(new_n671), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(G1971), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(G1971), .ZN(new_n681));
  NOR2_X1   g256(.A1(G16), .A2(G23), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G288), .B2(new_n671), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n676), .A2(new_n680), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(KEYINPUT34), .ZN(new_n688));
  MUX2_X1   g263(.A(G24), .B(G290), .S(G16), .Z(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G1986), .Z(new_n690));
  NAND2_X1  g265(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(G25), .A2(G29), .ZN(new_n693));
  NOR2_X1   g268(.A1(G95), .A2(G2105), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT87), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n695), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT88), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n491), .A2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n481), .A2(G119), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n693), .B1(new_n701), .B2(G29), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT35), .B(G1991), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n702), .A2(new_n704), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n692), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n688), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(KEYINPUT34), .B2(new_n687), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n709), .A2(KEYINPUT92), .A3(KEYINPUT36), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(KEYINPUT92), .B2(KEYINPUT36), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT31), .B(G11), .Z(new_n712));
  INV_X1    g287(.A(G28), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(KEYINPUT30), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NOR2_X1   g292(.A1(G171), .A2(new_n671), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(G5), .B2(new_n671), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n716), .B1(new_n717), .B2(new_n619), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n671), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n671), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT97), .Z(new_n724));
  AOI21_X1  g299(.A(new_n721), .B1(new_n724), .B2(G1966), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G1966), .B2(new_n724), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(KEYINPUT98), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n719), .A2(new_n720), .ZN(new_n728));
  INV_X1    g303(.A(G2078), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n509), .A2(new_n511), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n499), .A2(new_n501), .B1(new_n464), .B2(new_n503), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n717), .A2(G27), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n729), .B2(new_n735), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n481), .A2(G129), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT26), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n741), .A2(new_n742), .B1(G105), .B2(new_n471), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n491), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G29), .ZN(new_n748));
  NOR2_X1   g323(.A1(G29), .A2(G32), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(KEYINPUT96), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(KEYINPUT96), .B2(new_n748), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT27), .B(G1996), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT24), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n717), .B1(new_n753), .B2(G34), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n753), .B2(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G160), .B2(G29), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n751), .A2(new_n752), .B1(G2084), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n717), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n481), .A2(G128), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT93), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n491), .A2(G140), .ZN(new_n762));
  OAI221_X1 g337(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n461), .C2(G116), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(G29), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT94), .B(G2067), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G19), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n553), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1341), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n727), .A2(new_n737), .A3(new_n757), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(KEYINPUT98), .B2(new_n726), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G35), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G162), .B2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT99), .B(KEYINPUT29), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G2090), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n717), .A2(G33), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT25), .Z(new_n781));
  INV_X1    g356(.A(G139), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n490), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n787));
  OAI22_X1  g362(.A1(new_n785), .A2(new_n786), .B1(new_n461), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n779), .B1(new_n788), .B2(G29), .ZN(new_n789));
  INV_X1    g364(.A(G2072), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n671), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT23), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n751), .A2(new_n752), .B1(G2084), .B2(new_n756), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n791), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(G4), .A2(G16), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(new_n597), .B2(G16), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1348), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n790), .B2(new_n789), .ZN(new_n802));
  AND3_X1   g377(.A1(new_n778), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n710), .A2(new_n711), .A3(new_n773), .A4(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  NAND2_X1  g380(.A1(new_n597), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G93), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT101), .B(G55), .ZN(new_n810));
  OAI22_X1  g385(.A1(new_n533), .A2(new_n809), .B1(new_n520), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(new_n542), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n553), .B(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n808), .B(new_n816), .Z(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n818));
  INV_X1    g393(.A(G860), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(KEYINPUT39), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n814), .A2(new_n819), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(G145));
  XOR2_X1   g399(.A(new_n700), .B(KEYINPUT103), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n612), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n464), .A2(new_n503), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n500), .B1(new_n495), .B2(new_n498), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT102), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n502), .A2(new_n504), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n730), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n788), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n826), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n764), .B(new_n746), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n481), .A2(G130), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n461), .A2(G118), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(G142), .B2(new_n491), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n835), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n834), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n619), .B(G160), .ZN(new_n843));
  XNOR2_X1  g418(.A(G162), .B(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(G37), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n842), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(G395));
  XNOR2_X1  g423(.A(G288), .B(KEYINPUT106), .ZN(new_n849));
  XNOR2_X1  g424(.A(G303), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(G290), .B(new_n583), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT107), .ZN(new_n855));
  MUX2_X1   g430(.A(new_n854), .B(new_n855), .S(KEYINPUT42), .Z(new_n856));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n857));
  INV_X1    g432(.A(G299), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n596), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n858), .B2(new_n596), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n596), .B2(new_n858), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OR3_X1    g437(.A1(new_n860), .A2(KEYINPUT41), .A3(new_n861), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT41), .B1(new_n860), .B2(new_n861), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n605), .B(new_n816), .ZN(new_n867));
  MUX2_X1   g442(.A(new_n862), .B(new_n866), .S(new_n867), .Z(new_n868));
  XNOR2_X1  g443(.A(new_n856), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G868), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n815), .A2(new_n588), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(G295));
  NOR2_X1   g447(.A1(G295), .A2(KEYINPUT108), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n870), .B2(new_n871), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(new_n875), .ZN(G331));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n877));
  NOR2_X1   g452(.A1(G168), .A2(G171), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n572), .B2(G171), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(new_n816), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n816), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n879), .A2(KEYINPUT109), .A3(new_n816), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n883), .A2(new_n864), .A3(new_n863), .A4(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT110), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n865), .A2(KEYINPUT110), .A3(new_n884), .A4(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n880), .A2(new_n881), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n862), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n887), .A2(new_n855), .A3(new_n888), .A4(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n892), .B2(KEYINPUT111), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n890), .B1(new_n885), .B2(new_n886), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT111), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n855), .A4(new_n888), .ZN(new_n896));
  INV_X1    g471(.A(new_n855), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n862), .B1(new_n883), .B2(new_n884), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n865), .A2(new_n889), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n893), .A2(new_n896), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n877), .B1(new_n901), .B2(KEYINPUT43), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n892), .A2(KEYINPUT111), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n897), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n896), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n902), .B1(KEYINPUT43), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n893), .A2(new_n910), .A3(new_n896), .A4(new_n900), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT112), .B1(new_n912), .B2(new_n877), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n914));
  AOI211_X1 g489(.A(new_n914), .B(KEYINPUT44), .C1(new_n909), .C2(new_n911), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n908), .B1(new_n913), .B2(new_n915), .ZN(G397));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n832), .A2(new_n917), .ZN(new_n918));
  XOR2_X1   g493(.A(KEYINPUT113), .B(KEYINPUT45), .Z(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G40), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n469), .A2(new_n921), .A3(new_n477), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G2067), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n764), .B(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G1996), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n746), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n924), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(KEYINPUT114), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n701), .A2(new_n703), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n700), .A2(new_n704), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n923), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G290), .B(G1986), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n923), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G8), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT45), .B1(new_n832), .B2(new_n917), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n466), .A2(new_n468), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n479), .ZN(new_n940));
  INV_X1    g515(.A(new_n477), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(G40), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT117), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT117), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n509), .A2(new_n511), .B1(new_n731), .B2(new_n830), .ZN(new_n945));
  AOI21_X1  g520(.A(G1384), .B1(new_n945), .B2(new_n829), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n944), .B(new_n922), .C1(new_n946), .C2(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n732), .A2(new_n917), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n948), .A2(new_n919), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n943), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1966), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G2084), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n832), .A2(new_n954), .A3(new_n917), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n922), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n937), .B1(new_n952), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(G168), .A2(new_n937), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n959), .A2(KEYINPUT51), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT123), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n952), .B2(new_n958), .ZN(new_n963));
  AOI211_X1 g538(.A(KEYINPUT123), .B(new_n957), .C1(new_n950), .C2(new_n951), .ZN(new_n964));
  OAI21_X1  g539(.A(G8), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT124), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT124), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(G8), .C1(new_n963), .C2(new_n964), .ZN(new_n968));
  INV_X1    g543(.A(new_n960), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n961), .B1(new_n970), .B2(KEYINPUT51), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT125), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT62), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT125), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n960), .B1(new_n965), .B2(KEYINPUT124), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n978), .B2(new_n968), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n976), .B(new_n972), .C1(new_n979), .C2(new_n961), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n974), .A2(new_n975), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n975), .B1(new_n974), .B2(new_n980), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n942), .A2(new_n918), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n983), .A2(new_n937), .ZN(new_n984));
  INV_X1    g559(.A(G1976), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(G288), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT52), .ZN(new_n987));
  NOR2_X1   g562(.A1(G305), .A2(G1981), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n989));
  AND2_X1   g564(.A1(G305), .A2(G1981), .ZN(new_n990));
  OR3_X1    g565(.A1(new_n988), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n988), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n984), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(G288), .B2(new_n985), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n984), .B(new_n994), .C1(new_n985), .C2(G288), .ZN(new_n995));
  AND3_X1   g570(.A1(new_n987), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n956), .A2(new_n922), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n955), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n999), .B2(G2090), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n942), .B1(KEYINPUT45), .B2(new_n946), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n948), .A2(new_n919), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1971), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G2090), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n998), .A2(KEYINPUT115), .A3(new_n1006), .A4(new_n955), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(G303), .A2(G8), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT55), .Z(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(G8), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n996), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1010), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n942), .B1(KEYINPUT50), .B2(new_n918), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1014), .A2(KEYINPUT116), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n948), .A2(KEYINPUT50), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1016), .B1(new_n1014), .B2(KEYINPUT116), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1005), .B1(new_n1018), .B2(G2090), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1012), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n950), .A2(G2078), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT126), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n1024), .B2(new_n1023), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1001), .A2(new_n729), .A3(new_n1002), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1027), .A2(new_n1022), .B1(new_n999), .B2(new_n720), .ZN(new_n1028));
  AOI21_X1  g603(.A(G301), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1021), .A2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n981), .A2(new_n982), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n974), .A2(new_n980), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n920), .A2(new_n1022), .A3(G2078), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1001), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G171), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1033), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1026), .A2(G301), .A3(new_n1028), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1033), .B1(new_n1036), .B2(G171), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1021), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1001), .A2(new_n927), .A3(new_n1002), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT58), .B(G1341), .Z(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n942), .B2(new_n918), .ZN(new_n1045));
  AOI211_X1 g620(.A(new_n552), .B(new_n551), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1047));
  XNOR2_X1  g622(.A(new_n1046), .B(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1348), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n999), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n983), .A2(new_n925), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n597), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1052), .A2(KEYINPUT60), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n597), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1053), .B(new_n1056), .C1(new_n1054), .C2(new_n597), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1048), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1001), .A2(new_n1002), .A3(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g637(.A(new_n1062), .B(KEYINPUT118), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1956), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(G299), .B(KEYINPUT57), .Z(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT120), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1064), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1062), .B(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1066), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1070), .A3(new_n1066), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1067), .A2(new_n1073), .A3(KEYINPUT61), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1065), .A2(new_n1076), .A3(new_n1066), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(KEYINPUT119), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1071), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1060), .B(new_n1075), .C1(KEYINPUT61), .C2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1067), .A2(new_n1073), .A3(new_n1053), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1042), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1032), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n993), .ZN(new_n1086));
  NOR3_X1   g661(.A1(new_n1086), .A2(G1976), .A3(G288), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n984), .B1(new_n1087), .B2(new_n988), .ZN(new_n1088));
  INV_X1    g663(.A(new_n996), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1011), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1021), .A2(new_n572), .A3(new_n959), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1010), .B1(new_n1008), .B2(G8), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1012), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n572), .A3(new_n959), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1085), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n936), .B1(new_n1031), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n930), .A2(new_n932), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n764), .A2(G2067), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n924), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n924), .A2(G1986), .A3(G290), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT48), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n934), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n923), .A2(new_n927), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT46), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n926), .A2(new_n747), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(new_n924), .ZN(new_n1109));
  XOR2_X1   g684(.A(new_n1109), .B(KEYINPUT47), .Z(new_n1110));
  NOR3_X1   g685(.A1(new_n1102), .A2(new_n1105), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT127), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1099), .A2(new_n1112), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g688(.A1(new_n653), .A2(G319), .ZN(new_n1115));
  NOR3_X1   g689(.A1(G229), .A2(G401), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g690(.A1(new_n846), .A2(new_n912), .A3(new_n1116), .ZN(G225));
  INV_X1    g691(.A(G225), .ZN(G308));
endmodule


