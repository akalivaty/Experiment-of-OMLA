

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744;

  AND2_X1 U361 ( .A1(n414), .A2(n408), .ZN(n406) );
  XOR2_X1 U362 ( .A(G131), .B(G113), .Z(n482) );
  BUF_X1 U363 ( .A(G107), .Z(n340) );
  XNOR2_X1 U364 ( .A(n418), .B(KEYINPUT3), .ZN(n456) );
  XNOR2_X1 U365 ( .A(n394), .B(G122), .ZN(n494) );
  XNOR2_X1 U366 ( .A(n490), .B(KEYINPUT4), .ZN(n465) );
  XNOR2_X1 U367 ( .A(n416), .B(G101), .ZN(n470) );
  NOR2_X2 U368 ( .A1(n625), .A2(n717), .ZN(n627) );
  NOR2_X2 U369 ( .A1(n639), .A2(n717), .ZN(n640) );
  XNOR2_X1 U370 ( .A(n341), .B(n514), .ZN(n520) );
  NAND2_X1 U371 ( .A1(n361), .A2(n363), .ZN(n341) );
  XNOR2_X2 U372 ( .A(n424), .B(n342), .ZN(n527) );
  XNOR2_X1 U373 ( .A(G122), .B(G104), .ZN(n481) );
  XNOR2_X1 U374 ( .A(G146), .B(n340), .ZN(n472) );
  INV_X1 U375 ( .A(n662), .ZN(n576) );
  NOR2_X2 U376 ( .A1(n631), .A2(n717), .ZN(n632) );
  NOR2_X2 U377 ( .A1(n612), .A2(n717), .ZN(n614) );
  NOR2_X2 U378 ( .A1(n527), .A2(n679), .ZN(n570) );
  NOR2_X1 U379 ( .A1(G953), .A2(G237), .ZN(n485) );
  NOR2_X1 U380 ( .A1(n557), .A2(n558), .ZN(n652) );
  NOR2_X2 U381 ( .A1(n556), .A2(n433), .ZN(n435) );
  NAND2_X1 U382 ( .A1(n344), .A2(n665), .ZN(n354) );
  XNOR2_X1 U383 ( .A(n537), .B(KEYINPUT42), .ZN(n744) );
  NOR2_X1 U384 ( .A1(n693), .A2(n557), .ZN(n537) );
  XNOR2_X1 U385 ( .A(n590), .B(n528), .ZN(n684) );
  XNOR2_X1 U386 ( .A(n364), .B(n476), .ZN(n536) );
  XNOR2_X1 U387 ( .A(n451), .B(n391), .ZN(n665) );
  NOR2_X1 U388 ( .A1(n609), .A2(G902), .ZN(n451) );
  XNOR2_X1 U389 ( .A(n634), .B(n636), .ZN(n637) );
  XNOR2_X1 U390 ( .A(n356), .B(n345), .ZN(n516) );
  XOR2_X1 U391 ( .A(n628), .B(KEYINPUT59), .Z(n629) );
  XNOR2_X1 U392 ( .A(n454), .B(KEYINPUT21), .ZN(n666) );
  XNOR2_X1 U393 ( .A(n450), .B(KEYINPUT20), .ZN(n453) );
  XNOR2_X1 U394 ( .A(n494), .B(n417), .ZN(n369) );
  XNOR2_X1 U395 ( .A(n456), .B(n470), .ZN(n370) );
  XNOR2_X1 U396 ( .A(n377), .B(n421), .ZN(n600) );
  XOR2_X1 U397 ( .A(KEYINPUT16), .B(KEYINPUT74), .Z(n417) );
  INV_X1 U398 ( .A(G953), .ZN(n436) );
  XNOR2_X1 U399 ( .A(G902), .B(KEYINPUT85), .ZN(n377) );
  XNOR2_X1 U400 ( .A(n465), .B(n464), .ZN(n469) );
  XNOR2_X1 U401 ( .A(G134), .B(G131), .ZN(n463) );
  XNOR2_X1 U402 ( .A(n390), .B(n389), .ZN(n573) );
  INV_X1 U403 ( .A(KEYINPUT70), .ZN(n389) );
  NOR2_X1 U404 ( .A1(n665), .A2(n534), .ZN(n390) );
  XNOR2_X1 U405 ( .A(n536), .B(KEYINPUT1), .ZN(n662) );
  XNOR2_X1 U406 ( .A(n384), .B(G146), .ZN(n448) );
  INV_X1 U407 ( .A(G125), .ZN(n384) );
  NAND2_X1 U408 ( .A1(G237), .A2(G234), .ZN(n429) );
  INV_X1 U409 ( .A(G210), .ZN(n422) );
  NOR2_X1 U410 ( .A1(n544), .A2(n543), .ZN(n560) );
  OR2_X1 U411 ( .A1(n714), .A2(G902), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n488), .B(n387), .ZN(n517) );
  XNOR2_X1 U413 ( .A(n487), .B(G475), .ZN(n387) );
  XNOR2_X1 U414 ( .A(n379), .B(n378), .ZN(n391) );
  XNOR2_X1 U415 ( .A(n452), .B(KEYINPUT77), .ZN(n378) );
  XNOR2_X1 U416 ( .A(n466), .B(n469), .ZN(n622) );
  XNOR2_X1 U417 ( .A(n494), .B(KEYINPUT9), .ZN(n495) );
  XNOR2_X1 U418 ( .A(n439), .B(n438), .ZN(n489) );
  XNOR2_X1 U419 ( .A(n437), .B(KEYINPUT81), .ZN(n439) );
  NAND2_X1 U420 ( .A1(G234), .A2(n436), .ZN(n437) );
  XNOR2_X1 U421 ( .A(n448), .B(n383), .ZN(n729) );
  XNOR2_X1 U422 ( .A(KEYINPUT10), .B(G140), .ZN(n383) );
  XNOR2_X1 U423 ( .A(n343), .B(n483), .ZN(n381) );
  INV_X1 U424 ( .A(KEYINPUT64), .ZN(n607) );
  XNOR2_X1 U425 ( .A(n512), .B(KEYINPUT33), .ZN(n363) );
  BUF_X1 U426 ( .A(n603), .Z(n733) );
  XNOR2_X1 U427 ( .A(n360), .B(KEYINPUT41), .ZN(n693) );
  NOR2_X1 U428 ( .A1(n678), .A2(n684), .ZN(n360) );
  INV_X1 U429 ( .A(KEYINPUT32), .ZN(n402) );
  NOR2_X1 U430 ( .A1(n499), .A2(n376), .ZN(n375) );
  OR2_X1 U431 ( .A1(n708), .A2(G902), .ZN(n364) );
  BUF_X1 U432 ( .A(n665), .Z(n355) );
  XNOR2_X1 U433 ( .A(n551), .B(n349), .ZN(n552) );
  NAND2_X1 U434 ( .A1(n652), .A2(n559), .ZN(n569) );
  INV_X1 U435 ( .A(KEYINPUT15), .ZN(n421) );
  INV_X1 U436 ( .A(KEYINPUT65), .ZN(n412) );
  NAND2_X1 U437 ( .A1(n411), .A2(n409), .ZN(n408) );
  NAND2_X1 U438 ( .A1(n601), .A2(n410), .ZN(n409) );
  NAND2_X1 U439 ( .A1(n413), .A2(n412), .ZN(n411) );
  NAND2_X1 U440 ( .A1(KEYINPUT2), .A2(n412), .ZN(n410) );
  INV_X1 U441 ( .A(n601), .ZN(n413) );
  OR2_X1 U442 ( .A1(G237), .A2(G902), .ZN(n425) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n682) );
  INV_X1 U444 ( .A(KEYINPUT99), .ZN(n385) );
  NOR2_X1 U445 ( .A1(n516), .A2(n517), .ZN(n386) );
  NAND2_X1 U446 ( .A1(n453), .A2(G217), .ZN(n379) );
  XNOR2_X1 U447 ( .A(G116), .B(G101), .ZN(n457) );
  XNOR2_X1 U448 ( .A(n419), .B(KEYINPUT18), .ZN(n367) );
  NAND2_X1 U449 ( .A1(n682), .A2(n586), .ZN(n678) );
  NAND2_X1 U450 ( .A1(n682), .A2(n344), .ZN(n376) );
  INV_X1 U451 ( .A(G902), .ZN(n467) );
  XNOR2_X1 U452 ( .A(n365), .B(n718), .ZN(n633) );
  XNOR2_X1 U453 ( .A(n368), .B(n366), .ZN(n365) );
  XNOR2_X1 U454 ( .A(n420), .B(n367), .ZN(n366) );
  XNOR2_X1 U455 ( .A(n465), .B(n448), .ZN(n368) );
  AND2_X1 U456 ( .A1(n697), .A2(n605), .ZN(n699) );
  INV_X1 U457 ( .A(KEYINPUT102), .ZN(n373) );
  XNOR2_X1 U458 ( .A(n427), .B(KEYINPUT19), .ZN(n428) );
  NAND2_X1 U459 ( .A1(n358), .A2(n538), .ZN(n557) );
  XNOR2_X1 U460 ( .A(n359), .B(KEYINPUT28), .ZN(n358) );
  NOR2_X1 U461 ( .A1(n573), .A2(n535), .ZN(n359) );
  BUF_X1 U462 ( .A(n670), .Z(n372) );
  XNOR2_X1 U463 ( .A(n622), .B(n621), .ZN(n623) );
  BUF_X1 U464 ( .A(n436), .Z(n734) );
  XNOR2_X1 U465 ( .A(n449), .B(n729), .ZN(n609) );
  XNOR2_X1 U466 ( .A(n357), .B(n493), .ZN(n714) );
  XNOR2_X1 U467 ( .A(n495), .B(n492), .ZN(n357) );
  XNOR2_X1 U468 ( .A(n382), .B(n380), .ZN(n628) );
  XNOR2_X1 U469 ( .A(n381), .B(n484), .ZN(n380) );
  XNOR2_X1 U470 ( .A(n486), .B(n729), .ZN(n382) );
  XNOR2_X1 U471 ( .A(n731), .B(n475), .ZN(n708) );
  INV_X1 U472 ( .A(n693), .ZN(n362) );
  NAND2_X1 U473 ( .A1(n398), .A2(n397), .ZN(n396) );
  NOR2_X1 U474 ( .A1(n505), .A2(n402), .ZN(n397) );
  AND2_X1 U475 ( .A1(n401), .A2(n400), .ZN(n399) );
  XNOR2_X1 U476 ( .A(n393), .B(n392), .ZN(n658) );
  INV_X1 U477 ( .A(KEYINPUT31), .ZN(n392) );
  XNOR2_X1 U478 ( .A(n552), .B(n353), .ZN(G33) );
  OR2_X1 U479 ( .A1(n423), .A2(n422), .ZN(n342) );
  AND2_X1 U480 ( .A1(n485), .A2(G214), .ZN(n343) );
  XOR2_X1 U481 ( .A(n666), .B(KEYINPUT92), .Z(n344) );
  XOR2_X1 U482 ( .A(KEYINPUT97), .B(G478), .Z(n345) );
  OR2_X1 U483 ( .A1(n686), .A2(n685), .ZN(n346) );
  BUF_X1 U484 ( .A(n527), .Z(n590) );
  NAND2_X1 U485 ( .A1(n509), .A2(n572), .ZN(n506) );
  AND2_X1 U486 ( .A1(n346), .A2(n363), .ZN(n347) );
  AND2_X1 U487 ( .A1(n395), .A2(n396), .ZN(n348) );
  XOR2_X1 U488 ( .A(n550), .B(KEYINPUT40), .Z(n349) );
  XNOR2_X1 U489 ( .A(KEYINPUT36), .B(KEYINPUT84), .ZN(n350) );
  XOR2_X1 U490 ( .A(n500), .B(KEYINPUT66), .Z(n351) );
  XNOR2_X1 U491 ( .A(n370), .B(n369), .ZN(n718) );
  AND2_X1 U492 ( .A1(n601), .A2(n412), .ZN(n352) );
  XNOR2_X1 U493 ( .A(G131), .B(KEYINPUT126), .ZN(n353) );
  XNOR2_X1 U494 ( .A(n548), .B(n547), .ZN(n595) );
  XNOR2_X2 U495 ( .A(n354), .B(n455), .ZN(n539) );
  NAND2_X1 U496 ( .A1(n404), .A2(n606), .ZN(n608) );
  XNOR2_X2 U497 ( .A(G143), .B(G128), .ZN(n490) );
  INV_X1 U498 ( .A(n513), .ZN(n361) );
  AND2_X1 U499 ( .A1(n363), .A2(n362), .ZN(n694) );
  XNOR2_X1 U500 ( .A(n371), .B(n350), .ZN(n577) );
  AND2_X1 U501 ( .A1(n588), .A2(n570), .ZN(n371) );
  XNOR2_X1 U502 ( .A(n374), .B(n373), .ZN(n574) );
  NOR2_X1 U503 ( .A1(n572), .A2(n573), .ZN(n374) );
  XNOR2_X1 U504 ( .A(n375), .B(n351), .ZN(n509) );
  XNOR2_X2 U505 ( .A(n435), .B(n434), .ZN(n499) );
  NAND2_X1 U506 ( .A1(n617), .A2(n388), .ZN(n568) );
  NAND2_X1 U507 ( .A1(n569), .A2(KEYINPUT47), .ZN(n388) );
  NOR2_X1 U508 ( .A1(n499), .A2(n673), .ZN(n393) );
  XNOR2_X2 U509 ( .A(G116), .B(G107), .ZN(n394) );
  NOR2_X2 U510 ( .A1(n619), .A2(n403), .ZN(n523) );
  INV_X1 U511 ( .A(n618), .ZN(n395) );
  NAND2_X1 U512 ( .A1(n348), .A2(n399), .ZN(n403) );
  XNOR2_X2 U513 ( .A(n468), .B(G472), .ZN(n670) );
  NAND2_X1 U514 ( .A1(n407), .A2(n352), .ZN(n405) );
  NOR2_X1 U515 ( .A1(n497), .A2(n680), .ZN(n498) );
  NAND2_X1 U516 ( .A1(n399), .A2(n396), .ZN(n743) );
  INV_X1 U517 ( .A(n506), .ZN(n398) );
  NAND2_X1 U518 ( .A1(n505), .A2(n402), .ZN(n400) );
  NAND2_X1 U519 ( .A1(n506), .A2(n402), .ZN(n401) );
  NAND2_X1 U520 ( .A1(n406), .A2(n405), .ZN(n404) );
  INV_X1 U521 ( .A(n599), .ZN(n407) );
  NAND2_X1 U522 ( .A1(n599), .A2(n415), .ZN(n414) );
  AND2_X1 U523 ( .A1(n604), .A2(KEYINPUT65), .ZN(n415) );
  INV_X1 U524 ( .A(KEYINPUT17), .ZN(n419) );
  XNOR2_X1 U525 ( .A(n522), .B(n521), .ZN(n619) );
  INV_X1 U526 ( .A(KEYINPUT121), .ZN(n613) );
  BUF_X1 U527 ( .A(n619), .Z(n620) );
  XNOR2_X2 U528 ( .A(G110), .B(G104), .ZN(n416) );
  XNOR2_X2 U529 ( .A(G119), .B(G113), .ZN(n418) );
  NAND2_X1 U530 ( .A1(G224), .A2(n734), .ZN(n420) );
  NAND2_X1 U531 ( .A1(n633), .A2(n413), .ZN(n424) );
  INV_X1 U532 ( .A(n425), .ZN(n423) );
  NAND2_X1 U533 ( .A1(n425), .A2(G214), .ZN(n426) );
  XOR2_X1 U534 ( .A(KEYINPUT86), .B(n426), .Z(n679) );
  XOR2_X1 U535 ( .A(KEYINPUT76), .B(KEYINPUT67), .Z(n427) );
  XNOR2_X1 U536 ( .A(n570), .B(n428), .ZN(n556) );
  XNOR2_X1 U537 ( .A(n429), .B(KEYINPUT14), .ZN(n430) );
  NAND2_X1 U538 ( .A1(G952), .A2(n430), .ZN(n692) );
  NOR2_X1 U539 ( .A1(n692), .A2(G953), .ZN(n532) );
  NAND2_X1 U540 ( .A1(G902), .A2(n430), .ZN(n529) );
  INV_X1 U541 ( .A(G898), .ZN(n723) );
  NAND2_X1 U542 ( .A1(G953), .A2(n723), .ZN(n719) );
  NOR2_X1 U543 ( .A1(n529), .A2(n719), .ZN(n431) );
  NOR2_X1 U544 ( .A1(n532), .A2(n431), .ZN(n432) );
  XOR2_X1 U545 ( .A(KEYINPUT87), .B(n432), .Z(n433) );
  INV_X1 U546 ( .A(KEYINPUT0), .ZN(n434) );
  XOR2_X1 U547 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n438) );
  NAND2_X1 U548 ( .A1(n489), .A2(G221), .ZN(n447) );
  XOR2_X1 U549 ( .A(G137), .B(G128), .Z(n441) );
  XNOR2_X1 U550 ( .A(G110), .B(G119), .ZN(n440) );
  XNOR2_X1 U551 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U552 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n443) );
  XNOR2_X1 U553 ( .A(KEYINPUT90), .B(KEYINPUT91), .ZN(n442) );
  XNOR2_X1 U554 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U555 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U556 ( .A(n447), .B(n446), .ZN(n449) );
  NAND2_X1 U557 ( .A1(G234), .A2(n600), .ZN(n450) );
  INV_X1 U558 ( .A(KEYINPUT25), .ZN(n452) );
  NAND2_X1 U559 ( .A1(n453), .A2(G221), .ZN(n454) );
  INV_X1 U560 ( .A(KEYINPUT68), .ZN(n455) );
  INV_X1 U561 ( .A(n539), .ZN(n663) );
  XNOR2_X1 U562 ( .A(n456), .B(n457), .ZN(n462) );
  XOR2_X1 U563 ( .A(G146), .B(KEYINPUT5), .Z(n459) );
  NAND2_X1 U564 ( .A1(n485), .A2(G210), .ZN(n458) );
  XNOR2_X1 U565 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U566 ( .A(n460), .B(KEYINPUT93), .Z(n461) );
  XNOR2_X1 U567 ( .A(n461), .B(n462), .ZN(n466) );
  XNOR2_X1 U568 ( .A(n463), .B(G137), .ZN(n464) );
  NAND2_X1 U569 ( .A1(n622), .A2(n467), .ZN(n468) );
  INV_X1 U570 ( .A(n670), .ZN(n535) );
  NOR2_X1 U571 ( .A1(n663), .A2(n535), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n469), .B(KEYINPUT89), .ZN(n731) );
  NAND2_X1 U573 ( .A1(n734), .A2(G227), .ZN(n471) );
  XNOR2_X1 U574 ( .A(n471), .B(G140), .ZN(n473) );
  XNOR2_X1 U575 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U576 ( .A(n470), .B(n474), .ZN(n475) );
  INV_X1 U577 ( .A(G469), .ZN(n476) );
  NAND2_X1 U578 ( .A1(n477), .A2(n576), .ZN(n673) );
  XNOR2_X1 U579 ( .A(n499), .B(KEYINPUT88), .ZN(n513) );
  NOR2_X1 U580 ( .A1(n372), .A2(n536), .ZN(n478) );
  NAND2_X1 U581 ( .A1(n539), .A2(n478), .ZN(n479) );
  NOR2_X1 U582 ( .A1(n513), .A2(n479), .ZN(n644) );
  NOR2_X1 U583 ( .A1(n658), .A2(n644), .ZN(n480) );
  XNOR2_X1 U584 ( .A(n480), .B(KEYINPUT94), .ZN(n497) );
  XNOR2_X1 U585 ( .A(n482), .B(n481), .ZN(n486) );
  XOR2_X1 U586 ( .A(KEYINPUT95), .B(KEYINPUT11), .Z(n484) );
  XNOR2_X1 U587 ( .A(G143), .B(KEYINPUT12), .ZN(n483) );
  NOR2_X1 U588 ( .A1(G902), .A2(n628), .ZN(n488) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n487) );
  NAND2_X1 U590 ( .A1(n489), .A2(G217), .ZN(n493) );
  XNOR2_X1 U591 ( .A(G134), .B(KEYINPUT7), .ZN(n491) );
  XNOR2_X1 U592 ( .A(n490), .B(n491), .ZN(n492) );
  INV_X1 U593 ( .A(n516), .ZN(n496) );
  OR2_X1 U594 ( .A1(n517), .A2(n496), .ZN(n594) );
  NAND2_X1 U595 ( .A1(n517), .A2(n496), .ZN(n571) );
  AND2_X1 U596 ( .A1(n594), .A2(n571), .ZN(n680) );
  XNOR2_X1 U597 ( .A(n498), .B(KEYINPUT98), .ZN(n504) );
  XNOR2_X1 U598 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n500) );
  XNOR2_X1 U599 ( .A(n670), .B(KEYINPUT6), .ZN(n572) );
  NOR2_X1 U600 ( .A1(n506), .A2(n576), .ZN(n502) );
  INV_X1 U601 ( .A(KEYINPUT83), .ZN(n501) );
  XNOR2_X1 U602 ( .A(n502), .B(n501), .ZN(n503) );
  AND2_X1 U603 ( .A1(n503), .A2(n355), .ZN(n641) );
  NOR2_X1 U604 ( .A1(n504), .A2(n641), .ZN(n525) );
  OR2_X1 U605 ( .A1(n662), .A2(n355), .ZN(n505) );
  NOR2_X1 U606 ( .A1(n355), .A2(n372), .ZN(n507) );
  AND2_X1 U607 ( .A1(n507), .A2(n662), .ZN(n508) );
  AND2_X1 U608 ( .A1(n509), .A2(n508), .ZN(n618) );
  INV_X1 U609 ( .A(n572), .ZN(n510) );
  AND2_X1 U610 ( .A1(n539), .A2(n510), .ZN(n511) );
  NAND2_X1 U611 ( .A1(n511), .A2(n576), .ZN(n512) );
  INV_X1 U612 ( .A(KEYINPUT34), .ZN(n514) );
  NAND2_X1 U613 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U614 ( .A(n518), .B(KEYINPUT100), .ZN(n565) );
  XNOR2_X1 U615 ( .A(n565), .B(KEYINPUT79), .ZN(n519) );
  NAND2_X1 U616 ( .A1(n520), .A2(n519), .ZN(n522) );
  XNOR2_X1 U617 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n521) );
  XNOR2_X1 U618 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  NAND2_X1 U619 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U620 ( .A(n526), .B(KEYINPUT45), .ZN(n602) );
  INV_X1 U621 ( .A(KEYINPUT38), .ZN(n528) );
  INV_X1 U622 ( .A(n679), .ZN(n586) );
  OR2_X1 U623 ( .A1(n734), .A2(n529), .ZN(n530) );
  NOR2_X1 U624 ( .A1(n530), .A2(G900), .ZN(n531) );
  NOR2_X1 U625 ( .A1(n532), .A2(n531), .ZN(n543) );
  NOR2_X1 U626 ( .A1(n666), .A2(n543), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n533), .B(KEYINPUT71), .ZN(n534) );
  INV_X1 U628 ( .A(n536), .ZN(n538) );
  INV_X1 U629 ( .A(n744), .ZN(n553) );
  NAND2_X1 U630 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U631 ( .A(KEYINPUT104), .ZN(n540) );
  XNOR2_X1 U632 ( .A(n541), .B(n540), .ZN(n561) );
  NAND2_X1 U633 ( .A1(n670), .A2(n586), .ZN(n542) );
  XNOR2_X1 U634 ( .A(n542), .B(KEYINPUT30), .ZN(n544) );
  INV_X1 U635 ( .A(n684), .ZN(n545) );
  AND2_X1 U636 ( .A1(n545), .A2(n560), .ZN(n546) );
  NAND2_X1 U637 ( .A1(n561), .A2(n546), .ZN(n548) );
  XNOR2_X1 U638 ( .A(KEYINPUT72), .B(KEYINPUT39), .ZN(n547) );
  INV_X1 U639 ( .A(n571), .ZN(n549) );
  NAND2_X1 U640 ( .A1(n595), .A2(n549), .ZN(n551) );
  INV_X1 U641 ( .A(KEYINPUT106), .ZN(n550) );
  NAND2_X1 U642 ( .A1(n553), .A2(n552), .ZN(n555) );
  INV_X1 U643 ( .A(KEYINPUT46), .ZN(n554) );
  XNOR2_X1 U644 ( .A(n555), .B(n554), .ZN(n582) );
  BUF_X1 U645 ( .A(n556), .Z(n558) );
  INV_X1 U646 ( .A(n680), .ZN(n559) );
  AND2_X1 U647 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U648 ( .A(n590), .ZN(n562) );
  NAND2_X1 U649 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n564), .B(KEYINPUT105), .ZN(n567) );
  INV_X1 U651 ( .A(n565), .ZN(n566) );
  NAND2_X1 U652 ( .A1(n567), .A2(n566), .ZN(n617) );
  XNOR2_X1 U653 ( .A(n568), .B(KEYINPUT80), .ZN(n580) );
  OR2_X1 U654 ( .A1(n569), .A2(KEYINPUT47), .ZN(n578) );
  XNOR2_X1 U655 ( .A(n571), .B(KEYINPUT101), .ZN(n655) );
  INV_X1 U656 ( .A(n655), .ZN(n575) );
  NOR2_X1 U657 ( .A1(n575), .A2(n574), .ZN(n588) );
  NAND2_X1 U658 ( .A1(n577), .A2(n576), .ZN(n660) );
  NAND2_X1 U659 ( .A1(n578), .A2(n660), .ZN(n579) );
  NOR2_X1 U660 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n585) );
  INV_X1 U662 ( .A(KEYINPUT82), .ZN(n583) );
  XNOR2_X1 U663 ( .A(n583), .B(KEYINPUT48), .ZN(n584) );
  XNOR2_X1 U664 ( .A(n585), .B(n584), .ZN(n597) );
  AND2_X1 U665 ( .A1(n662), .A2(n586), .ZN(n587) );
  NAND2_X1 U666 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U667 ( .A(n589), .B(KEYINPUT43), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n593) );
  INV_X1 U669 ( .A(KEYINPUT103), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n593), .B(n592), .ZN(n742) );
  INV_X1 U671 ( .A(n594), .ZN(n657) );
  NAND2_X1 U672 ( .A1(n595), .A2(n657), .ZN(n615) );
  AND2_X1 U673 ( .A1(n742), .A2(n615), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT75), .ZN(n598) );
  NAND2_X1 U676 ( .A1(n602), .A2(n598), .ZN(n599) );
  INV_X1 U677 ( .A(KEYINPUT2), .ZN(n604) );
  INV_X1 U678 ( .A(n600), .ZN(n601) );
  BUF_X1 U679 ( .A(n602), .Z(n697) );
  NOR2_X1 U680 ( .A1(n733), .A2(n604), .ZN(n605) );
  INV_X1 U681 ( .A(n699), .ZN(n606) );
  XNOR2_X2 U682 ( .A(n608), .B(n607), .ZN(n705) );
  NAND2_X1 U683 ( .A1(n705), .A2(G217), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(n609), .ZN(n612) );
  INV_X1 U685 ( .A(G952), .ZN(n611) );
  AND2_X1 U686 ( .A1(n611), .A2(G953), .ZN(n717) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(G66) );
  XNOR2_X1 U688 ( .A(n615), .B(G134), .ZN(G36) );
  XNOR2_X1 U689 ( .A(G143), .B(KEYINPUT112), .ZN(n616) );
  XNOR2_X1 U690 ( .A(n617), .B(n616), .ZN(G45) );
  XOR2_X1 U691 ( .A(n618), .B(G110), .Z(G12) );
  XOR2_X1 U692 ( .A(n620), .B(G122), .Z(G24) );
  NAND2_X1 U693 ( .A1(n705), .A2(G472), .ZN(n624) );
  XNOR2_X1 U694 ( .A(KEYINPUT107), .B(KEYINPUT62), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(n625) );
  XOR2_X1 U696 ( .A(KEYINPUT108), .B(KEYINPUT63), .Z(n626) );
  XNOR2_X1 U697 ( .A(n627), .B(n626), .ZN(G57) );
  NAND2_X1 U698 ( .A1(n705), .A2(G475), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n632), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U701 ( .A1(n705), .A2(G210), .ZN(n638) );
  BUF_X1 U702 ( .A(n633), .Z(n634) );
  XNOR2_X1 U703 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n635) );
  XNOR2_X1 U704 ( .A(n635), .B(KEYINPUT55), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n640), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U707 ( .A(G101), .B(n641), .ZN(n642) );
  XNOR2_X1 U708 ( .A(n642), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U709 ( .A1(n644), .A2(n655), .ZN(n643) );
  XNOR2_X1 U710 ( .A(n643), .B(G104), .ZN(G6) );
  XNOR2_X1 U711 ( .A(n340), .B(KEYINPUT27), .ZN(n648) );
  XOR2_X1 U712 ( .A(KEYINPUT26), .B(KEYINPUT110), .Z(n646) );
  NAND2_X1 U713 ( .A1(n644), .A2(n657), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n648), .B(n647), .ZN(G9) );
  XOR2_X1 U716 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n650) );
  NAND2_X1 U717 ( .A1(n652), .A2(n657), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U719 ( .A(G128), .B(n651), .Z(G30) );
  XOR2_X1 U720 ( .A(G146), .B(KEYINPUT113), .Z(n654) );
  NAND2_X1 U721 ( .A1(n652), .A2(n655), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(G48) );
  NAND2_X1 U723 ( .A1(n658), .A2(n655), .ZN(n656) );
  XNOR2_X1 U724 ( .A(n656), .B(G113), .ZN(G15) );
  NAND2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n659), .B(G116), .ZN(G18) );
  XOR2_X1 U727 ( .A(G125), .B(n660), .Z(n661) );
  XNOR2_X1 U728 ( .A(n661), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U729 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n676) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n664), .B(KEYINPUT50), .ZN(n672) );
  INV_X1 U732 ( .A(n355), .ZN(n667) );
  NAND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U734 ( .A(KEYINPUT49), .B(n668), .ZN(n669) );
  NOR2_X1 U735 ( .A1(n372), .A2(n669), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U738 ( .A(n676), .B(n675), .Z(n677) );
  NOR2_X1 U739 ( .A1(n693), .A2(n677), .ZN(n688) );
  INV_X1 U740 ( .A(n678), .ZN(n686) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U744 ( .A(KEYINPUT115), .B(n347), .Z(n687) );
  NOR2_X1 U745 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U746 ( .A(KEYINPUT52), .B(n689), .Z(n690) );
  XOR2_X1 U747 ( .A(KEYINPUT116), .B(n690), .Z(n691) );
  NOR2_X1 U748 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U749 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U750 ( .A(KEYINPUT117), .B(n696), .Z(n702) );
  INV_X1 U751 ( .A(n697), .ZN(n720) );
  NOR2_X1 U752 ( .A1(n720), .A2(n733), .ZN(n698) );
  NOR2_X1 U753 ( .A1(n698), .A2(KEYINPUT2), .ZN(n700) );
  OR2_X1 U754 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U755 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U756 ( .A1(n703), .A2(G953), .ZN(n704) );
  XNOR2_X1 U757 ( .A(n704), .B(KEYINPUT53), .ZN(G75) );
  BUF_X1 U758 ( .A(n705), .Z(n713) );
  NAND2_X1 U759 ( .A1(n713), .A2(G469), .ZN(n711) );
  XOR2_X1 U760 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n707) );
  XNOR2_X1 U761 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n706) );
  XNOR2_X1 U762 ( .A(n707), .B(n706), .ZN(n709) );
  XOR2_X1 U763 ( .A(n709), .B(n708), .Z(n710) );
  XNOR2_X1 U764 ( .A(n711), .B(n710), .ZN(n712) );
  NOR2_X1 U765 ( .A1(n717), .A2(n712), .ZN(G54) );
  NAND2_X1 U766 ( .A1(n713), .A2(G478), .ZN(n715) );
  XNOR2_X1 U767 ( .A(n714), .B(n715), .ZN(n716) );
  NOR2_X1 U768 ( .A1(n717), .A2(n716), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n719), .A2(n718), .ZN(n728) );
  NOR2_X1 U770 ( .A1(n720), .A2(G953), .ZN(n726) );
  XOR2_X1 U771 ( .A(KEYINPUT122), .B(KEYINPUT61), .Z(n722) );
  NAND2_X1 U772 ( .A1(G224), .A2(G953), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n722), .B(n721), .ZN(n724) );
  NOR2_X1 U774 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U775 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U776 ( .A(n728), .B(n727), .ZN(G69) );
  XNOR2_X1 U777 ( .A(n729), .B(KEYINPUT123), .ZN(n730) );
  XNOR2_X1 U778 ( .A(n731), .B(n730), .ZN(n736) );
  XNOR2_X1 U779 ( .A(n736), .B(KEYINPUT124), .ZN(n732) );
  XNOR2_X1 U780 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U781 ( .A1(n735), .A2(n734), .ZN(n740) );
  XNOR2_X1 U782 ( .A(G227), .B(n736), .ZN(n737) );
  NAND2_X1 U783 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U784 ( .A1(G953), .A2(n738), .ZN(n739) );
  NAND2_X1 U785 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U786 ( .A(KEYINPUT125), .B(n741), .Z(G72) );
  XNOR2_X1 U787 ( .A(G140), .B(n742), .ZN(G42) );
  XOR2_X1 U788 ( .A(G119), .B(n743), .Z(G21) );
  XOR2_X1 U789 ( .A(n744), .B(G137), .Z(G39) );
endmodule

