

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U323 ( .A(KEYINPUT65), .B(KEYINPUT10), .Z(n291) );
  INV_X1 U324 ( .A(KEYINPUT45), .ZN(n416) );
  XNOR2_X1 U325 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U326 ( .A(n306), .B(n374), .ZN(n307) );
  XNOR2_X1 U327 ( .A(n308), .B(n307), .ZN(n309) );
  NOR2_X1 U328 ( .A1(n531), .A2(n447), .ZN(n563) );
  XNOR2_X1 U329 ( .A(n328), .B(n327), .ZN(n531) );
  XNOR2_X1 U330 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n448) );
  XNOR2_X1 U331 ( .A(n449), .B(n448), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n293) );
  XNOR2_X1 U333 ( .A(G43GAT), .B(G29GAT), .ZN(n292) );
  XNOR2_X1 U334 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U335 ( .A(KEYINPUT69), .B(n294), .Z(n361) );
  XOR2_X1 U336 ( .A(G92GAT), .B(G106GAT), .Z(n296) );
  XNOR2_X1 U337 ( .A(G134GAT), .B(G218GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n299) );
  XNOR2_X1 U339 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n291), .B(n297), .ZN(n298) );
  XOR2_X1 U341 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U342 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n301) );
  NAND2_X1 U343 ( .A1(G232GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U345 ( .A(KEYINPUT75), .B(n302), .ZN(n303) );
  XNOR2_X1 U346 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n331) );
  XOR2_X1 U348 ( .A(G36GAT), .B(G190GAT), .Z(n352) );
  XOR2_X1 U349 ( .A(n331), .B(n352), .Z(n306) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(G85GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n305), .B(KEYINPUT72), .ZN(n374) );
  XNOR2_X1 U352 ( .A(n361), .B(n309), .ZN(n554) );
  XOR2_X1 U353 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n311) );
  XNOR2_X1 U354 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT87), .B(n312), .Z(n353) );
  XOR2_X1 U357 ( .A(KEYINPUT0), .B(G134GAT), .Z(n314) );
  XNOR2_X1 U358 ( .A(KEYINPUT83), .B(G127GAT), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U360 ( .A(G113GAT), .B(n315), .Z(n435) );
  XNOR2_X1 U361 ( .A(n353), .B(n435), .ZN(n328) );
  XOR2_X1 U362 ( .A(KEYINPUT86), .B(G99GAT), .Z(n317) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U365 ( .A(G176GAT), .B(KEYINPUT20), .Z(n319) );
  XNOR2_X1 U366 ( .A(KEYINPUT85), .B(KEYINPUT84), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U368 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U369 ( .A(G120GAT), .B(G71GAT), .Z(n384) );
  XOR2_X1 U370 ( .A(G15GAT), .B(n384), .Z(n323) );
  NAND2_X1 U371 ( .A1(G227GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U373 ( .A(G169GAT), .B(n324), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U375 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n330) );
  XNOR2_X1 U376 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n329) );
  XNOR2_X1 U377 ( .A(n330), .B(n329), .ZN(n335) );
  XOR2_X1 U378 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n333) );
  XOR2_X1 U379 ( .A(G141GAT), .B(G22GAT), .Z(n365) );
  XNOR2_X1 U380 ( .A(n365), .B(n331), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U382 ( .A(n335), .B(n334), .Z(n337) );
  NAND2_X1 U383 ( .A1(G228GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U384 ( .A(n337), .B(n336), .ZN(n340) );
  XOR2_X1 U385 ( .A(G155GAT), .B(KEYINPUT2), .Z(n339) );
  XNOR2_X1 U386 ( .A(KEYINPUT3), .B(KEYINPUT90), .ZN(n338) );
  XNOR2_X1 U387 ( .A(n339), .B(n338), .ZN(n438) );
  XOR2_X1 U388 ( .A(n340), .B(n438), .Z(n347) );
  XNOR2_X1 U389 ( .A(G211GAT), .B(G218GAT), .ZN(n341) );
  XNOR2_X1 U390 ( .A(n341), .B(KEYINPUT89), .ZN(n342) );
  XOR2_X1 U391 ( .A(n342), .B(KEYINPUT21), .Z(n344) );
  XNOR2_X1 U392 ( .A(G197GAT), .B(G204GAT), .ZN(n343) );
  XNOR2_X1 U393 ( .A(n344), .B(n343), .ZN(n351) );
  XNOR2_X1 U394 ( .A(G106GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U395 ( .A(n345), .B(G148GAT), .ZN(n375) );
  XNOR2_X1 U396 ( .A(n351), .B(n375), .ZN(n346) );
  XNOR2_X1 U397 ( .A(n347), .B(n346), .ZN(n456) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(G92GAT), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n348), .B(G64GAT), .ZN(n380) );
  XOR2_X1 U400 ( .A(KEYINPUT95), .B(n380), .Z(n350) );
  NAND2_X1 U401 ( .A1(G226GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n357) );
  XOR2_X1 U403 ( .A(n352), .B(n351), .Z(n355) );
  XOR2_X1 U404 ( .A(G169GAT), .B(G8GAT), .Z(n362) );
  XNOR2_X1 U405 ( .A(n362), .B(n353), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U407 ( .A(n357), .B(n356), .Z(n520) );
  XOR2_X1 U408 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n359) );
  XNOR2_X1 U409 ( .A(G113GAT), .B(G197GAT), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n361), .B(n360), .ZN(n373) );
  XOR2_X1 U412 ( .A(G50GAT), .B(G36GAT), .Z(n364) );
  XOR2_X1 U413 ( .A(G15GAT), .B(G1GAT), .Z(n406) );
  XNOR2_X1 U414 ( .A(n362), .B(n406), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n366) );
  XOR2_X1 U416 ( .A(n366), .B(n365), .Z(n371) );
  XOR2_X1 U417 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n368) );
  NAND2_X1 U418 ( .A1(G229GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U420 ( .A(KEYINPUT67), .B(n369), .ZN(n370) );
  XNOR2_X1 U421 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U422 ( .A(n373), .B(n372), .ZN(n567) );
  XNOR2_X1 U423 ( .A(n375), .B(n374), .ZN(n388) );
  XOR2_X1 U424 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n377) );
  NAND2_X1 U425 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U426 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U427 ( .A(n378), .B(KEYINPUT73), .Z(n382) );
  XNOR2_X1 U428 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n379) );
  XNOR2_X1 U429 ( .A(n379), .B(KEYINPUT71), .ZN(n405) );
  XNOR2_X1 U430 ( .A(n380), .B(n405), .ZN(n381) );
  XNOR2_X1 U431 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U432 ( .A(n383), .B(KEYINPUT32), .Z(n386) );
  XNOR2_X1 U433 ( .A(n384), .B(G204GAT), .ZN(n385) );
  XNOR2_X1 U434 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U435 ( .A(n388), .B(n387), .ZN(n572) );
  XOR2_X1 U436 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n389) );
  XNOR2_X1 U437 ( .A(n572), .B(n389), .ZN(n560) );
  NAND2_X1 U438 ( .A1(n567), .A2(n560), .ZN(n391) );
  XNOR2_X1 U439 ( .A(KEYINPUT114), .B(KEYINPUT46), .ZN(n390) );
  XNOR2_X1 U440 ( .A(n391), .B(n390), .ZN(n413) );
  XOR2_X1 U441 ( .A(G155GAT), .B(G78GAT), .Z(n393) );
  XNOR2_X1 U442 ( .A(G127GAT), .B(G211GAT), .ZN(n392) );
  XNOR2_X1 U443 ( .A(n393), .B(n392), .ZN(n397) );
  XOR2_X1 U444 ( .A(KEYINPUT81), .B(G64GAT), .Z(n395) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(G8GAT), .ZN(n394) );
  XNOR2_X1 U446 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U447 ( .A(n397), .B(n396), .Z(n402) );
  XOR2_X1 U448 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n399) );
  NAND2_X1 U449 ( .A1(G231GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U451 ( .A(KEYINPUT12), .B(n400), .ZN(n401) );
  XNOR2_X1 U452 ( .A(n402), .B(n401), .ZN(n412) );
  XOR2_X1 U453 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n404) );
  XNOR2_X1 U454 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n403) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n410) );
  XOR2_X1 U456 ( .A(n405), .B(G71GAT), .Z(n408) );
  XNOR2_X1 U457 ( .A(n406), .B(G183GAT), .ZN(n407) );
  XNOR2_X1 U458 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U459 ( .A(n410), .B(n409), .Z(n411) );
  XNOR2_X1 U460 ( .A(n412), .B(n411), .ZN(n486) );
  NAND2_X1 U461 ( .A1(n413), .A2(n486), .ZN(n414) );
  NOR2_X1 U462 ( .A1(n554), .A2(n414), .ZN(n415) );
  XOR2_X1 U463 ( .A(KEYINPUT47), .B(n415), .Z(n423) );
  INV_X1 U464 ( .A(n554), .ZN(n467) );
  XNOR2_X1 U465 ( .A(n467), .B(KEYINPUT36), .ZN(n581) );
  NOR2_X1 U466 ( .A1(n581), .A2(n486), .ZN(n417) );
  NOR2_X1 U467 ( .A1(n572), .A2(n418), .ZN(n419) );
  XNOR2_X1 U468 ( .A(n419), .B(KEYINPUT115), .ZN(n420) );
  NOR2_X1 U469 ( .A1(n567), .A2(n420), .ZN(n421) );
  XNOR2_X1 U470 ( .A(KEYINPUT116), .B(n421), .ZN(n422) );
  NOR2_X1 U471 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U472 ( .A(KEYINPUT48), .B(n424), .ZN(n528) );
  NOR2_X1 U473 ( .A1(n520), .A2(n528), .ZN(n425) );
  XNOR2_X1 U474 ( .A(n425), .B(KEYINPUT54), .ZN(n444) );
  XOR2_X1 U475 ( .A(G162GAT), .B(G148GAT), .Z(n427) );
  XNOR2_X1 U476 ( .A(G141GAT), .B(G120GAT), .ZN(n426) );
  XNOR2_X1 U477 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U478 ( .A(KEYINPUT94), .B(KEYINPUT6), .Z(n429) );
  XNOR2_X1 U479 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n428) );
  XNOR2_X1 U480 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U481 ( .A(n431), .B(n430), .Z(n437) );
  XOR2_X1 U482 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n433) );
  XNOR2_X1 U483 ( .A(KEYINPUT1), .B(G57GAT), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U486 ( .A(n437), .B(n436), .ZN(n443) );
  XOR2_X1 U487 ( .A(G85GAT), .B(n438), .Z(n440) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U489 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U490 ( .A(G29GAT), .B(n441), .Z(n442) );
  XNOR2_X1 U491 ( .A(n443), .B(n442), .ZN(n518) );
  NAND2_X1 U492 ( .A1(n444), .A2(n518), .ZN(n565) );
  NOR2_X1 U493 ( .A1(n456), .A2(n565), .ZN(n446) );
  XNOR2_X1 U494 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n445) );
  XNOR2_X1 U495 ( .A(n446), .B(n445), .ZN(n447) );
  NAND2_X1 U496 ( .A1(n554), .A2(n563), .ZN(n449) );
  XOR2_X1 U497 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n475) );
  XNOR2_X1 U498 ( .A(n456), .B(KEYINPUT66), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n450), .B(KEYINPUT28), .ZN(n535) );
  INV_X1 U500 ( .A(n518), .ZN(n473) );
  XOR2_X1 U501 ( .A(n520), .B(KEYINPUT27), .Z(n460) );
  NAND2_X1 U502 ( .A1(n473), .A2(n460), .ZN(n529) );
  NOR2_X1 U503 ( .A1(n535), .A2(n529), .ZN(n451) );
  NAND2_X1 U504 ( .A1(n531), .A2(n451), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n452), .B(KEYINPUT96), .ZN(n466) );
  NOR2_X1 U506 ( .A1(n531), .A2(n520), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n453), .B(KEYINPUT98), .ZN(n454) );
  NOR2_X1 U508 ( .A1(n456), .A2(n454), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n455), .B(KEYINPUT25), .ZN(n462) );
  XOR2_X1 U510 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n458) );
  NAND2_X1 U511 ( .A1(n456), .A2(n531), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n566) );
  INV_X1 U513 ( .A(n566), .ZN(n459) );
  NAND2_X1 U514 ( .A1(n460), .A2(n459), .ZN(n461) );
  NAND2_X1 U515 ( .A1(n462), .A2(n461), .ZN(n463) );
  XOR2_X1 U516 ( .A(KEYINPUT99), .B(n463), .Z(n464) );
  NAND2_X1 U517 ( .A1(n464), .A2(n518), .ZN(n465) );
  NAND2_X1 U518 ( .A1(n466), .A2(n465), .ZN(n485) );
  XOR2_X1 U519 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n469) );
  INV_X1 U520 ( .A(n486), .ZN(n575) );
  NAND2_X1 U521 ( .A1(n575), .A2(n467), .ZN(n468) );
  XNOR2_X1 U522 ( .A(n469), .B(n468), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n485), .A2(n470), .ZN(n471) );
  XOR2_X1 U524 ( .A(KEYINPUT100), .B(n471), .Z(n503) );
  INV_X1 U525 ( .A(n567), .ZN(n501) );
  NOR2_X1 U526 ( .A1(n572), .A2(n501), .ZN(n489) );
  NAND2_X1 U527 ( .A1(n503), .A2(n489), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT101), .ZN(n482) );
  NAND2_X1 U529 ( .A1(n482), .A2(n473), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U531 ( .A(G1GAT), .B(n476), .Z(G1324GAT) );
  INV_X1 U532 ( .A(n520), .ZN(n477) );
  NAND2_X1 U533 ( .A1(n477), .A2(n482), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT35), .Z(n481) );
  INV_X1 U536 ( .A(n531), .ZN(n479) );
  NAND2_X1 U537 ( .A1(n482), .A2(n479), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  XOR2_X1 U539 ( .A(G22GAT), .B(KEYINPUT103), .Z(n484) );
  NAND2_X1 U540 ( .A1(n482), .A2(n535), .ZN(n483) );
  XNOR2_X1 U541 ( .A(n484), .B(n483), .ZN(G1327GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT38), .B(KEYINPUT105), .Z(n491) );
  NAND2_X1 U543 ( .A1(n486), .A2(n485), .ZN(n487) );
  NOR2_X1 U544 ( .A1(n581), .A2(n487), .ZN(n488) );
  XOR2_X1 U545 ( .A(KEYINPUT37), .B(n488), .Z(n517) );
  NAND2_X1 U546 ( .A1(n517), .A2(n489), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n491), .B(n490), .ZN(n499) );
  NOR2_X1 U548 ( .A1(n499), .A2(n518), .ZN(n493) );
  XNOR2_X1 U549 ( .A(KEYINPUT104), .B(KEYINPUT39), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U551 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n520), .A2(n499), .ZN(n495) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  XNOR2_X1 U554 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n497) );
  NOR2_X1 U555 ( .A1(n531), .A2(n499), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U557 ( .A(G43GAT), .B(n498), .Z(G1330GAT) );
  INV_X1 U558 ( .A(n535), .ZN(n524) );
  NOR2_X1 U559 ( .A1(n499), .A2(n524), .ZN(n500) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n500), .Z(G1331GAT) );
  NAND2_X1 U561 ( .A1(n560), .A2(n501), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(KEYINPUT107), .ZN(n516) );
  NAND2_X1 U563 ( .A1(n516), .A2(n503), .ZN(n512) );
  NOR2_X1 U564 ( .A1(n518), .A2(n512), .ZN(n506) );
  XOR2_X1 U565 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n504) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n520), .A2(n512), .ZN(n508) );
  XNOR2_X1 U569 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n509), .ZN(G1333GAT) );
  NOR2_X1 U572 ( .A1(n531), .A2(n512), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(KEYINPUT111), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1334GAT) );
  NOR2_X1 U575 ( .A1(n524), .A2(n512), .ZN(n514) );
  XNOR2_X1 U576 ( .A(KEYINPUT43), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n515), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n518), .A2(n523), .ZN(n519) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n520), .A2(n523), .ZN(n521) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U584 ( .A1(n531), .A2(n523), .ZN(n522) );
  XOR2_X1 U585 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X1 U587 ( .A(KEYINPUT113), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  INV_X1 U590 ( .A(KEYINPUT118), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U592 ( .A(n530), .B(KEYINPUT117), .ZN(n546) );
  NOR2_X1 U593 ( .A1(n531), .A2(n546), .ZN(n532) );
  XNOR2_X1 U594 ( .A(n533), .B(n532), .ZN(n534) );
  NOR2_X1 U595 ( .A1(n535), .A2(n534), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n542), .A2(n567), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U599 ( .A1(n542), .A2(n560), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n540) );
  NAND2_X1 U602 ( .A1(n542), .A2(n575), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U606 ( .A1(n542), .A2(n554), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U609 ( .A1(n566), .A2(n546), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n567), .A2(n553), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U613 ( .A1(n553), .A2(n560), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n550), .ZN(G1345GAT) );
  XOR2_X1 U616 ( .A(G155GAT), .B(KEYINPUT121), .Z(n552) );
  NAND2_X1 U617 ( .A1(n553), .A2(n575), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1346GAT) );
  NAND2_X1 U619 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n567), .A2(n563), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT56), .B(n559), .Z(n562) );
  NAND2_X1 U627 ( .A1(n563), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n575), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT125), .Z(n569) );
  NOR2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n579) );
  NAND2_X1 U633 ( .A1(n579), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n578) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n583) );
  INV_X1 U645 ( .A(n579), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(n583), .B(n582), .Z(G1355GAT) );
endmodule

