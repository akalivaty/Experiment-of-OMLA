//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G68), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n213), .A2(new_n214), .B1(new_n202), .B2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n212), .B(new_n216), .C1(G107), .C2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  AND2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(G58), .A2(G232), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(G58), .A2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n209), .B(new_n227), .C1(new_n230), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G264), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n238), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G97), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G107), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n247), .B(new_n252), .ZN(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT64), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G41), .B2(G45), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n256), .B1(new_n255), .B2(new_n258), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G226), .ZN(new_n262));
  INV_X1    g0062(.A(G274), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(KEYINPUT65), .A3(new_n228), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT65), .ZN(new_n267));
  AND2_X1   g0067(.A1(G1), .A2(G13), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n254), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G222), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G223), .A2(G1698), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n270), .B(new_n275), .C1(G77), .C2(new_n271), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n262), .A2(new_n264), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G200), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n229), .B1(new_n231), .B2(new_n220), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(G150), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT66), .A2(G58), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT66), .A2(G58), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT8), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n286), .B1(KEYINPUT8), .B2(G58), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n229), .A2(G33), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(new_n228), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n257), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n289), .A2(new_n291), .B1(new_n220), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n291), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n257), .A2(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT9), .ZN(new_n301));
  OAI221_X1 g0101(.A(new_n278), .B1(new_n279), .B2(new_n277), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n301), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT10), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n277), .A2(new_n279), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n294), .A2(new_n299), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(KEYINPUT9), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT10), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(new_n303), .A4(new_n278), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n277), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n300), .B(new_n313), .C1(G179), .C2(new_n277), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n316), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n317));
  XOR2_X1   g0117(.A(KEYINPUT15), .B(G87), .Z(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n288), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n291), .B1(new_n222), .B2(new_n293), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n298), .A2(G77), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n261), .A2(G244), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G238), .A2(G1698), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n271), .B(new_n325), .C1(new_n240), .C2(G1698), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n270), .B(new_n326), .C1(G107), .C2(new_n271), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n324), .A2(new_n264), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT67), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n329), .A3(G190), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n324), .A2(new_n264), .A3(new_n327), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT67), .B1(new_n331), .B2(new_n279), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n323), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n331), .A2(G200), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n311), .A2(new_n314), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n271), .B2(G20), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT70), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT3), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  INV_X1    g0141(.A(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n343));
  OAI211_X1 g0143(.A(KEYINPUT7), .B(new_n229), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(G33), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n348), .A2(KEYINPUT70), .A3(KEYINPUT7), .A4(new_n229), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(G68), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT66), .B(G58), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n232), .B1(new_n351), .B2(new_n210), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(G20), .B1(G159), .B2(new_n281), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n231), .B1(new_n285), .B2(G68), .ZN(new_n357));
  INV_X1    g0157(.A(G159), .ZN(new_n358));
  INV_X1    g0158(.A(new_n281), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n357), .A2(new_n229), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n210), .B1(new_n338), .B2(new_n344), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n295), .B1(new_n362), .B2(KEYINPUT16), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n255), .A2(new_n258), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n264), .B1(new_n365), .B2(new_n240), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(G223), .A2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n221), .A2(G1698), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n346), .A2(new_n368), .A3(new_n347), .A4(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n342), .B2(new_n213), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n270), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G200), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n371), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT71), .B1(new_n371), .B2(new_n270), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n367), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n375), .B1(new_n378), .B2(G190), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n287), .A2(new_n292), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n287), .B2(new_n298), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n364), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n381), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n356), .B2(new_n363), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n379), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n338), .A2(new_n344), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n390), .A2(new_n353), .A3(KEYINPUT16), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n291), .ZN(new_n392));
  AOI21_X1  g0192(.A(KEYINPUT16), .B1(new_n350), .B2(new_n353), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n381), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n366), .B1(new_n270), .B2(new_n371), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(G169), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT71), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n372), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n371), .A2(KEYINPUT71), .A3(new_n270), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n366), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G179), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n396), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n394), .A2(new_n402), .A3(KEYINPUT18), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT18), .B1(new_n394), .B2(new_n402), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n328), .A2(new_n401), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n331), .A2(new_n312), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n323), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n388), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G238), .B1(new_n259), .B2(new_n260), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G97), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n240), .A2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G226), .B2(G1698), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n412), .B1(new_n414), .B2(new_n348), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n270), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n411), .A2(new_n416), .A3(new_n264), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT68), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT13), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n411), .A2(new_n416), .A3(new_n420), .A4(new_n264), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(KEYINPUT68), .A3(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(G169), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT14), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n422), .A2(new_n426), .A3(G169), .A4(new_n423), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n418), .A2(G179), .A3(new_n421), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n425), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n359), .A2(new_n220), .B1(new_n229), .B2(G68), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n288), .A2(new_n222), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n291), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g0232(.A(new_n432), .B(KEYINPUT11), .Z(new_n433));
  INV_X1    g0233(.A(KEYINPUT12), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n293), .B2(new_n210), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n292), .A2(KEYINPUT12), .A3(G68), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n435), .A2(new_n436), .B1(new_n297), .B2(new_n210), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n429), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT69), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n422), .A2(G200), .A3(new_n423), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n418), .A2(G190), .A3(new_n421), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(new_n438), .A3(new_n443), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n441), .B1(new_n440), .B2(new_n444), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n336), .B(new_n410), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n271), .B1(G257), .B2(new_n272), .ZN(new_n448));
  NOR2_X1   g0248(.A1(G250), .A2(G1698), .ZN(new_n449));
  INV_X1    g0249(.A(G294), .ZN(new_n450));
  OAI22_X1  g0250(.A1(new_n448), .A2(new_n449), .B1(new_n342), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n270), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT75), .ZN(new_n453));
  INV_X1    g0253(.A(G41), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT5), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(KEYINPUT75), .B2(G41), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(new_n460), .A2(new_n255), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G264), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n455), .A2(new_n457), .A3(new_n459), .A4(G274), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G169), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n451), .A2(new_n270), .B1(G264), .B2(new_n461), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(G179), .A3(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n257), .A2(G33), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n292), .A2(new_n470), .A3(new_n228), .A4(new_n290), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n473), .A2(new_n474), .A3(new_n203), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n346), .A2(new_n347), .A3(new_n229), .A4(G87), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT22), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n271), .A2(new_n478), .A3(new_n229), .A4(G87), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT80), .B1(new_n229), .B2(G107), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n484));
  OAI211_X1 g0284(.A(KEYINPUT80), .B(KEYINPUT23), .C1(new_n229), .C2(G107), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT24), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT24), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n480), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n475), .B1(new_n491), .B2(new_n291), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n292), .A2(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT25), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n469), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n480), .A2(new_n489), .A3(new_n486), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n489), .B1(new_n480), .B2(new_n486), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n291), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n475), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n469), .A3(new_n499), .A4(new_n494), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n468), .B1(new_n495), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n498), .A2(new_n499), .A3(new_n494), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n374), .B1(new_n466), .B2(new_n463), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n464), .A2(new_n279), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n293), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g0309(.A1(new_n471), .A2(new_n508), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(new_n229), .C1(G33), .C2(new_n202), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n291), .C1(new_n229), .C2(G116), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT20), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n509), .B(new_n510), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G264), .A2(G1698), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n271), .B(new_n519), .C1(new_n215), .C2(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n270), .B(new_n520), .C1(G303), .C2(new_n271), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n461), .A2(G270), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n522), .A3(new_n463), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G200), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n518), .B(new_n524), .C1(new_n279), .C2(new_n523), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n517), .A2(G169), .A3(new_n523), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n523), .A2(new_n401), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n517), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n517), .A2(new_n523), .A3(KEYINPUT21), .A4(G169), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n525), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n502), .A2(new_n507), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n345), .A2(G107), .A3(new_n349), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT6), .ZN(new_n538));
  INV_X1    g0338(.A(new_n204), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n202), .A2(new_n203), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n538), .B2(new_n248), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(G20), .B1(G77), .B2(new_n281), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n345), .A2(KEYINPUT72), .A3(G107), .A4(new_n349), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n291), .ZN(new_n546));
  OAI21_X1  g0346(.A(G97), .B1(new_n473), .B2(new_n474), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n547), .B(KEYINPUT74), .C1(G97), .C2(new_n293), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT74), .ZN(new_n549));
  OR2_X1    g0349(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n202), .B1(new_n550), .B2(new_n472), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n293), .A2(G97), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n546), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n346), .A2(new_n347), .A3(G244), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT4), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n557), .A2(G1698), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n271), .A2(G244), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n560), .A3(new_n511), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n271), .A2(G250), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n272), .B1(new_n562), .B2(KEYINPUT4), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n270), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n460), .A2(G257), .A3(new_n255), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n463), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT76), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(KEYINPUT76), .A3(new_n463), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n312), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n564), .A2(new_n568), .A3(new_n401), .A4(new_n569), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n555), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT79), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n271), .A2(new_n229), .A3(G68), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n288), .B2(new_n202), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n412), .A2(new_n577), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(G20), .ZN(new_n580));
  OR2_X1    g0380(.A1(KEYINPUT77), .A2(G87), .ZN(new_n581));
  NAND2_X1  g0381(.A1(KEYINPUT77), .A2(G87), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n204), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n576), .B(new_n578), .C1(new_n580), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n291), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n550), .A2(new_n318), .A3(new_n472), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n319), .A2(new_n293), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n211), .A2(new_n272), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n223), .A2(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n346), .A2(new_n589), .A3(new_n347), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(G33), .A2(G116), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n270), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n214), .B1(new_n458), .B2(G1), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n257), .A2(new_n263), .A3(G45), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n255), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n312), .ZN(new_n599));
  INV_X1    g0399(.A(new_n597), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n593), .B2(new_n270), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n401), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n588), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT65), .B1(new_n265), .B2(new_n228), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n268), .A2(new_n267), .A3(new_n254), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n592), .B2(new_n591), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT78), .ZN(new_n608));
  NOR4_X1   g0408(.A1(new_n607), .A2(new_n608), .A3(new_n279), .A4(new_n600), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT78), .B1(new_n598), .B2(G200), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n594), .A2(G190), .A3(new_n597), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n550), .A2(G87), .A3(new_n472), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n585), .A2(new_n613), .A3(new_n587), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n575), .B(new_n603), .C1(new_n612), .C2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n611), .B(new_n608), .C1(new_n374), .C2(new_n601), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n601), .A2(KEYINPUT78), .A3(G190), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n588), .A2(new_n599), .A3(new_n602), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT79), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n570), .A2(G200), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n564), .A2(new_n568), .A3(G190), .A4(new_n569), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n546), .A2(new_n554), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n574), .A2(new_n615), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n447), .A2(new_n534), .A3(new_n624), .ZN(G372));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n403), .A2(new_n404), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT18), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n378), .A2(G179), .B1(G169), .B2(new_n395), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n628), .B1(new_n386), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n394), .A2(new_n402), .A3(KEYINPUT18), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT87), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n627), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n444), .A2(new_n409), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n388), .B1(new_n440), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n311), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n314), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT82), .B1(new_n601), .B2(G169), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT82), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n641), .B(new_n312), .C1(new_n607), .C2(new_n600), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n640), .A2(new_n642), .A3(new_n602), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT83), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n640), .A2(new_n642), .A3(KEYINPUT83), .A4(new_n602), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n588), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n546), .A2(new_n554), .A3(new_n621), .A4(new_n622), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n545), .A2(new_n291), .B1(new_n553), .B2(new_n548), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n571), .A2(new_n572), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n468), .A2(new_n503), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n612), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n614), .A2(KEYINPUT84), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT84), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n584), .A2(new_n291), .B1(new_n293), .B2(new_n319), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n613), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n647), .A2(new_n588), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n653), .A2(new_n507), .A3(new_n656), .A4(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n555), .A2(KEYINPUT85), .A3(new_n573), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT85), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n650), .B2(new_n651), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT26), .B1(new_n668), .B2(new_n663), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n620), .A2(new_n615), .ZN(new_n670));
  XNOR2_X1  g0470(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n670), .A2(new_n574), .A3(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n648), .B(new_n664), .C1(new_n669), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n639), .B1(new_n447), .B2(new_n674), .ZN(G369));
  INV_X1    g0475(.A(new_n468), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n503), .A2(KEYINPUT81), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n676), .B1(new_n677), .B2(new_n500), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n506), .ZN(new_n679));
  INV_X1    g0479(.A(G13), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G20), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n257), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(KEYINPUT27), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(G213), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT88), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G343), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n495), .B2(new_n501), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n679), .A2(new_n689), .B1(new_n678), .B2(new_n688), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n654), .B2(new_n688), .ZN(new_n691));
  INV_X1    g0491(.A(G330), .ZN(new_n692));
  OR3_X1    g0492(.A1(new_n654), .A2(new_n518), .A3(new_n687), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n533), .B1(new_n518), .B2(new_n687), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n654), .A2(new_n688), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n679), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n468), .A2(new_n503), .A3(new_n687), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  NAND2_X1  g0502(.A1(new_n583), .A2(new_n508), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n207), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(G1), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n233), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT85), .B1(new_n555), .B2(new_n573), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n650), .A2(new_n651), .A3(new_n666), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT26), .B(new_n663), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT90), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n671), .B1(new_n670), .B2(new_n574), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT90), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n668), .A2(new_n716), .A3(KEYINPUT26), .A4(new_n663), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n648), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n507), .A2(new_n663), .A3(new_n574), .A4(new_n623), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n502), .A2(new_n654), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .A3(new_n687), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n673), .A2(new_n687), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n564), .A2(new_n568), .A3(new_n569), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(new_n529), .A3(new_n466), .A4(new_n601), .ZN(new_n730));
  NOR2_X1   g0530(.A1(KEYINPUT89), .A2(KEYINPUT30), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n730), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n570), .A2(new_n464), .A3(new_n401), .A4(new_n523), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n601), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n687), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n534), .A2(new_n624), .A3(new_n688), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT31), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n730), .B(new_n731), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT31), .B(new_n688), .C1(new_n742), .C2(new_n735), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G330), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n728), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n710), .B1(new_n747), .B2(G1), .ZN(G364));
  INV_X1    g0548(.A(KEYINPUT91), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n695), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n681), .A2(G45), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n707), .A2(G1), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n693), .A2(new_n694), .A3(new_n692), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n750), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n228), .B1(G20), .B2(new_n312), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n374), .A2(G179), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n229), .A2(G190), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n203), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT93), .ZN(new_n762));
  INV_X1    g0562(.A(new_n758), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G159), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT32), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n401), .A2(new_n374), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n758), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n760), .B(new_n766), .C1(G68), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(G20), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n401), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n758), .A2(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n773), .A2(new_n220), .B1(new_n775), .B2(new_n222), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n772), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n776), .B1(new_n285), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT92), .ZN(new_n780));
  OAI21_X1  g0580(.A(G20), .B1(new_n762), .B2(new_n279), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G97), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n757), .A2(new_n772), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n581), .A3(new_n582), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n770), .A2(new_n271), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n759), .A2(new_n788), .B1(new_n777), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT33), .B(G317), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(new_n769), .B2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G326), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n793), .B2(new_n773), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n271), .B1(new_n764), .B2(G329), .ZN(new_n795));
  INV_X1    g0595(.A(new_n781), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n450), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n775), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n794), .B(new_n797), .C1(G311), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G303), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n784), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n756), .B1(new_n787), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n693), .A2(new_n694), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n234), .A2(new_n458), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n705), .A2(new_n271), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n807), .B(new_n808), .C1(new_n247), .C2(new_n458), .ZN(new_n809));
  INV_X1    g0609(.A(G355), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n271), .A2(new_n207), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(G116), .B2(new_n207), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n805), .A2(new_n755), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n752), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n806), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n754), .B1(new_n802), .B2(new_n816), .ZN(G396));
  AOI21_X1  g0617(.A(new_n348), .B1(new_n781), .B2(new_n285), .ZN(new_n818));
  INV_X1    g0618(.A(G132), .ZN(new_n819));
  INV_X1    g0619(.A(new_n764), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n220), .B2(new_n784), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G150), .A2(new_n769), .B1(new_n778), .B2(G143), .ZN(new_n822));
  INV_X1    g0622(.A(new_n773), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G137), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n358), .C2(new_n775), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT34), .Z(new_n826));
  INV_X1    g0626(.A(new_n759), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n821), .B(new_n826), .C1(G68), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G311), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n782), .B1(new_n450), .B2(new_n777), .C1(new_n829), .C2(new_n820), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n271), .B1(new_n769), .B2(G283), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n831), .B1(new_n508), .B2(new_n775), .C1(new_n800), .C2(new_n773), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n759), .A2(new_n213), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n784), .A2(new_n203), .ZN(new_n834));
  NOR4_X1   g0634(.A1(new_n830), .A2(new_n832), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n755), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n755), .A2(new_n803), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n836), .B(new_n815), .C1(G77), .C2(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT94), .Z(new_n840));
  NAND2_X1  g0640(.A1(new_n688), .A2(new_n323), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n409), .B1(new_n335), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n408), .A2(new_n688), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n840), .B1(new_n803), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT95), .Z(new_n847));
  NAND3_X1  g0647(.A1(new_n673), .A2(new_n687), .A3(new_n844), .ZN(new_n848));
  INV_X1    g0648(.A(new_n725), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT96), .ZN(new_n850));
  INV_X1    g0650(.A(new_n843), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n335), .A2(new_n841), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n409), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT96), .B1(new_n842), .B2(new_n843), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n848), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(new_n745), .Z(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n752), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n847), .A2(new_n858), .ZN(G384));
  NOR2_X1   g0659(.A1(new_n438), .A2(new_n687), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n860), .A2(KEYINPUT98), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n861), .A2(new_n444), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n860), .A2(KEYINPUT98), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT97), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n429), .A2(new_n864), .A3(new_n439), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n429), .B2(new_n439), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n862), .B(new_n863), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n429), .A2(new_n439), .A3(new_n688), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n678), .A2(new_n506), .A3(new_n532), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n623), .B1(new_n650), .B2(new_n651), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(new_n670), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n872), .A3(new_n687), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n737), .B1(new_n873), .B2(KEYINPUT31), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n743), .A2(KEYINPUT102), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n733), .A2(new_n736), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT102), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT31), .A4(new_n688), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n869), .B(new_n844), .C1(new_n874), .C2(new_n879), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n384), .A2(new_n387), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n627), .B2(new_n632), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n394), .A2(new_n686), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n394), .A2(new_n402), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n382), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  XOR2_X1   g0687(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n888), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n382), .A2(new_n886), .A3(new_n883), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(KEYINPUT38), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n686), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n391), .A2(new_n895), .A3(new_n291), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n629), .A2(new_n894), .B1(new_n381), .B2(new_n896), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n400), .A2(new_n279), .B1(new_n374), .B2(new_n373), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n394), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n891), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT100), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n896), .A2(new_n381), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n686), .B(new_n904), .C1(new_n388), .C2(new_n405), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n900), .A2(KEYINPUT100), .A3(new_n891), .ZN(new_n906));
  AND4_X1   g0706(.A1(KEYINPUT38), .A2(new_n903), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n893), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT40), .B1(new_n880), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n903), .A2(new_n905), .A3(KEYINPUT38), .A4(new_n906), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT40), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n845), .B1(new_n867), .B2(new_n868), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n875), .A2(new_n878), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n741), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n909), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n447), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(G330), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n919), .B2(new_n922), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT103), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n634), .A2(new_n894), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n848), .A2(new_n851), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n912), .A2(new_n913), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n928), .A3(new_n869), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n882), .A2(new_n884), .B1(new_n891), .B2(new_n889), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n913), .B1(new_n930), .B2(KEYINPUT38), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n932), .B2(new_n928), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n865), .A2(new_n866), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n688), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n926), .B(new_n929), .C1(new_n934), .C2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n925), .B(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n724), .A2(new_n920), .A3(new_n727), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT101), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT29), .B1(new_n673), .B2(new_n687), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n688), .B1(new_n718), .B2(new_n722), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n942), .B1(KEYINPUT29), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT101), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(new_n945), .A3(new_n920), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n638), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n939), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n257), .B2(new_n681), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n508), .B1(new_n542), .B2(KEYINPUT35), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n230), .C1(KEYINPUT35), .C2(new_n542), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n234), .B1(new_n351), .B2(new_n210), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n953), .A2(new_n222), .B1(G50), .B2(new_n210), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n680), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n949), .A2(new_n952), .A3(new_n955), .ZN(G367));
  NAND2_X1  g0756(.A1(new_n751), .A2(G1), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT106), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT45), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT105), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n653), .B1(new_n650), .B2(new_n687), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n652), .A2(new_n688), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n701), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n961), .B1(new_n701), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n967), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n699), .A2(new_n700), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n971), .A2(new_n962), .A3(new_n963), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n968), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n691), .A2(new_n699), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n696), .B1(new_n750), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n728), .A3(new_n745), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n959), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n979), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(KEYINPUT106), .A3(new_n975), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n746), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n706), .B(KEYINPUT41), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n958), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n699), .A2(new_n871), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT42), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n688), .B1(new_n661), .B2(new_n658), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n663), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n648), .A2(new_n989), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n574), .B1(new_n962), .B2(new_n502), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n687), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n988), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT104), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n993), .B1(new_n988), .B2(new_n995), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n992), .A2(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n696), .A2(new_n964), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1001), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n986), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n808), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n813), .B1(new_n207), .B2(new_n319), .C1(new_n238), .C2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n348), .B1(new_n773), .B2(new_n829), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n759), .A2(new_n202), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n784), .A2(new_n508), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1010), .A2(KEYINPUT46), .B1(new_n769), .B2(G294), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(KEYINPUT46), .B2(new_n1010), .C1(new_n800), .C2(new_n777), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1009), .B(new_n1012), .C1(G317), .C2(new_n764), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n203), .B2(new_n796), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1008), .B(new_n1014), .C1(G283), .C2(new_n798), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n764), .A2(G137), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n781), .A2(G68), .B1(G143), .B2(new_n823), .ZN(new_n1017));
  INV_X1    g0817(.A(G150), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n777), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT107), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n271), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1019), .A2(KEYINPUT107), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n827), .A2(G77), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n769), .A2(G159), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n798), .A2(G50), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1021), .B(new_n1026), .C1(new_n285), .C2(new_n785), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1015), .B1(new_n1016), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1028), .B(new_n1029), .Z(new_n1030));
  OAI211_X1 g0830(.A(new_n815), .B(new_n1007), .C1(new_n1030), .C2(new_n756), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n992), .A2(G20), .A3(new_n804), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1005), .A2(new_n1034), .ZN(G387));
  OAI22_X1  g0835(.A1(new_n287), .A2(new_n768), .B1(new_n210), .B2(new_n775), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT111), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1009), .B(new_n1037), .C1(G159), .C2(new_n823), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n778), .A2(G50), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n348), .B1(new_n785), .B2(G77), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(KEYINPUT110), .B(G150), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n781), .A2(new_n318), .B1(new_n764), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(G317), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n775), .A2(new_n800), .B1(new_n777), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT112), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n829), .B2(new_n768), .C1(new_n789), .C2(new_n773), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT48), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n788), .B2(new_n796), .C1(new_n450), .C2(new_n784), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n348), .B1(new_n508), .B2(new_n759), .C1(new_n820), .C2(new_n793), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1043), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n755), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n690), .A2(new_n805), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n815), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n243), .A2(G45), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT109), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n315), .A2(G50), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT50), .ZN(new_n1060));
  AOI21_X1  g0860(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1060), .A2(new_n704), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1058), .A2(new_n808), .A3(new_n1062), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1063), .B1(G107), .B2(new_n207), .C1(new_n704), .C2(new_n811), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1056), .B1(new_n813), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n957), .B2(new_n978), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n706), .B1(new_n747), .B2(new_n978), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1066), .B1(new_n981), .B2(new_n1067), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n980), .A2(new_n982), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT114), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n976), .A2(new_n1070), .A3(new_n696), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n696), .A2(new_n1070), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n697), .A2(KEYINPUT114), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n975), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1069), .B(new_n706), .C1(new_n1075), .C2(new_n981), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n962), .A2(new_n805), .A3(new_n963), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G150), .A2(new_n823), .B1(new_n778), .B2(G159), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n271), .B1(new_n768), .B2(new_n220), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n784), .A2(new_n210), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1081), .A2(new_n833), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n781), .A2(G77), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n798), .A2(new_n316), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1078), .A2(new_n1080), .B1(new_n764), .B2(G143), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n773), .A2(new_n1044), .B1(new_n777), .B2(new_n829), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT52), .Z(new_n1090));
  OAI21_X1  g0890(.A(new_n348), .B1(new_n784), .B2(new_n788), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1090), .A2(new_n760), .A3(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n789), .B2(new_n820), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n781), .A2(G116), .B1(G294), .B2(new_n798), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n800), .B2(new_n768), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT116), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1088), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n755), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n813), .B1(new_n202), .B2(new_n207), .C1(new_n252), .C2(new_n1006), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1077), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1075), .A2(new_n957), .B1(new_n815), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1076), .A2(new_n1101), .ZN(G390));
  INV_X1    g0902(.A(KEYINPUT120), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n922), .A2(G330), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n945), .B1(new_n944), .B2(new_n920), .ZN(new_n1106));
  AND4_X1   g0906(.A1(new_n945), .A2(new_n724), .A3(new_n920), .A4(new_n727), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n639), .B(new_n1105), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n744), .A2(G330), .A3(new_n844), .A4(new_n869), .ZN(new_n1109));
  OAI211_X1 g0909(.A(G330), .B(new_n855), .C1(new_n874), .C2(new_n879), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n869), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n842), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n843), .B1(new_n943), .B2(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1109), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  AND2_X1   g0915(.A1(new_n848), .A2(new_n851), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n743), .ZN(new_n1117));
  OAI211_X1 g0917(.A(G330), .B(new_n844), .C1(new_n874), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1111), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n917), .A2(G330), .A3(new_n915), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1104), .B1(new_n1108), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n937), .B1(new_n1116), .B2(new_n1111), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n934), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n688), .B(new_n842), .C1(new_n718), .C2(new_n722), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n869), .B1(new_n1126), .B2(new_n843), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n908), .A2(new_n936), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1125), .A2(new_n1129), .A3(new_n1109), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1124), .A2(new_n934), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n1120), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1109), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n1116), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1135), .A2(new_n947), .A3(KEYINPUT117), .A4(new_n1105), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1123), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1132), .B1(new_n1123), .B2(new_n1136), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n707), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n785), .A2(new_n1041), .ZN(new_n1140));
  XOR2_X1   g0940(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1141));
  OR2_X1    g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n271), .A3(new_n1143), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n781), .A2(G159), .B1(G137), .B2(new_n769), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n764), .A2(G125), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n819), .C2(new_n777), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  AOI211_X1 g0948(.A(new_n1144), .B(new_n1147), .C1(new_n798), .C2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n823), .A2(G128), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(new_n220), .C2(new_n759), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n759), .A2(new_n210), .B1(new_n777), .B2(new_n508), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n271), .B(new_n1152), .C1(G283), .C2(new_n823), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n764), .A2(G294), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n769), .A2(G107), .ZN(new_n1155));
  AND4_X1   g0955(.A1(new_n1085), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n213), .B2(new_n784), .C1(new_n202), .C2(new_n775), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n815), .B1(new_n1158), .B2(new_n756), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n287), .B2(new_n837), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT119), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n934), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n804), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1132), .B2(new_n958), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1103), .B1(new_n1139), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1123), .A2(new_n1136), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1132), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1123), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n706), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1164), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1170), .A2(KEYINPUT120), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1165), .A2(new_n1172), .ZN(G378));
  INV_X1    g0973(.A(KEYINPUT122), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n307), .A2(new_n894), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n311), .A2(new_n314), .ZN(new_n1177));
  XOR2_X1   g0977(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1176), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n919), .B2(G330), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n692), .B(new_n1185), .C1(new_n909), .C2(new_n918), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n938), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n929), .A2(new_n926), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1162), .B2(new_n936), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n880), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n917), .A2(new_n931), .A3(new_n915), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1192), .A2(new_n914), .B1(new_n1193), .B2(KEYINPUT40), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1185), .B1(new_n1194), .B2(new_n692), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n919), .A2(G330), .A3(new_n1186), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1191), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1174), .B1(new_n1189), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n938), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1195), .A2(new_n1191), .A3(new_n1196), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(KEYINPUT122), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n957), .A3(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(G41), .B(new_n271), .C1(new_n823), .C2(G116), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1203), .B1(new_n203), .B2(new_n777), .C1(new_n796), .C2(new_n210), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n319), .A2(new_n775), .B1(new_n222), .B2(new_n784), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n768), .A2(new_n202), .B1(new_n759), .B2(new_n351), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n788), .B2(new_n820), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT58), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n342), .A2(new_n454), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT121), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n220), .C1(G41), .C2(new_n271), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n781), .A2(G150), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n785), .A2(new_n1148), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G132), .A2(new_n769), .B1(new_n798), .B2(G137), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n823), .A2(G125), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G128), .B2(new_n778), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT59), .Z(new_n1219));
  AOI21_X1  g1019(.A(new_n1211), .B1(new_n764), .B2(G124), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n358), .B2(new_n759), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1209), .B(new_n1212), .C1(new_n1219), .C2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n752), .B1(new_n1222), .B2(new_n755), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(G50), .B2(new_n838), .C1(new_n1185), .C2(new_n804), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1202), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1201), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT122), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1108), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1168), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1189), .A2(new_n1197), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1108), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n706), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1226), .B1(new_n1232), .B2(new_n1237), .ZN(G375));
  NAND2_X1  g1038(.A1(new_n1135), .A2(new_n957), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1111), .A2(new_n803), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n837), .A2(new_n210), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n775), .A2(new_n1018), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n773), .A2(new_n819), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n348), .B(new_n1243), .C1(new_n769), .C2(new_n1148), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n781), .A2(G50), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n764), .A2(G128), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n285), .A2(new_n827), .B1(new_n778), .B2(G137), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1242), .B(new_n1248), .C1(G159), .C2(new_n785), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n781), .A2(new_n318), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n764), .A2(G303), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n769), .A2(G116), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1023), .A4(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n773), .A2(new_n450), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n784), .A2(new_n202), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n348), .B1(new_n777), .B2(new_n788), .C1(new_n203), .C2(new_n775), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n755), .B1(new_n1249), .B2(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1240), .A2(new_n815), .A3(new_n1241), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1239), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1108), .A2(new_n1122), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(KEYINPUT123), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT123), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1108), .A2(new_n1122), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n985), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1166), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1260), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(G381));
  AOI21_X1  g1068(.A(new_n707), .B1(new_n1231), .B2(new_n1234), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1198), .A2(new_n1201), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1233), .B1(new_n1270), .B2(new_n1236), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1225), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1139), .A2(new_n1164), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1033), .B1(new_n986), .B2(new_n1004), .ZN(new_n1275));
  INV_X1    g1075(.A(G390), .ZN(new_n1276));
  INV_X1    g1076(.A(G384), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(G393), .A2(G396), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  OR3_X1    g1079(.A1(new_n1274), .A2(G381), .A3(new_n1279), .ZN(G407));
  INV_X1    g1080(.A(G343), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(G213), .ZN(new_n1282));
  XOR2_X1   g1082(.A(new_n1282), .B(KEYINPUT124), .Z(new_n1283));
  OAI211_X1 g1083(.A(G407), .B(G213), .C1(new_n1274), .C2(new_n1283), .ZN(G409));
  OAI21_X1  g1084(.A(KEYINPUT126), .B1(G387), .B2(new_n1276), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G390), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(G387), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT126), .B1(new_n1076), .B2(new_n1101), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1275), .B2(KEYINPUT125), .ZN(new_n1291));
  XOR2_X1   g1091(.A(G393), .B(G396), .Z(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1285), .A2(new_n1289), .A3(new_n1291), .A4(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(G387), .A2(new_n1276), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1275), .A2(G390), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1292), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1294), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1199), .A2(new_n1200), .A3(new_n957), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1198), .B(new_n1201), .C1(new_n1138), .C2(new_n1108), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1224), .B(new_n1300), .C1(new_n1301), .C2(new_n985), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1273), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1172), .ZN(new_n1304));
  AOI21_X1  g1104(.A(KEYINPUT120), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1303), .B1(new_n1306), .B2(G375), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(new_n1283), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1108), .A2(new_n1122), .A3(KEYINPUT60), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n1136), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n707), .B(new_n1310), .C1(new_n1311), .C2(new_n1312), .ZN(new_n1313));
  NOR3_X1   g1113(.A1(new_n1313), .A2(new_n1277), .A3(new_n1260), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1315), .A2(new_n706), .A3(new_n1309), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1260), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1314), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1314), .A2(new_n1318), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1307), .A2(new_n1282), .A3(new_n1321), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1308), .A2(new_n1320), .B1(new_n1322), .B2(new_n1319), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1282), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(G2897), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1314), .A2(new_n1318), .A3(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(G2897), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1283), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1277), .B1(new_n1313), .B2(new_n1260), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1316), .A2(G384), .A3(new_n1317), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1329), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1327), .A2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1324), .B1(new_n1308), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1299), .B1(new_n1323), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1297), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G378), .A2(new_n1272), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1325), .B1(new_n1338), .B2(new_n1303), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1337), .B1(new_n1339), .B2(new_n1333), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT63), .B1(new_n1339), .B2(new_n1321), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND4_X1  g1142(.A1(new_n1307), .A2(KEYINPUT63), .A3(new_n1283), .A4(new_n1321), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1336), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1298), .A2(new_n1324), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1307), .A2(new_n1282), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1330), .A2(G2897), .A3(new_n1325), .A4(new_n1331), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1347), .B1(new_n1321), .B2(new_n1329), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1345), .B1(new_n1346), .B2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT63), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1322), .A2(new_n1350), .ZN(new_n1351));
  AND4_X1   g1151(.A1(new_n1336), .A2(new_n1349), .A3(new_n1351), .A4(new_n1343), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1335), .B1(new_n1344), .B2(new_n1352), .ZN(G405));
  INV_X1    g1153(.A(new_n1273), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1338), .B1(new_n1354), .B2(new_n1272), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1355), .B(new_n1321), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1299), .ZN(G402));
endmodule


