

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n402, n403, n404, n405,
         n406, n407, n408, n409, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749;

  INV_X1 U373 ( .A(n712), .ZN(n353) );
  INV_X1 U374 ( .A(KEYINPUT56), .ZN(n351) );
  NOR2_X1 U375 ( .A1(n533), .A2(n664), .ZN(n534) );
  OR2_X1 U376 ( .A1(n719), .A2(G902), .ZN(n452) );
  XNOR2_X1 U377 ( .A(n516), .B(n438), .ZN(n409) );
  XNOR2_X1 U378 ( .A(n434), .B(n437), .ZN(n438) );
  XNOR2_X1 U379 ( .A(n411), .B(G101), .ZN(n503) );
  XNOR2_X1 U380 ( .A(n439), .B(G119), .ZN(n436) );
  XNOR2_X1 U381 ( .A(KEYINPUT3), .B(KEYINPUT72), .ZN(n435) );
  XNOR2_X1 U382 ( .A(G107), .B(G116), .ZN(n434) );
  INV_X1 U383 ( .A(KEYINPUT71), .ZN(n439) );
  XNOR2_X1 U384 ( .A(KEYINPUT15), .B(G902), .ZN(n621) );
  XNOR2_X2 U385 ( .A(n350), .B(n525), .ZN(n702) );
  XNOR2_X2 U386 ( .A(n725), .B(n520), .ZN(n350) );
  XNOR2_X1 U387 ( .A(n352), .B(n351), .ZN(G51) );
  NAND2_X1 U388 ( .A1(n408), .A2(n418), .ZN(n352) );
  XNOR2_X2 U389 ( .A(n384), .B(n589), .ZN(n747) );
  NAND2_X2 U390 ( .A1(n747), .A2(n746), .ZN(n432) );
  XNOR2_X1 U391 ( .A(n354), .B(n353), .ZN(G60) );
  NAND2_X1 U392 ( .A1(n407), .A2(n418), .ZN(n354) );
  INV_X1 U393 ( .A(G953), .ZN(n735) );
  XNOR2_X2 U394 ( .A(n383), .B(n382), .ZN(n746) );
  NOR2_X1 U395 ( .A1(n601), .A2(n692), .ZN(n593) );
  XNOR2_X2 U396 ( .A(n535), .B(KEYINPUT1), .ZN(n665) );
  XNOR2_X1 U397 ( .A(n371), .B(n370), .ZN(n744) );
  OR2_X1 U398 ( .A1(n532), .A2(n587), .ZN(n371) );
  XNOR2_X1 U399 ( .A(n571), .B(n556), .ZN(n677) );
  XNOR2_X1 U400 ( .A(n561), .B(KEYINPUT108), .ZN(n679) );
  INV_X1 U401 ( .A(n543), .ZN(n571) );
  XOR2_X2 U402 ( .A(KEYINPUT10), .B(n522), .Z(n733) );
  AND2_X1 U403 ( .A1(n555), .A2(n744), .ZN(n375) );
  INV_X1 U404 ( .A(n562), .ZN(n391) );
  XNOR2_X1 U405 ( .A(n558), .B(KEYINPUT39), .ZN(n572) );
  INV_X1 U406 ( .A(n378), .ZN(n377) );
  NAND2_X1 U407 ( .A1(n649), .A2(n652), .ZN(n680) );
  XNOR2_X1 U408 ( .A(n680), .B(KEYINPUT89), .ZN(n539) );
  XOR2_X1 U409 ( .A(KEYINPUT78), .B(KEYINPUT100), .Z(n509) );
  XNOR2_X1 U410 ( .A(G146), .B(G137), .ZN(n508) );
  XOR2_X1 U411 ( .A(KEYINPUT5), .B(KEYINPUT101), .Z(n507) );
  XNOR2_X1 U412 ( .A(n372), .B(n447), .ZN(n374) );
  INV_X1 U413 ( .A(KEYINPUT48), .ZN(n447) );
  XNOR2_X1 U414 ( .A(n519), .B(n456), .ZN(n511) );
  XNOR2_X1 U415 ( .A(G131), .B(G134), .ZN(n456) );
  XNOR2_X1 U416 ( .A(n477), .B(n412), .ZN(n519) );
  XNOR2_X1 U417 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n412) );
  XOR2_X1 U418 ( .A(G113), .B(G104), .Z(n517) );
  INV_X1 U419 ( .A(KEYINPUT93), .ZN(n431) );
  XNOR2_X1 U420 ( .A(n526), .B(KEYINPUT85), .ZN(n527) );
  XNOR2_X1 U421 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U422 ( .A(n503), .B(n444), .ZN(n521) );
  XNOR2_X1 U423 ( .A(G110), .B(KEYINPUT73), .ZN(n444) );
  XNOR2_X1 U424 ( .A(n521), .B(n441), .ZN(n524) );
  XNOR2_X1 U425 ( .A(n443), .B(n442), .ZN(n441) );
  XNOR2_X1 U426 ( .A(KEYINPUT82), .B(KEYINPUT17), .ZN(n443) );
  NAND2_X1 U427 ( .A1(n735), .A2(G224), .ZN(n442) );
  XNOR2_X1 U428 ( .A(n591), .B(KEYINPUT33), .ZN(n692) );
  NAND2_X1 U429 ( .A1(n388), .A2(n387), .ZN(n386) );
  NOR2_X1 U430 ( .A1(n679), .A2(n392), .ZN(n387) );
  NAND2_X1 U431 ( .A1(n679), .A2(n392), .ZN(n389) );
  NAND2_X1 U432 ( .A1(n681), .A2(n392), .ZN(n390) );
  INV_X1 U433 ( .A(KEYINPUT36), .ZN(n530) );
  NOR2_X1 U434 ( .A1(n446), .A2(n666), .ZN(n445) );
  XNOR2_X1 U435 ( .A(n430), .B(n429), .ZN(n559) );
  XNOR2_X1 U436 ( .A(n472), .B(G475), .ZN(n429) );
  OR2_X1 U437 ( .A1(n710), .A2(G902), .ZN(n430) );
  INV_X1 U438 ( .A(G472), .ZN(n512) );
  OR2_X1 U439 ( .A1(n679), .A2(n582), .ZN(n583) );
  XNOR2_X1 U440 ( .A(n486), .B(n487), .ZN(n719) );
  XNOR2_X1 U441 ( .A(n449), .B(n448), .ZN(n485) );
  NOR2_X1 U442 ( .A1(G953), .A2(G237), .ZN(n505) );
  OR2_X1 U443 ( .A1(G902), .A2(G237), .ZN(n528) );
  INV_X1 U444 ( .A(KEYINPUT67), .ZN(n411) );
  INV_X1 U445 ( .A(G122), .ZN(n437) );
  NAND2_X1 U446 ( .A1(G237), .A2(G234), .ZN(n492) );
  INV_X1 U447 ( .A(n539), .ZN(n609) );
  INV_X1 U448 ( .A(KEYINPUT41), .ZN(n392) );
  NAND2_X1 U449 ( .A1(n677), .A2(n676), .ZN(n681) );
  XNOR2_X1 U450 ( .A(n380), .B(n358), .ZN(n535) );
  OR2_X1 U451 ( .A1(n705), .A2(G902), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n357), .B(n510), .ZN(n394) );
  XNOR2_X1 U453 ( .A(n393), .B(n511), .ZN(n373) );
  XNOR2_X1 U454 ( .A(n450), .B(KEYINPUT23), .ZN(n449) );
  XNOR2_X1 U455 ( .A(KEYINPUT24), .B(G128), .ZN(n450) );
  XNOR2_X1 U456 ( .A(G119), .B(G110), .ZN(n448) );
  XOR2_X1 U457 ( .A(G137), .B(G140), .Z(n483) );
  XOR2_X1 U458 ( .A(KEYINPUT9), .B(G134), .Z(n480) );
  XNOR2_X1 U459 ( .A(n470), .B(n471), .ZN(n710) );
  XNOR2_X1 U460 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U461 ( .A(G131), .B(G122), .Z(n468) );
  XNOR2_X1 U462 ( .A(n511), .B(n483), .ZN(n732) );
  XNOR2_X1 U463 ( .A(G104), .B(G107), .ZN(n460) );
  INV_X1 U464 ( .A(G146), .ZN(n457) );
  INV_X1 U465 ( .A(n654), .ZN(n573) );
  XNOR2_X1 U466 ( .A(n491), .B(n359), .ZN(n451) );
  INV_X1 U467 ( .A(KEYINPUT6), .ZN(n405) );
  NOR2_X1 U468 ( .A1(n415), .A2(n720), .ZN(n414) );
  NOR2_X1 U469 ( .A1(n365), .A2(G472), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n732), .B(n381), .ZN(n705) );
  XNOR2_X1 U471 ( .A(n461), .B(n459), .ZN(n381) );
  XNOR2_X1 U472 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U473 ( .A(n521), .B(n460), .ZN(n461) );
  XNOR2_X1 U474 ( .A(KEYINPUT113), .B(KEYINPUT42), .ZN(n563) );
  XNOR2_X1 U475 ( .A(n403), .B(n402), .ZN(n749) );
  INV_X1 U476 ( .A(KEYINPUT40), .ZN(n402) );
  INV_X1 U477 ( .A(KEYINPUT115), .ZN(n370) );
  INV_X1 U478 ( .A(KEYINPUT35), .ZN(n397) );
  NOR2_X1 U479 ( .A1(n559), .A2(n552), .ZN(n646) );
  NAND2_X1 U480 ( .A1(n361), .A2(n379), .ZN(n378) );
  INV_X1 U481 ( .A(KEYINPUT109), .ZN(n382) );
  NOR2_X1 U482 ( .A1(n590), .A2(n424), .ZN(n423) );
  INV_X1 U483 ( .A(n719), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n378), .B(G143), .ZN(G45) );
  AND2_X1 U485 ( .A1(n390), .A2(n389), .ZN(n355) );
  NAND2_X1 U486 ( .A1(n654), .A2(n433), .ZN(n356) );
  XNOR2_X1 U487 ( .A(n605), .B(n405), .ZN(n613) );
  XOR2_X1 U488 ( .A(n507), .B(n506), .Z(n357) );
  XOR2_X1 U489 ( .A(KEYINPUT70), .B(G469), .Z(n358) );
  XOR2_X1 U490 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n359) );
  XOR2_X1 U491 ( .A(n594), .B(KEYINPUT83), .Z(n360) );
  INV_X1 U492 ( .A(n586), .ZN(n424) );
  AND2_X1 U493 ( .A1(n557), .A2(n594), .ZN(n361) );
  AND2_X1 U494 ( .A1(n386), .A2(n391), .ZN(n362) );
  AND2_X1 U495 ( .A1(n600), .A2(n550), .ZN(n363) );
  OR2_X1 U496 ( .A1(n587), .A2(n424), .ZN(n364) );
  NOR2_X2 U497 ( .A1(n562), .A2(n400), .ZN(n647) );
  XOR2_X1 U498 ( .A(n630), .B(n454), .Z(n365) );
  XOR2_X1 U499 ( .A(n710), .B(n709), .Z(n366) );
  XOR2_X1 U500 ( .A(n702), .B(n701), .Z(n367) );
  AND2_X1 U501 ( .A1(n365), .A2(G472), .ZN(n368) );
  NOR2_X1 U502 ( .A1(G952), .A2(n735), .ZN(n720) );
  INV_X1 U503 ( .A(n720), .ZN(n418) );
  NOR2_X1 U504 ( .A1(n715), .A2(n365), .ZN(n417) );
  NAND2_X1 U505 ( .A1(n715), .A2(n368), .ZN(n416) );
  NAND2_X1 U506 ( .A1(n715), .A2(G217), .ZN(n428) );
  XNOR2_X1 U507 ( .A(n537), .B(KEYINPUT19), .ZN(n369) );
  XNOR2_X1 U508 ( .A(n537), .B(KEYINPUT19), .ZN(n580) );
  INV_X1 U509 ( .A(n571), .ZN(n379) );
  NAND2_X1 U510 ( .A1(n375), .A2(n376), .ZN(n372) );
  XNOR2_X1 U511 ( .A(n373), .B(n394), .ZN(n630) );
  NAND2_X1 U512 ( .A1(n374), .A2(n655), .ZN(n419) );
  XNOR2_X1 U513 ( .A(n565), .B(KEYINPUT46), .ZN(n376) );
  NOR2_X1 U514 ( .A1(n553), .A2(n377), .ZN(n554) );
  NAND2_X1 U515 ( .A1(n611), .A2(n423), .ZN(n383) );
  NAND2_X1 U516 ( .A1(n611), .A2(n385), .ZN(n384) );
  NOR2_X1 U517 ( .A1(n364), .A2(n613), .ZN(n385) );
  XNOR2_X2 U518 ( .A(n585), .B(n584), .ZN(n611) );
  NAND2_X1 U519 ( .A1(n355), .A2(n386), .ZN(n691) );
  NAND2_X1 U520 ( .A1(n362), .A2(n355), .ZN(n564) );
  INV_X1 U521 ( .A(n681), .ZN(n388) );
  XNOR2_X1 U522 ( .A(n516), .B(n504), .ZN(n393) );
  NAND2_X1 U523 ( .A1(n572), .A2(n641), .ZN(n654) );
  NAND2_X1 U524 ( .A1(n395), .A2(n625), .ZN(n626) );
  NAND2_X1 U525 ( .A1(n395), .A2(n735), .ZN(n724) );
  NAND2_X1 U526 ( .A1(n421), .A2(n395), .ZN(n420) );
  NAND2_X1 U527 ( .A1(n734), .A2(n395), .ZN(n657) );
  XNOR2_X2 U528 ( .A(n404), .B(KEYINPUT45), .ZN(n395) );
  NOR2_X2 U529 ( .A1(n396), .A2(n583), .ZN(n585) );
  NOR2_X1 U530 ( .A1(n671), .A2(n396), .ZN(n607) );
  XNOR2_X1 U531 ( .A(n396), .B(n592), .ZN(n601) );
  XNOR2_X2 U532 ( .A(n581), .B(KEYINPUT0), .ZN(n396) );
  XNOR2_X1 U533 ( .A(n745), .B(n596), .ZN(n597) );
  XNOR2_X2 U534 ( .A(n398), .B(n397), .ZN(n745) );
  NAND2_X1 U535 ( .A1(n399), .A2(n360), .ZN(n398) );
  XNOR2_X1 U536 ( .A(n593), .B(KEYINPUT34), .ZN(n399) );
  INV_X1 U537 ( .A(n369), .ZN(n400) );
  XNOR2_X1 U538 ( .A(n419), .B(KEYINPUT92), .ZN(n623) );
  NOR2_X1 U539 ( .A1(n749), .A2(n748), .ZN(n565) );
  NAND2_X1 U540 ( .A1(n620), .A2(n619), .ZN(n404) );
  NAND2_X1 U541 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U542 ( .A1(n572), .A2(n646), .ZN(n403) );
  NAND2_X2 U543 ( .A1(n543), .A2(n676), .ZN(n537) );
  NOR2_X1 U544 ( .A1(n529), .A2(n537), .ZN(n531) );
  XNOR2_X2 U545 ( .A(n513), .B(n512), .ZN(n605) );
  XNOR2_X1 U546 ( .A(n406), .B(n481), .ZN(n714) );
  XNOR2_X1 U547 ( .A(n479), .B(n480), .ZN(n406) );
  NOR2_X1 U548 ( .A1(n623), .A2(n356), .ZN(n421) );
  INV_X1 U549 ( .A(n438), .ZN(n515) );
  XNOR2_X1 U550 ( .A(n711), .B(n366), .ZN(n407) );
  XNOR2_X1 U551 ( .A(n703), .B(n367), .ZN(n408) );
  XNOR2_X2 U552 ( .A(n409), .B(n518), .ZN(n725) );
  AND2_X4 U553 ( .A1(n629), .A2(n628), .ZN(n715) );
  NOR2_X1 U554 ( .A1(n417), .A2(n413), .ZN(n631) );
  NOR2_X1 U555 ( .A1(n617), .A2(n618), .ZN(n619) );
  NAND2_X1 U556 ( .A1(n605), .A2(n676), .ZN(n547) );
  NAND2_X1 U557 ( .A1(n548), .A2(n363), .ZN(n446) );
  XNOR2_X2 U558 ( .A(G128), .B(G143), .ZN(n477) );
  NAND2_X1 U559 ( .A1(n416), .A2(n414), .ZN(n413) );
  XNOR2_X1 U560 ( .A(n420), .B(KEYINPUT90), .ZN(n422) );
  NAND2_X1 U561 ( .A1(n422), .A2(n453), .ZN(n629) );
  XNOR2_X1 U562 ( .A(n425), .B(KEYINPUT125), .ZN(G66) );
  NAND2_X1 U563 ( .A1(n426), .A2(n418), .ZN(n425) );
  XNOR2_X1 U564 ( .A(n428), .B(n427), .ZN(n426) );
  NAND2_X1 U565 ( .A1(n432), .A2(KEYINPUT44), .ZN(n616) );
  XNOR2_X1 U566 ( .A(n432), .B(n431), .ZN(n595) );
  NOR2_X1 U567 ( .A1(n627), .A2(n573), .ZN(n734) );
  INV_X1 U568 ( .A(n621), .ZN(n433) );
  XNOR2_X2 U569 ( .A(n436), .B(n435), .ZN(n516) );
  XNOR2_X2 U570 ( .A(n440), .B(n527), .ZN(n543) );
  NAND2_X1 U571 ( .A1(n702), .A2(n621), .ZN(n440) );
  NAND2_X1 U572 ( .A1(n557), .A2(n677), .ZN(n558) );
  XNOR2_X1 U573 ( .A(n445), .B(n551), .ZN(n557) );
  XNOR2_X2 U574 ( .A(n544), .B(KEYINPUT68), .ZN(n666) );
  XNOR2_X2 U575 ( .A(n452), .B(n451), .ZN(n661) );
  OR2_X1 U576 ( .A1(n656), .A2(n622), .ZN(n453) );
  XNOR2_X1 U577 ( .A(KEYINPUT62), .B(KEYINPUT94), .ZN(n454) );
  AND2_X1 U578 ( .A1(n484), .A2(G221), .ZN(n455) );
  INV_X1 U579 ( .A(n658), .ZN(n628) );
  XNOR2_X1 U580 ( .A(n503), .B(n502), .ZN(n504) );
  INV_X1 U581 ( .A(KEYINPUT44), .ZN(n596) );
  INV_X1 U582 ( .A(n519), .ZN(n520) );
  INV_X1 U583 ( .A(KEYINPUT25), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n567), .B(KEYINPUT114), .ZN(n529) );
  INV_X1 U585 ( .A(KEYINPUT79), .ZN(n551) );
  XNOR2_X1 U586 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U587 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U588 ( .A(n564), .B(n563), .ZN(n748) );
  NAND2_X1 U589 ( .A1(G227), .A2(n735), .ZN(n458) );
  XOR2_X1 U590 ( .A(n665), .B(KEYINPUT95), .Z(n587) );
  XOR2_X2 U591 ( .A(G125), .B(G146), .Z(n522) );
  XNOR2_X1 U592 ( .A(n733), .B(n517), .ZN(n471) );
  XOR2_X1 U593 ( .A(KEYINPUT12), .B(KEYINPUT105), .Z(n463) );
  XNOR2_X1 U594 ( .A(G140), .B(G143), .ZN(n462) );
  XNOR2_X1 U595 ( .A(n463), .B(n462), .ZN(n467) );
  XOR2_X1 U596 ( .A(KEYINPUT104), .B(KEYINPUT11), .Z(n465) );
  NAND2_X1 U597 ( .A1(n505), .A2(G214), .ZN(n464) );
  XNOR2_X1 U598 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U599 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U600 ( .A(KEYINPUT13), .B(KEYINPUT106), .ZN(n472) );
  XOR2_X1 U601 ( .A(KEYINPUT107), .B(KEYINPUT7), .Z(n476) );
  NAND2_X1 U602 ( .A1(n735), .A2(G234), .ZN(n474) );
  XNOR2_X1 U603 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n473) );
  XNOR2_X1 U604 ( .A(n474), .B(n473), .ZN(n484) );
  NAND2_X1 U605 ( .A1(G217), .A2(n484), .ZN(n475) );
  XNOR2_X1 U606 ( .A(n476), .B(n475), .ZN(n481) );
  INV_X1 U607 ( .A(n477), .ZN(n478) );
  XNOR2_X1 U608 ( .A(n515), .B(n478), .ZN(n479) );
  NOR2_X1 U609 ( .A1(G902), .A2(n714), .ZN(n482) );
  XOR2_X1 U610 ( .A(G478), .B(n482), .Z(n552) );
  XNOR2_X1 U611 ( .A(n733), .B(n483), .ZN(n487) );
  XNOR2_X1 U612 ( .A(n485), .B(n455), .ZN(n486) );
  NAND2_X1 U613 ( .A1(G234), .A2(n621), .ZN(n488) );
  XNOR2_X1 U614 ( .A(KEYINPUT20), .B(n488), .ZN(n499) );
  NAND2_X1 U615 ( .A1(n499), .A2(G217), .ZN(n490) );
  XNOR2_X1 U616 ( .A(n492), .B(KEYINPUT14), .ZN(n493) );
  XNOR2_X1 U617 ( .A(KEYINPUT76), .B(n493), .ZN(n495) );
  NAND2_X1 U618 ( .A1(G952), .A2(n495), .ZN(n690) );
  NOR2_X1 U619 ( .A1(G953), .A2(n690), .ZN(n494) );
  XOR2_X1 U620 ( .A(KEYINPUT97), .B(n494), .Z(n574) );
  AND2_X1 U621 ( .A1(n495), .A2(G953), .ZN(n496) );
  NAND2_X1 U622 ( .A1(G902), .A2(n496), .ZN(n575) );
  NOR2_X1 U623 ( .A1(G900), .A2(n575), .ZN(n497) );
  NOR2_X1 U624 ( .A1(n574), .A2(n497), .ZN(n498) );
  XNOR2_X1 U625 ( .A(KEYINPUT86), .B(n498), .ZN(n549) );
  NOR2_X1 U626 ( .A1(n661), .A2(n549), .ZN(n501) );
  NAND2_X1 U627 ( .A1(n499), .A2(G221), .ZN(n500) );
  XOR2_X1 U628 ( .A(KEYINPUT21), .B(n500), .Z(n660) );
  NAND2_X1 U629 ( .A1(n501), .A2(n660), .ZN(n533) );
  XNOR2_X1 U630 ( .A(G113), .B(G116), .ZN(n502) );
  NAND2_X1 U631 ( .A1(n505), .A2(G210), .ZN(n506) );
  XNOR2_X1 U632 ( .A(n509), .B(n508), .ZN(n510) );
  NOR2_X1 U633 ( .A1(n630), .A2(G902), .ZN(n513) );
  INV_X1 U634 ( .A(n613), .ZN(n588) );
  NOR2_X1 U635 ( .A1(n533), .A2(n588), .ZN(n514) );
  NAND2_X1 U636 ( .A1(n646), .A2(n514), .ZN(n567) );
  XNOR2_X1 U637 ( .A(KEYINPUT16), .B(n517), .ZN(n518) );
  XNOR2_X1 U638 ( .A(n522), .B(KEYINPUT18), .ZN(n523) );
  XNOR2_X1 U639 ( .A(n524), .B(n523), .ZN(n525) );
  NAND2_X1 U640 ( .A1(n528), .A2(G210), .ZN(n526) );
  NAND2_X1 U641 ( .A1(G214), .A2(n528), .ZN(n676) );
  XNOR2_X1 U642 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U643 ( .A(n646), .ZN(n649) );
  NAND2_X1 U644 ( .A1(n559), .A2(n552), .ZN(n652) );
  INV_X1 U645 ( .A(n605), .ZN(n664) );
  XNOR2_X1 U646 ( .A(n534), .B(KEYINPUT28), .ZN(n536) );
  INV_X1 U647 ( .A(n535), .ZN(n600) );
  NAND2_X1 U648 ( .A1(n536), .A2(n600), .ZN(n562) );
  NAND2_X1 U649 ( .A1(n680), .A2(n647), .ZN(n538) );
  NAND2_X1 U650 ( .A1(n538), .A2(KEYINPUT47), .ZN(n542) );
  NOR2_X1 U651 ( .A1(KEYINPUT47), .A2(n539), .ZN(n540) );
  NAND2_X1 U652 ( .A1(n540), .A2(n647), .ZN(n541) );
  NAND2_X1 U653 ( .A1(n542), .A2(n541), .ZN(n553) );
  NAND2_X1 U654 ( .A1(n661), .A2(n660), .ZN(n544) );
  XNOR2_X1 U655 ( .A(KEYINPUT112), .B(KEYINPUT30), .ZN(n545) );
  XNOR2_X1 U656 ( .A(n545), .B(KEYINPUT111), .ZN(n546) );
  XNOR2_X1 U657 ( .A(n547), .B(n546), .ZN(n548) );
  INV_X1 U658 ( .A(n549), .ZN(n550) );
  INV_X1 U659 ( .A(n552), .ZN(n560) );
  NOR2_X1 U660 ( .A1(n559), .A2(n560), .ZN(n594) );
  XOR2_X1 U661 ( .A(KEYINPUT75), .B(n554), .Z(n555) );
  XOR2_X1 U662 ( .A(KEYINPUT38), .B(KEYINPUT77), .Z(n556) );
  NAND2_X1 U663 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n676), .A2(n665), .ZN(n566) );
  NOR2_X1 U665 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U666 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n568) );
  XNOR2_X1 U667 ( .A(n569), .B(n568), .ZN(n570) );
  NAND2_X1 U668 ( .A1(n571), .A2(n570), .ZN(n655) );
  INV_X1 U669 ( .A(n652), .ZN(n641) );
  INV_X1 U670 ( .A(n574), .ZN(n578) );
  NOR2_X1 U671 ( .A1(G898), .A2(n575), .ZN(n576) );
  XOR2_X1 U672 ( .A(KEYINPUT98), .B(n576), .Z(n577) );
  NAND2_X1 U673 ( .A1(n578), .A2(n577), .ZN(n579) );
  INV_X1 U674 ( .A(n660), .ZN(n582) );
  XNOR2_X1 U675 ( .A(KEYINPUT22), .B(KEYINPUT74), .ZN(n584) );
  INV_X1 U676 ( .A(n661), .ZN(n586) );
  XNOR2_X1 U677 ( .A(KEYINPUT32), .B(KEYINPUT84), .ZN(n589) );
  NAND2_X1 U678 ( .A1(n665), .A2(n664), .ZN(n590) );
  NOR2_X1 U679 ( .A1(n666), .A2(n665), .ZN(n604) );
  AND2_X1 U680 ( .A1(n613), .A2(n604), .ZN(n591) );
  INV_X1 U681 ( .A(KEYINPUT99), .ZN(n592) );
  NAND2_X1 U682 ( .A1(n595), .A2(n745), .ZN(n598) );
  NAND2_X1 U683 ( .A1(n598), .A2(n597), .ZN(n620) );
  INV_X1 U684 ( .A(n666), .ZN(n599) );
  AND2_X1 U685 ( .A1(n600), .A2(n599), .ZN(n603) );
  NOR2_X1 U686 ( .A1(n605), .A2(n601), .ZN(n602) );
  NAND2_X1 U687 ( .A1(n603), .A2(n602), .ZN(n635) );
  NAND2_X1 U688 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U689 ( .A(KEYINPUT102), .B(n606), .ZN(n671) );
  XOR2_X1 U690 ( .A(KEYINPUT103), .B(n607), .Z(n608) );
  XNOR2_X1 U691 ( .A(KEYINPUT31), .B(n608), .ZN(n651) );
  NAND2_X1 U692 ( .A1(n635), .A2(n651), .ZN(n610) );
  NAND2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n661), .A2(n611), .ZN(n612) );
  NOR2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n614), .A2(n665), .ZN(n632) );
  NAND2_X1 U697 ( .A1(n615), .A2(n632), .ZN(n618) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT65), .ZN(n617) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n656) );
  XOR2_X1 U700 ( .A(KEYINPUT91), .B(n621), .Z(n622) );
  BUF_X1 U701 ( .A(n623), .Z(n627) );
  NAND2_X1 U702 ( .A1(KEYINPUT2), .A2(n654), .ZN(n624) );
  XNOR2_X1 U703 ( .A(KEYINPUT87), .B(n624), .ZN(n625) );
  NOR2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n658) );
  XOR2_X1 U705 ( .A(KEYINPUT63), .B(n631), .Z(G57) );
  XNOR2_X1 U706 ( .A(G101), .B(n632), .ZN(G3) );
  NOR2_X1 U707 ( .A1(n649), .A2(n635), .ZN(n633) );
  XOR2_X1 U708 ( .A(KEYINPUT116), .B(n633), .Z(n634) );
  XNOR2_X1 U709 ( .A(G104), .B(n634), .ZN(G6) );
  NOR2_X1 U710 ( .A1(n652), .A2(n635), .ZN(n640) );
  XOR2_X1 U711 ( .A(KEYINPUT27), .B(KEYINPUT118), .Z(n637) );
  XNOR2_X1 U712 ( .A(G107), .B(KEYINPUT117), .ZN(n636) );
  XNOR2_X1 U713 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U714 ( .A(KEYINPUT26), .B(n638), .ZN(n639) );
  XNOR2_X1 U715 ( .A(n640), .B(n639), .ZN(G9) );
  XOR2_X1 U716 ( .A(KEYINPUT29), .B(KEYINPUT120), .Z(n643) );
  NAND2_X1 U717 ( .A1(n647), .A2(n641), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(n645) );
  XOR2_X1 U719 ( .A(G128), .B(KEYINPUT119), .Z(n644) );
  XNOR2_X1 U720 ( .A(n645), .B(n644), .ZN(G30) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n648), .B(G146), .ZN(G48) );
  NOR2_X1 U723 ( .A1(n649), .A2(n651), .ZN(n650) );
  XOR2_X1 U724 ( .A(G113), .B(n650), .Z(G15) );
  NOR2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U726 ( .A(G116), .B(n653), .Z(G18) );
  XNOR2_X1 U727 ( .A(G134), .B(n654), .ZN(G36) );
  XNOR2_X1 U728 ( .A(G140), .B(n655), .ZN(G42) );
  NAND2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n659), .A2(n628), .ZN(n696) );
  NOR2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(KEYINPUT49), .ZN(n663) );
  NAND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n669) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U735 ( .A(KEYINPUT50), .B(n667), .Z(n668) );
  NOR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U737 ( .A(KEYINPUT121), .B(n670), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT122), .ZN(n674) );
  XNOR2_X1 U740 ( .A(n674), .B(KEYINPUT51), .ZN(n675) );
  NOR2_X1 U741 ( .A1(n691), .A2(n675), .ZN(n687) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n684) );
  INV_X1 U744 ( .A(n680), .ZN(n682) );
  NOR2_X1 U745 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U746 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n685), .A2(n692), .ZN(n686) );
  NOR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT52), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U751 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U752 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n697), .A2(G953), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n698), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U756 ( .A1(n715), .A2(G210), .ZN(n703) );
  XOR2_X1 U757 ( .A(KEYINPUT88), .B(KEYINPUT55), .Z(n700) );
  XNOR2_X1 U758 ( .A(KEYINPUT123), .B(KEYINPUT54), .ZN(n699) );
  XNOR2_X1 U759 ( .A(n700), .B(n699), .ZN(n701) );
  NAND2_X1 U760 ( .A1(n715), .A2(G469), .ZN(n707) );
  XOR2_X1 U761 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n704) );
  NOR2_X1 U762 ( .A1(n720), .A2(n708), .ZN(G54) );
  NAND2_X1 U763 ( .A1(n715), .A2(G475), .ZN(n711) );
  XOR2_X1 U764 ( .A(KEYINPUT59), .B(KEYINPUT96), .Z(n709) );
  XNOR2_X1 U765 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n714), .B(KEYINPUT124), .ZN(n717) );
  NAND2_X1 U767 ( .A1(G478), .A2(n715), .ZN(n716) );
  XNOR2_X1 U768 ( .A(n717), .B(n716), .ZN(n718) );
  NOR2_X1 U769 ( .A1(n720), .A2(n718), .ZN(G63) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n721) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n721), .ZN(n722) );
  NAND2_X1 U772 ( .A1(n722), .A2(G898), .ZN(n723) );
  NAND2_X1 U773 ( .A1(n724), .A2(n723), .ZN(n731) );
  XNOR2_X1 U774 ( .A(n725), .B(G101), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n726), .B(KEYINPUT126), .ZN(n727) );
  XNOR2_X1 U776 ( .A(n727), .B(G110), .ZN(n729) );
  NOR2_X1 U777 ( .A1(n735), .A2(G898), .ZN(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U779 ( .A(n731), .B(n730), .ZN(G69) );
  XOR2_X1 U780 ( .A(n733), .B(n732), .Z(n737) );
  XNOR2_X1 U781 ( .A(n737), .B(n734), .ZN(n736) );
  NAND2_X1 U782 ( .A1(n736), .A2(n735), .ZN(n742) );
  XNOR2_X1 U783 ( .A(n737), .B(G227), .ZN(n738) );
  XNOR2_X1 U784 ( .A(n738), .B(KEYINPUT127), .ZN(n739) );
  NAND2_X1 U785 ( .A1(n739), .A2(G900), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n740), .A2(G953), .ZN(n741) );
  NAND2_X1 U787 ( .A1(n742), .A2(n741), .ZN(G72) );
  XOR2_X1 U788 ( .A(G125), .B(KEYINPUT37), .Z(n743) );
  XNOR2_X1 U789 ( .A(n744), .B(n743), .ZN(G27) );
  XNOR2_X1 U790 ( .A(n745), .B(G122), .ZN(G24) );
  XNOR2_X1 U791 ( .A(n746), .B(G110), .ZN(G12) );
  XNOR2_X1 U792 ( .A(n747), .B(G119), .ZN(G21) );
  XOR2_X1 U793 ( .A(n748), .B(G137), .Z(G39) );
  XOR2_X1 U794 ( .A(n749), .B(G131), .Z(G33) );
endmodule

