//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT65), .Z(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n213), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  INV_X1    g0027(.A(new_n202), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT66), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n229), .A2(G50), .A3(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n211), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n216), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(KEYINPUT73), .ZN(new_n253));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n233), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n255), .B1(new_n210), .B2(G20), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G50), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(G50), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n211), .A2(G33), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  INV_X1    g0063(.A(G58), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT69), .B(G58), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n263), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n261), .B1(new_n262), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n259), .B1(new_n268), .B2(new_n255), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G41), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G1), .A3(G13), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G274), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n210), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND2_X1   g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G41), .A2(G45), .ZN(new_n280));
  OAI22_X1  g0080(.A1(new_n279), .A2(new_n233), .B1(new_n280), .B2(G1), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n272), .A2(KEYINPUT68), .A3(new_n274), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n278), .B1(new_n285), .B2(G226), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(G222), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(G223), .A3(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G77), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n289), .ZN(new_n294));
  INV_X1    g0094(.A(new_n272), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n286), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n286), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n270), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT9), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n270), .A2(new_n303), .B1(G200), .B2(new_n297), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(new_n297), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n255), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT8), .B(G58), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n314), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT15), .B(G87), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(new_n262), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n312), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n258), .A2(G77), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(new_n256), .B2(G77), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT71), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G20), .A2(G77), .ZN(new_n323));
  INV_X1    g0123(.A(new_n260), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n323), .B1(new_n316), .B2(new_n262), .C1(new_n324), .C2(new_n313), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n255), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT71), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(new_n320), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n278), .B1(new_n285), .B2(G244), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n289), .A2(G232), .A3(new_n290), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n289), .A2(G238), .A3(G1698), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n331), .B(new_n332), .C1(new_n207), .C2(new_n289), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n295), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n298), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT72), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n328), .A2(new_n322), .B1(new_n335), .B2(new_n298), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n330), .A2(new_n334), .A3(new_n300), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n338), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n329), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT70), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n330), .A2(new_n334), .A3(new_n345), .A4(G190), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT70), .B1(new_n335), .B2(G200), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n335), .A2(new_n306), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n344), .B(new_n346), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n253), .B1(new_n311), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n310), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n308), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n343), .A2(new_n349), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n353), .A2(KEYINPUT73), .A3(new_n302), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n267), .A2(new_n258), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n256), .B2(new_n267), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n228), .B1(new_n266), .B2(new_n218), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n211), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  NOR4_X1   g0165(.A1(new_n361), .A2(new_n362), .A3(new_n365), .A4(G20), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n360), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n312), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n360), .A2(new_n367), .A3(KEYINPUT16), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n358), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n276), .A2(new_n277), .ZN(new_n373));
  INV_X1    g0173(.A(G274), .ZN(new_n374));
  INV_X1    g0174(.A(new_n233), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n271), .ZN(new_n376));
  AND2_X1   g0176(.A1(new_n272), .A2(new_n274), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n373), .A2(new_n376), .B1(new_n377), .B2(G232), .ZN(new_n378));
  OR2_X1    g0178(.A1(G223), .A2(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G226), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n379), .B(new_n381), .C1(new_n361), .C2(new_n362), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n295), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n298), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT79), .ZN(new_n388));
  INV_X1    g0188(.A(new_n383), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G223), .A2(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n380), .B2(G1698), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n391), .B2(new_n289), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n388), .B1(new_n392), .B2(new_n272), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n384), .A2(KEYINPUT79), .A3(new_n295), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n378), .A2(new_n300), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n387), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT18), .B1(new_n372), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n264), .A2(KEYINPUT69), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT69), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G58), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n202), .B1(new_n402), .B2(G68), .ZN(new_n403));
  INV_X1    g0203(.A(G159), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n403), .A2(new_n211), .B1(new_n404), .B2(new_n324), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n287), .A2(new_n211), .A3(new_n288), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n365), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n218), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n369), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(new_n255), .A3(new_n371), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n357), .ZN(new_n412));
  INV_X1    g0212(.A(new_n395), .ZN(new_n413));
  INV_X1    g0213(.A(new_n396), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n413), .A2(new_n414), .B1(new_n298), .B2(new_n386), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n412), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n398), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT80), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n393), .A2(new_n378), .A3(new_n394), .A4(new_n306), .ZN(new_n420));
  INV_X1    g0220(.A(G200), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n373), .A2(new_n376), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n377), .A2(G232), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n272), .B1(new_n382), .B2(new_n383), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n419), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n420), .A2(new_n426), .A3(new_n419), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n372), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT81), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT17), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n372), .B(new_n434), .C1(new_n427), .C2(new_n428), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n418), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n351), .A2(new_n355), .A3(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n293), .B2(new_n262), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n255), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT11), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT75), .A3(new_n443), .ZN(new_n444));
  OR3_X1    g0244(.A1(new_n258), .A2(KEYINPUT12), .A3(G68), .ZN(new_n445));
  OAI21_X1  g0245(.A(KEYINPUT12), .B1(new_n258), .B2(G68), .ZN(new_n446));
  AOI22_X1  g0246(.A1(G68), .A2(new_n256), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT75), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n442), .A2(new_n443), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT76), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT13), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT74), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n219), .B1(new_n283), .B2(new_n284), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n278), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n272), .A2(KEYINPUT68), .A3(new_n274), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT68), .B1(new_n272), .B2(new_n274), .ZN(new_n459));
  OAI21_X1  g0259(.A(G238), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(KEYINPUT74), .A3(new_n422), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n380), .A2(new_n290), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n289), .B(new_n463), .C1(G232), .C2(new_n290), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G97), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n272), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n454), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  AOI211_X1 g0268(.A(KEYINPUT13), .B(new_n466), .C1(new_n457), .C2(new_n461), .ZN(new_n469));
  OAI21_X1  g0269(.A(G200), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n468), .A2(new_n469), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G190), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n453), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT78), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n474), .A3(G179), .ZN(new_n475));
  NOR3_X1   g0275(.A1(new_n456), .A2(new_n455), .A3(new_n278), .ZN(new_n476));
  AOI21_X1  g0276(.A(KEYINPUT74), .B1(new_n460), .B2(new_n422), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n467), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT13), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n462), .A2(new_n454), .A3(new_n467), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(G179), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT78), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n298), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT14), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(KEYINPUT77), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT77), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n488), .B(KEYINPUT14), .C1(new_n471), .C2(new_n298), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n483), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n453), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n473), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n437), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n210), .A2(G45), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G257), .A3(new_n272), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n376), .A2(new_n496), .A3(new_n494), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G244), .B(new_n290), .C1(new_n361), .C2(new_n362), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n289), .A2(KEYINPUT4), .A3(G244), .A4(new_n290), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n295), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT83), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT83), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n507), .A2(new_n510), .A3(new_n295), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n500), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT84), .B1(new_n512), .B2(new_n421), .ZN(new_n513));
  INV_X1    g0313(.A(new_n500), .ZN(new_n514));
  INV_X1    g0314(.A(new_n511), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n510), .B1(new_n507), .B2(new_n295), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(G200), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n210), .A2(G33), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n258), .A2(new_n520), .A3(new_n233), .A4(new_n254), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G97), .ZN(new_n522));
  INV_X1    g0322(.A(new_n258), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(G97), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT82), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n522), .B(new_n526), .C1(G97), .C2(new_n523), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n529), .A2(new_n206), .A3(G107), .ZN(new_n530));
  XNOR2_X1  g0330(.A(G97), .B(G107), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n530), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n532), .A2(new_n211), .B1(new_n293), .B2(new_n324), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n207), .B1(new_n407), .B2(new_n408), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n255), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n500), .B1(new_n295), .B2(new_n507), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(G190), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n513), .A2(new_n519), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n508), .A2(new_n514), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n298), .B1(new_n528), .B2(new_n535), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n517), .B2(G179), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT85), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n495), .A2(G250), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(new_n295), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n272), .A2(KEYINPUT85), .A3(G250), .A4(new_n495), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n545), .A2(new_n546), .B1(new_n496), .B2(new_n376), .ZN(new_n547));
  OAI211_X1 g0347(.A(G244), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n548));
  OAI211_X1 g0348(.A(G238), .B(new_n290), .C1(new_n361), .C2(new_n362), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G116), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n295), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n521), .A2(new_n220), .ZN(new_n555));
  INV_X1    g0355(.A(new_n316), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(new_n258), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n289), .A2(new_n211), .A3(G68), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n211), .B1(new_n465), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(G87), .B2(new_n208), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n559), .B1(new_n262), .B2(new_n206), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI211_X1 g0363(.A(new_n555), .B(new_n557), .C1(new_n563), .C2(new_n255), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n554), .B(new_n564), .C1(new_n306), .C2(new_n553), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n557), .B1(new_n563), .B2(new_n255), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n521), .B2(new_n316), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n553), .A2(new_n298), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n547), .A2(new_n300), .A3(new_n552), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n539), .A2(new_n542), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n523), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n521), .B2(new_n573), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n573), .A2(G20), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT86), .B1(new_n255), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n255), .A2(KEYINPUT86), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n506), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT20), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n580), .ZN(new_n584));
  OAI211_X1 g0384(.A(KEYINPUT20), .B(new_n582), .C1(new_n584), .C2(new_n578), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n576), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G264), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n588));
  OAI211_X1 g0388(.A(G257), .B(new_n290), .C1(new_n361), .C2(new_n362), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n287), .A2(G303), .A3(new_n288), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n295), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n497), .A2(G270), .A3(new_n272), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n499), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n587), .A2(G179), .A3(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n595), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n298), .B1(new_n598), .B2(new_n592), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n587), .A2(KEYINPUT21), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n582), .B1(new_n584), .B2(new_n578), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n575), .B1(new_n604), .B2(new_n585), .ZN(new_n605));
  OAI21_X1  g0405(.A(G169), .B1(new_n593), .B2(new_n595), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n601), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n597), .A2(new_n600), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n497), .A2(G264), .A3(new_n272), .ZN(new_n609));
  OAI211_X1 g0409(.A(G257), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n610));
  NAND2_X1  g0410(.A1(G33), .A2(G294), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n221), .A2(G1698), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n361), .B2(new_n362), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT88), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT88), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n289), .A2(new_n616), .A3(new_n613), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n612), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n295), .B1(new_n618), .B2(KEYINPUT89), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n617), .ZN(new_n620));
  INV_X1    g0420(.A(new_n612), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT89), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n499), .B(new_n609), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n298), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n621), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT89), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n618), .A2(KEYINPUT89), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n295), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(new_n300), .A3(new_n499), .A4(new_n609), .ZN(new_n630));
  OR3_X1    g0430(.A1(new_n258), .A2(KEYINPUT25), .A3(G107), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT25), .B1(new_n258), .B2(G107), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n631), .B(new_n632), .C1(new_n207), .C2(new_n521), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT87), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n550), .A2(G20), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT23), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n211), .B2(G107), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n636), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n211), .B(G87), .C1(new_n361), .C2(new_n362), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n642), .A2(KEYINPUT22), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(KEYINPUT22), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT24), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n255), .B1(new_n645), .B2(KEYINPUT24), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n635), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n624), .A2(new_n630), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n623), .A2(G200), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n633), .B(KEYINPUT87), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n643), .A2(new_n644), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n640), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT24), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n312), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n652), .B1(new_n656), .B2(new_n646), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n629), .A2(G190), .A3(new_n499), .A4(new_n609), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n651), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n598), .A2(new_n592), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(G200), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n661), .B(new_n605), .C1(new_n306), .C2(new_n660), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n608), .A2(new_n650), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n493), .A2(new_n572), .A3(new_n663), .ZN(G372));
  INV_X1    g0464(.A(new_n302), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n372), .A2(KEYINPUT18), .A3(new_n397), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n416), .B1(new_n412), .B2(new_n415), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n474), .B1(new_n471), .B2(G179), .ZN(new_n669));
  NOR4_X1   g0469(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT78), .A4(new_n300), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n486), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n487), .A2(new_n489), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n491), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(new_n343), .ZN(new_n674));
  INV_X1    g0474(.A(new_n473), .ZN(new_n675));
  INV_X1    g0475(.A(new_n427), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n420), .A2(new_n426), .A3(new_n419), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n412), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n435), .B1(new_n678), .B2(new_n430), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n668), .B1(new_n674), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n665), .B1(new_n681), .B2(new_n353), .ZN(new_n682));
  INV_X1    g0482(.A(new_n570), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n512), .A2(new_n300), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n571), .A2(KEYINPUT26), .A3(new_n684), .A4(new_n541), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n565), .A2(new_n570), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n542), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n683), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n597), .A2(new_n600), .A3(new_n607), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n597), .A2(new_n600), .A3(new_n607), .A4(KEYINPUT90), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n657), .B1(new_n298), .B2(new_n623), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n692), .A2(new_n693), .B1(new_n694), .B2(new_n630), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n539), .A2(new_n542), .A3(new_n571), .A4(new_n659), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n689), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n682), .B1(new_n493), .B2(new_n698), .ZN(G369));
  NAND3_X1  g0499(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT27), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(G213), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G343), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n587), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n692), .B2(new_n693), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n690), .A2(new_n706), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n662), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n650), .A2(new_n705), .ZN(new_n712));
  INV_X1    g0512(.A(new_n705), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n659), .B1(new_n657), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n712), .B1(new_n714), .B2(new_n650), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n690), .A2(new_n713), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT91), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n712), .B1(new_n720), .B2(new_n715), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n718), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n214), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n231), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT94), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n690), .B1(new_n694), .B2(new_n630), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n689), .B1(new_n731), .B2(new_n696), .ZN(new_n732));
  AND4_X1   g0532(.A1(new_n730), .A2(new_n732), .A3(KEYINPUT29), .A4(new_n713), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n732), .A2(new_n713), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n730), .B1(new_n734), .B2(KEYINPUT29), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n698), .B2(new_n705), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n733), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G330), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n547), .A2(new_n552), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n740), .A2(new_n596), .A3(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(new_n517), .A3(new_n623), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n740), .B(new_n609), .C1(new_n619), .C2(new_n622), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT92), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT92), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n629), .A2(new_n746), .A3(new_n740), .A4(new_n609), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n596), .A2(new_n537), .A3(G179), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT30), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n748), .B1(new_n744), .B2(KEYINPUT92), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT30), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n753), .A3(new_n747), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n743), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n713), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n755), .A2(KEYINPUT93), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT93), .ZN(new_n760));
  AND4_X1   g0560(.A1(new_n753), .A2(new_n745), .A3(new_n747), .A4(new_n749), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n753), .B1(new_n752), .B2(new_n747), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n742), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(new_n763), .B2(new_n757), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT31), .B1(new_n763), .B2(new_n705), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n572), .A2(new_n663), .A3(new_n705), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n739), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n738), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n729), .B1(new_n771), .B2(G1), .ZN(G364));
  INV_X1    g0572(.A(G13), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n210), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n724), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n739), .B1(new_n707), .B2(new_n709), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n711), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n723), .A2(new_n363), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G355), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G116), .B2(new_n214), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n723), .A2(new_n289), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G45), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n232), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n251), .A2(G45), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G13), .A2(G33), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n233), .B1(G20), .B2(new_n298), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n777), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n211), .A2(G179), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n797), .A2(new_n306), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n207), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n211), .A2(new_n300), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n797), .A2(G190), .A3(G200), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n803), .A2(new_n218), .B1(new_n804), .B2(new_n220), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n801), .A2(new_n306), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n799), .B(new_n805), .C1(G50), .C2(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n306), .A2(G179), .A3(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n211), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT95), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G97), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G190), .A2(G200), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n797), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n404), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n800), .A2(new_n812), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n800), .A2(G190), .A3(new_n421), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n289), .B1(new_n816), .B2(new_n293), .C1(new_n266), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n807), .A2(new_n811), .A3(new_n815), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(KEYINPUT33), .B(G317), .ZN(new_n821));
  INV_X1    g0621(.A(new_n817), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n802), .A2(new_n821), .B1(new_n822), .B2(G322), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT96), .Z(new_n824));
  INV_X1    g0624(.A(G311), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n816), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n813), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n289), .B(new_n826), .C1(G329), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n809), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(G294), .ZN(new_n830));
  INV_X1    g0630(.A(new_n798), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(G283), .ZN(new_n832));
  INV_X1    g0632(.A(new_n804), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n806), .A2(G326), .B1(new_n833), .B2(G303), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n828), .A2(new_n830), .A3(new_n832), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n820), .B1(new_n824), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n796), .B1(new_n836), .B2(new_n793), .ZN(new_n837));
  INV_X1    g0637(.A(new_n792), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n837), .B1(new_n710), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n780), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  INV_X1    g0641(.A(new_n793), .ZN(new_n842));
  INV_X1    g0642(.A(new_n816), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n822), .A2(G143), .B1(new_n843), .B2(G159), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  INV_X1    g0646(.A(new_n806), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n844), .B1(new_n803), .B2(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT34), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n798), .A2(new_n218), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n363), .B(new_n852), .C1(G132), .C2(new_n827), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n829), .A2(new_n402), .B1(new_n833), .B2(G50), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n850), .A2(new_n851), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G294), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n817), .A2(new_n856), .B1(new_n816), .B2(new_n573), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n289), .B(new_n857), .C1(G311), .C2(new_n827), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n802), .A2(G283), .B1(new_n806), .B2(G303), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n833), .A2(G107), .B1(new_n831), .B2(G87), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n858), .A2(new_n811), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n842), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n793), .A2(new_n790), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n778), .B(new_n862), .C1(new_n293), .C2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n329), .A2(new_n705), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n342), .B1(new_n339), .B2(new_n340), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n337), .A2(KEYINPUT72), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n349), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT97), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n343), .A2(new_n865), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n343), .A2(KEYINPUT97), .A3(new_n349), .A4(new_n865), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n864), .B1(new_n873), .B2(new_n791), .ZN(new_n874));
  INV_X1    g0674(.A(new_n873), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n698), .B2(new_n705), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n697), .A2(new_n873), .A3(new_n713), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n770), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n778), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n770), .A2(new_n878), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n874), .B1(new_n880), .B2(new_n881), .ZN(G384));
  NOR2_X1   g0682(.A1(new_n774), .A2(new_n210), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n412), .A2(new_n415), .ZN(new_n884));
  INV_X1    g0684(.A(new_n703), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n412), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n429), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n429), .A2(new_n889), .A3(new_n884), .A4(new_n886), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT99), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n890), .A2(KEYINPUT98), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n890), .B2(KEYINPUT98), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(KEYINPUT98), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT99), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n890), .A2(KEYINPUT98), .A3(new_n891), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n679), .A2(new_n668), .ZN(new_n900));
  INV_X1    g0700(.A(new_n886), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n894), .A2(new_n899), .A3(KEYINPUT38), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n888), .A2(new_n890), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT101), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n900), .A2(new_n901), .B1(new_n888), .B2(new_n890), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT101), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT38), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n903), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n491), .A2(new_n705), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n673), .A2(new_n675), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n491), .B(new_n705), .C1(new_n490), .C2(new_n473), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n875), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n756), .B1(new_n755), .B2(new_n713), .ZN(new_n916));
  INV_X1    g0716(.A(new_n572), .ZN(new_n917));
  AND4_X1   g0717(.A1(new_n608), .A2(new_n650), .A3(new_n659), .A4(new_n662), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n918), .A3(new_n713), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n763), .A2(new_n757), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n911), .A2(KEYINPUT40), .A3(new_n915), .A4(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT102), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n915), .A2(new_n921), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n905), .A2(KEYINPUT101), .A3(new_n906), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n909), .B1(new_n908), .B2(KEYINPUT38), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n926), .B1(new_n929), .B2(new_n903), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n925), .A2(new_n930), .A3(KEYINPUT102), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n436), .A2(new_n886), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n896), .A2(new_n898), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n934), .B2(new_n888), .ZN(new_n935));
  AOI21_X1  g0735(.A(KEYINPUT38), .B1(new_n935), .B2(new_n899), .ZN(new_n936));
  INV_X1    g0736(.A(new_n903), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n915), .B(new_n921), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n926), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n437), .A2(new_n492), .A3(new_n921), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n942), .A2(new_n943), .A3(new_n739), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT39), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n911), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n491), .B(new_n713), .C1(new_n671), .C2(new_n672), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT100), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n490), .A2(KEYINPUT100), .A3(new_n491), .A4(new_n713), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n894), .A2(new_n899), .A3(new_n902), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n906), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n947), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n343), .A2(new_n705), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n877), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n913), .A2(new_n914), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n954), .A2(new_n903), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n961), .A2(new_n962), .B1(new_n418), .B2(new_n703), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n682), .B1(new_n738), .B2(new_n493), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  AOI21_X1  g0766(.A(new_n883), .B1(new_n945), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n945), .ZN(new_n968));
  INV_X1    g0768(.A(new_n532), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT35), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(KEYINPUT35), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n970), .A2(G116), .A3(new_n234), .A4(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT36), .ZN(new_n973));
  OAI21_X1  g0773(.A(G77), .B1(new_n266), .B2(new_n218), .ZN(new_n974));
  INV_X1    g0774(.A(new_n201), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n231), .A2(new_n974), .B1(new_n218), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n976), .A2(G1), .A3(new_n773), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n968), .A2(new_n973), .A3(new_n977), .ZN(G367));
  NAND2_X1  g0778(.A1(new_n720), .A2(new_n715), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n536), .A2(new_n705), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n539), .A2(new_n542), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n684), .A2(new_n541), .A3(new_n705), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n979), .A2(KEYINPUT42), .A3(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n542), .B1(new_n981), .B2(new_n650), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n713), .ZN(new_n987));
  OAI21_X1  g0787(.A(KEYINPUT42), .B1(new_n979), .B2(new_n984), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n564), .A2(new_n713), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n571), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT103), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT103), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n570), .C2(new_n990), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n989), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT104), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT104), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n989), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT43), .B2(new_n994), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n997), .A2(new_n1002), .A3(new_n999), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n718), .A2(new_n984), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1004), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n724), .B(KEYINPUT41), .Z(new_n1008));
  XOR2_X1   g0808(.A(new_n711), .B(KEYINPUT107), .Z(new_n1009));
  OR2_X1    g0809(.A1(new_n720), .A2(new_n715), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(KEYINPUT106), .A3(new_n979), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT106), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n720), .A2(new_n715), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n711), .A2(KEYINPUT107), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1015), .B1(new_n1017), .B2(new_n1014), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n771), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT108), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n771), .A2(new_n1018), .A3(KEYINPUT108), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n721), .A2(new_n983), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT44), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n721), .A2(new_n983), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n1026));
  XNOR2_X1  g0826(.A(new_n1025), .B(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n717), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1024), .A2(new_n718), .A3(new_n1027), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1021), .A2(new_n1022), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1008), .B1(new_n1031), .B2(new_n771), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1007), .B1(new_n1032), .B2(new_n776), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n794), .B1(new_n214), .B2(new_n316), .C1(new_n785), .C2(new_n244), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1034), .A2(new_n777), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n798), .A2(new_n206), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n847), .A2(new_n825), .B1(new_n207), .B2(new_n809), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G294), .C2(new_n802), .ZN(new_n1038));
  INV_X1    g0838(.A(G283), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n363), .B1(new_n816), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(G303), .ZN(new_n1041));
  INV_X1    g0841(.A(G317), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n817), .A2(new_n1041), .B1(new_n813), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n804), .A2(new_n573), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1040), .B(new_n1043), .C1(KEYINPUT46), .C2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1038), .B(new_n1045), .C1(KEYINPUT46), .C2(new_n1044), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n810), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n218), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n817), .A2(new_n845), .B1(new_n816), .B2(new_n201), .ZN(new_n1049));
  AOI211_X1 g0849(.A(new_n363), .B(new_n1049), .C1(G137), .C2(new_n827), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n802), .A2(G159), .B1(new_n806), .B2(G143), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n798), .A2(new_n293), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n402), .B2(new_n833), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1046), .B1(new_n1048), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT109), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT47), .Z(new_n1057));
  OAI221_X1 g0857(.A(new_n1035), .B1(new_n838), .B2(new_n994), .C1(new_n1057), .C2(new_n842), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1033), .A2(new_n1058), .ZN(G387));
  NAND2_X1  g0859(.A1(new_n1018), .A2(new_n776), .ZN(new_n1060));
  INV_X1    g0860(.A(G50), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n817), .A2(new_n1061), .B1(new_n816), .B2(new_n218), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n363), .B(new_n1062), .C1(G150), .C2(new_n827), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n810), .A2(new_n556), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n804), .A2(new_n293), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1036), .B(new_n1065), .C1(G159), .C2(new_n806), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n803), .A2(new_n267), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n289), .B1(new_n827), .B2(G326), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n809), .A2(new_n1039), .B1(new_n804), .B2(new_n856), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n822), .A2(G317), .B1(new_n843), .B2(G303), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT110), .B(G322), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(new_n803), .B2(new_n825), .C1(new_n847), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1074), .B2(new_n1073), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT49), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1069), .B1(new_n573), .B2(new_n798), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1068), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n793), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n726), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n781), .A2(new_n1082), .B1(new_n207), .B2(new_n723), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n241), .A2(new_n786), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n314), .A2(new_n1061), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT50), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n726), .B(new_n786), .C1(new_n218), .C2(new_n293), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n784), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1083), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n778), .B1(new_n1089), .B2(new_n794), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1081), .B(new_n1090), .C1(new_n715), .C2(new_n838), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1019), .A2(new_n724), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n771), .A2(new_n1018), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1060), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(G393));
  NAND3_X1  g0894(.A1(new_n1029), .A2(KEYINPUT111), .A3(new_n1030), .ZN(new_n1095));
  OR3_X1    g0895(.A1(new_n1028), .A2(KEYINPUT111), .A3(new_n717), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1095), .A2(new_n1096), .A3(new_n1019), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1031), .A2(new_n1097), .A3(new_n724), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n829), .A2(G116), .B1(new_n843), .B2(G294), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1041), .B2(new_n803), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT112), .Z(new_n1101));
  OAI22_X1  g0901(.A1(new_n847), .A2(new_n1042), .B1(new_n825), .B2(new_n817), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n363), .B1(new_n813), .B2(new_n1072), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n799), .B(new_n1104), .C1(G283), .C2(new_n833), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n218), .A2(new_n804), .B1(new_n798), .B2(new_n220), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n363), .B1(new_n827), .B2(G143), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n313), .B2(new_n816), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(new_n975), .C2(new_n802), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n847), .A2(new_n845), .B1(new_n404), .B2(new_n817), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT51), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n810), .A2(G77), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1110), .A2(new_n1113), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n842), .B1(new_n1106), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n784), .A2(new_n248), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n795), .B1(G97), .B2(new_n723), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n778), .B(new_n1117), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT113), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n792), .B2(new_n984), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n776), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1098), .A2(new_n1124), .ZN(G390));
  AOI21_X1  g0925(.A(new_n960), .B1(new_n769), .B2(new_n873), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n739), .B1(new_n768), .B2(new_n920), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n915), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n959), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n769), .A2(new_n915), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n921), .A2(G330), .A3(new_n873), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n913), .A3(new_n914), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n732), .A2(new_n873), .A3(new_n713), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n958), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AND4_X1   g0935(.A1(KEYINPUT114), .A2(new_n1130), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n769), .B2(new_n915), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT114), .B1(new_n1137), .B2(new_n1132), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1129), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n437), .A2(new_n492), .A3(new_n1127), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n682), .B(new_n1140), .C1(new_n738), .C2(new_n493), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n954), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT39), .B1(new_n929), .B2(new_n903), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n1144), .A2(new_n1145), .B1(new_n952), .B2(new_n961), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1134), .A2(new_n960), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n952), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n911), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1130), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n952), .B1(new_n959), .B2(new_n960), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n947), .B2(new_n955), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1149), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1128), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1150), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1139), .A2(new_n1150), .A3(new_n1154), .A4(new_n1142), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n724), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1150), .A2(new_n1154), .A3(new_n776), .ZN(new_n1159));
  INV_X1    g0959(.A(G128), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1160), .A2(new_n847), .B1(new_n803), .B2(new_n846), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n975), .B2(new_n831), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n822), .A2(G132), .B1(new_n827), .B2(G125), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT54), .B(G143), .Z(new_n1164));
  AOI21_X1  g0964(.A(new_n363), .B1(new_n843), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n804), .A2(new_n845), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT53), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n810), .A2(G159), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1162), .A2(new_n1166), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n816), .A2(new_n206), .B1(new_n813), .B2(new_n856), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n289), .B(new_n1171), .C1(G116), .C2(new_n822), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n852), .B1(G87), .B2(new_n833), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n802), .A2(G107), .B1(new_n806), .B2(G283), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1172), .A2(new_n1114), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n842), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n778), .B(new_n1176), .C1(new_n267), .C2(new_n863), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n947), .A2(new_n955), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1177), .B1(new_n1179), .B2(new_n791), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1158), .A2(new_n1159), .A3(new_n1180), .ZN(G378));
  NAND2_X1  g0981(.A1(new_n270), .A2(new_n885), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT55), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n311), .B(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1186), .A2(new_n790), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n778), .B1(new_n201), .B2(new_n863), .ZN(new_n1188));
  OR2_X1    g0988(.A1(new_n289), .A2(G41), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1189), .B(new_n1061), .C1(G33), .C2(G41), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT115), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n817), .A2(new_n207), .B1(new_n813), .B2(new_n1039), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1189), .B(new_n1192), .C1(new_n556), .C2(new_n843), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1065), .B1(G97), .B2(new_n802), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n573), .B2(new_n847), .C1(new_n266), .C2(new_n798), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1194), .A2(new_n1196), .A3(new_n1048), .ZN(new_n1197));
  XOR2_X1   g0997(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1191), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT117), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n817), .A2(new_n1160), .B1(new_n816), .B2(new_n846), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G132), .B2(new_n802), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n806), .A2(G125), .B1(new_n833), .B2(new_n1164), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n1047), .C2(new_n845), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n827), .C2(G124), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n404), .B2(new_n798), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1205), .B2(KEYINPUT59), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1206), .A2(new_n1209), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1210));
  AND2_X1   g1010(.A1(new_n1201), .A2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1188), .B1(new_n1211), .B2(new_n842), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1187), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT120), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n956), .A2(new_n963), .A3(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n956), .B2(new_n963), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n739), .B1(new_n938), .B2(new_n926), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT119), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1186), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n932), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n932), .B2(new_n1218), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1217), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n922), .A2(new_n923), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT102), .B1(new_n925), .B2(new_n930), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1218), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1220), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n932), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n964), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1223), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1213), .B1(new_n1231), .B2(new_n776), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1157), .B2(new_n1142), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1228), .A2(new_n964), .A3(new_n1229), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n964), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(new_n724), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1157), .A2(new_n1142), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT57), .B1(new_n1231), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1232), .B1(new_n1238), .B2(new_n1240), .ZN(G375));
  INV_X1    g1041(.A(new_n1008), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1141), .B(new_n1129), .C1(new_n1136), .C2(new_n1138), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1143), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n913), .A2(new_n914), .A3(new_n790), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n793), .A2(G68), .A3(new_n790), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n816), .A2(new_n207), .B1(new_n813), .B2(new_n1041), .ZN(new_n1247));
  AOI211_X1 g1047(.A(new_n289), .B(new_n1247), .C1(G283), .C2(new_n822), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1052), .B1(G116), .B2(new_n802), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n806), .A2(G294), .B1(new_n833), .B2(G97), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1248), .A2(new_n1064), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT121), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n817), .A2(new_n846), .B1(new_n813), .B2(new_n1160), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n363), .B(new_n1254), .C1(G150), .C2(new_n843), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n810), .A2(G50), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G159), .A2(new_n833), .B1(new_n831), .B2(new_n402), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G132), .A2(new_n806), .B1(new_n802), .B2(new_n1164), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1253), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n778), .B(new_n1246), .C1(new_n1261), .C2(new_n793), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1139), .A2(new_n776), .B1(new_n1245), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1244), .A2(new_n1263), .ZN(G381));
  OR4_X1    g1064(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(new_n1265), .A2(G387), .A3(G378), .A4(G381), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(G375), .B(KEYINPUT122), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(KEYINPUT123), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(KEYINPUT123), .ZN(new_n1270));
  OR2_X1    g1070(.A1(new_n1269), .A2(new_n1270), .ZN(G407));
  INV_X1    g1071(.A(G378), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1267), .A2(G213), .A3(new_n704), .A4(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G213), .B(new_n1273), .C1(new_n1269), .C2(new_n1270), .ZN(G409));
  XNOR2_X1  g1074(.A(G393), .B(new_n840), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1033), .A2(new_n1058), .A3(G390), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G390), .B1(new_n1033), .B2(new_n1058), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(G390), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G387), .A2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1033), .A2(G390), .A3(new_n1058), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(new_n1275), .A3(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1279), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT125), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT125), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1279), .A2(new_n1283), .A3(new_n1287), .A4(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1232), .C1(new_n1238), .C2(new_n1240), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n776), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1213), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI221_X4 g1093(.A(new_n1008), .B1(new_n1157), .B2(new_n1142), .C1(new_n1223), .C2(new_n1230), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1272), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1290), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n704), .A2(G213), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT60), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1243), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1137), .A2(new_n1132), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT114), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1137), .A2(KEYINPUT114), .A3(new_n1132), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(KEYINPUT60), .A3(new_n1141), .A4(new_n1129), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1299), .A2(new_n1305), .A3(new_n724), .A4(new_n1143), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1263), .ZN(new_n1307));
  INV_X1    g1107(.A(G384), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1306), .A2(G384), .A3(new_n1263), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1296), .A2(new_n1297), .A3(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(KEYINPUT63), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT63), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1306), .A2(G384), .A3(new_n1263), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G384), .B1(new_n1306), .B2(new_n1263), .ZN(new_n1319));
  OAI21_X1  g1119(.A(KEYINPUT124), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n704), .A2(G213), .A3(G2897), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(KEYINPUT124), .B(new_n1321), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT124), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n1323), .A2(new_n1324), .B1(new_n1312), .B2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1316), .B1(new_n1317), .B2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1289), .B(new_n1315), .C1(new_n1314), .C2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1312), .A2(new_n1325), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1321), .B1(new_n1311), .B2(KEYINPUT124), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1324), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1329), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  AOI22_X1  g1132(.A1(new_n1290), .A2(new_n1295), .B1(G213), .B2(new_n704), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1284), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT62), .ZN(new_n1335));
  AND4_X1   g1135(.A1(new_n1335), .A2(new_n1296), .A3(new_n1297), .A4(new_n1312), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT126), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT61), .B1(new_n1317), .B2(new_n1326), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1333), .A2(new_n1335), .A3(new_n1312), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1340), .A2(new_n1338), .A3(KEYINPUT126), .A4(new_n1341), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1279), .A2(new_n1283), .A3(KEYINPUT127), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT127), .B1(new_n1279), .B2(new_n1283), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1328), .B1(new_n1339), .B2(new_n1346), .ZN(G405));
  NAND2_X1  g1147(.A1(G375), .A2(new_n1272), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(new_n1290), .ZN(new_n1349));
  XNOR2_X1  g1149(.A(new_n1349), .B(new_n1311), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1351));
  XOR2_X1   g1151(.A(new_n1350), .B(new_n1351), .Z(G402));
endmodule


