

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  INV_X1 U322 ( .A(G99GAT), .ZN(n311) );
  XNOR2_X1 U323 ( .A(n323), .B(n322), .ZN(n325) );
  INV_X1 U324 ( .A(KEYINPUT18), .ZN(n322) );
  XNOR2_X1 U325 ( .A(n317), .B(n316), .ZN(n321) );
  XNOR2_X1 U326 ( .A(n312), .B(n311), .ZN(n317) );
  XNOR2_X1 U327 ( .A(n338), .B(n376), .ZN(n517) );
  NAND2_X1 U328 ( .A1(n510), .A2(n515), .ZN(n506) );
  OR2_X1 U329 ( .A1(n454), .A2(n453), .ZN(n455) );
  NOR2_X1 U330 ( .A1(n362), .A2(n361), .ZN(n363) );
  XOR2_X1 U331 ( .A(G127GAT), .B(KEYINPUT0), .Z(n313) );
  XNOR2_X1 U332 ( .A(n463), .B(KEYINPUT64), .ZN(n464) );
  XNOR2_X1 U333 ( .A(n331), .B(n435), .ZN(n332) );
  XNOR2_X1 U334 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U335 ( .A(n465), .B(n464), .ZN(n526) );
  XNOR2_X1 U336 ( .A(n333), .B(n332), .ZN(n335) );
  XNOR2_X1 U337 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U338 ( .A(n325), .B(n324), .ZN(n330) );
  XNOR2_X1 U339 ( .A(n358), .B(KEYINPUT26), .ZN(n568) );
  INV_X1 U340 ( .A(n568), .ZN(n544) );
  OR2_X1 U341 ( .A1(n482), .A2(n481), .ZN(n504) );
  XNOR2_X1 U342 ( .A(n473), .B(KEYINPUT123), .ZN(n563) );
  XOR2_X1 U343 ( .A(KEYINPUT108), .B(n505), .Z(n510) );
  XNOR2_X1 U344 ( .A(n327), .B(n326), .ZN(n527) );
  XNOR2_X1 U345 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U346 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U347 ( .A(n477), .B(n476), .ZN(G1349GAT) );
  XNOR2_X1 U348 ( .A(n450), .B(n449), .ZN(G1330GAT) );
  INV_X1 U349 ( .A(KEYINPUT37), .ZN(n415) );
  XOR2_X1 U350 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n291) );
  XNOR2_X1 U351 ( .A(G141GAT), .B(KEYINPUT4), .ZN(n290) );
  XNOR2_X1 U352 ( .A(n291), .B(n290), .ZN(n307) );
  XOR2_X1 U353 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n293) );
  NAND2_X1 U354 ( .A1(G225GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U355 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U356 ( .A(KEYINPUT94), .B(n294), .ZN(n305) );
  XOR2_X1 U357 ( .A(G148GAT), .B(G57GAT), .Z(n296) );
  XNOR2_X1 U358 ( .A(G120GAT), .B(G162GAT), .ZN(n295) );
  XNOR2_X1 U359 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U360 ( .A(n297), .B(G85GAT), .Z(n299) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(n313), .ZN(n298) );
  XNOR2_X1 U362 ( .A(n299), .B(n298), .ZN(n301) );
  XNOR2_X1 U363 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n300) );
  XNOR2_X1 U364 ( .A(n300), .B(KEYINPUT2), .ZN(n340) );
  XOR2_X1 U365 ( .A(n301), .B(n340), .Z(n303) );
  XOR2_X1 U366 ( .A(G113GAT), .B(G1GAT), .Z(n420) );
  XOR2_X1 U367 ( .A(G134GAT), .B(KEYINPUT81), .Z(n383) );
  XNOR2_X1 U368 ( .A(n420), .B(n383), .ZN(n302) );
  XNOR2_X1 U369 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U371 ( .A(n307), .B(n306), .ZN(n515) );
  INV_X1 U372 ( .A(n515), .ZN(n566) );
  XOR2_X1 U373 ( .A(KEYINPUT20), .B(G176GAT), .Z(n309) );
  XNOR2_X1 U374 ( .A(G15GAT), .B(G113GAT), .ZN(n308) );
  XNOR2_X1 U375 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U376 ( .A(G43GAT), .B(n310), .ZN(n312) );
  XOR2_X1 U377 ( .A(G190GAT), .B(G134GAT), .Z(n315) );
  XOR2_X1 U378 ( .A(G120GAT), .B(G71GAT), .Z(n439) );
  XNOR2_X1 U379 ( .A(n439), .B(n313), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U381 ( .A(KEYINPUT91), .B(KEYINPUT89), .Z(n319) );
  NAND2_X1 U382 ( .A1(G227GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U384 ( .A(n321), .B(n320), .Z(n327) );
  XNOR2_X1 U385 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n323) );
  XOR2_X1 U386 ( .A(G183GAT), .B(KEYINPUT19), .Z(n324) );
  XNOR2_X1 U387 ( .A(n330), .B(KEYINPUT90), .ZN(n326) );
  XOR2_X1 U388 ( .A(KEYINPUT21), .B(G211GAT), .Z(n329) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(G218GAT), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n348) );
  XNOR2_X1 U391 ( .A(n330), .B(G92GAT), .ZN(n333) );
  XOR2_X1 U392 ( .A(G8GAT), .B(KEYINPUT84), .Z(n396) );
  XOR2_X1 U393 ( .A(G204GAT), .B(n396), .Z(n331) );
  XOR2_X1 U394 ( .A(G176GAT), .B(G64GAT), .Z(n435) );
  AND2_X1 U395 ( .A1(G226GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n348), .B(n336), .ZN(n338) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(G190GAT), .ZN(n337) );
  XOR2_X1 U399 ( .A(n337), .B(KEYINPUT82), .Z(n376) );
  NAND2_X1 U400 ( .A1(n527), .A2(n517), .ZN(n339) );
  XNOR2_X1 U401 ( .A(KEYINPUT98), .B(n339), .ZN(n356) );
  XOR2_X1 U402 ( .A(G141GAT), .B(G22GAT), .Z(n421) );
  XOR2_X1 U403 ( .A(n340), .B(n421), .Z(n342) );
  NAND2_X1 U404 ( .A1(G228GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U406 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n344) );
  XNOR2_X1 U407 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U409 ( .A(n346), .B(n345), .Z(n350) );
  XNOR2_X1 U410 ( .A(G50GAT), .B(KEYINPUT75), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n347), .B(G162GAT), .ZN(n377) );
  XNOR2_X1 U412 ( .A(n377), .B(n348), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n355) );
  XOR2_X1 U414 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n352) );
  XNOR2_X1 U415 ( .A(G78GAT), .B(G148GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U417 ( .A(G106GAT), .B(G204GAT), .Z(n353) );
  XNOR2_X1 U418 ( .A(n354), .B(n353), .ZN(n446) );
  XNOR2_X1 U419 ( .A(n355), .B(n446), .ZN(n468) );
  NAND2_X1 U420 ( .A1(n356), .A2(n468), .ZN(n357) );
  XNOR2_X1 U421 ( .A(KEYINPUT25), .B(n357), .ZN(n362) );
  NOR2_X1 U422 ( .A1(n527), .A2(n468), .ZN(n358) );
  XNOR2_X1 U423 ( .A(KEYINPUT27), .B(KEYINPUT95), .ZN(n359) );
  XOR2_X1 U424 ( .A(n359), .B(n517), .Z(n366) );
  AND2_X1 U425 ( .A1(n568), .A2(n366), .ZN(n360) );
  XOR2_X1 U426 ( .A(n360), .B(KEYINPUT97), .Z(n361) );
  XNOR2_X1 U427 ( .A(n363), .B(KEYINPUT99), .ZN(n364) );
  AND2_X1 U428 ( .A1(n566), .A2(n364), .ZN(n365) );
  XNOR2_X1 U429 ( .A(n365), .B(KEYINPUT100), .ZN(n369) );
  NAND2_X1 U430 ( .A1(n515), .A2(n366), .ZN(n367) );
  XOR2_X1 U431 ( .A(KEYINPUT96), .B(n367), .Z(n542) );
  XNOR2_X1 U432 ( .A(n468), .B(KEYINPUT28), .ZN(n492) );
  NAND2_X1 U433 ( .A1(n542), .A2(n492), .ZN(n529) );
  NOR2_X1 U434 ( .A1(n529), .A2(n527), .ZN(n368) );
  NOR2_X1 U435 ( .A1(n369), .A2(n368), .ZN(n482) );
  XOR2_X1 U436 ( .A(KEYINPUT11), .B(KEYINPUT83), .Z(n371) );
  XNOR2_X1 U437 ( .A(G106GAT), .B(KEYINPUT77), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U439 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n373) );
  XNOR2_X1 U440 ( .A(KEYINPUT66), .B(KEYINPUT10), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U442 ( .A(n375), .B(n374), .Z(n379) );
  XOR2_X1 U443 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U444 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U445 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n381) );
  XNOR2_X1 U446 ( .A(G218GAT), .B(KEYINPUT78), .ZN(n380) );
  XNOR2_X1 U447 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U448 ( .A(n383), .B(n382), .Z(n385) );
  NAND2_X1 U449 ( .A1(G232GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U450 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U451 ( .A(n387), .B(n386), .Z(n393) );
  XOR2_X1 U452 ( .A(G29GAT), .B(G43GAT), .Z(n389) );
  XNOR2_X1 U453 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n389), .B(n388), .ZN(n429) );
  XOR2_X1 U455 ( .A(G85GAT), .B(G92GAT), .Z(n391) );
  XNOR2_X1 U456 ( .A(G99GAT), .B(KEYINPUT73), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n434) );
  XNOR2_X1 U458 ( .A(n429), .B(n434), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n478) );
  XNOR2_X1 U460 ( .A(n478), .B(KEYINPUT36), .ZN(n582) );
  XOR2_X1 U461 ( .A(G78GAT), .B(G64GAT), .Z(n395) );
  XNOR2_X1 U462 ( .A(G22GAT), .B(G1GAT), .ZN(n394) );
  XNOR2_X1 U463 ( .A(n395), .B(n394), .ZN(n397) );
  XOR2_X1 U464 ( .A(n397), .B(n396), .Z(n399) );
  XNOR2_X1 U465 ( .A(G15GAT), .B(G71GAT), .ZN(n398) );
  XNOR2_X1 U466 ( .A(n399), .B(n398), .ZN(n412) );
  XOR2_X1 U467 ( .A(KEYINPUT12), .B(G211GAT), .Z(n401) );
  NAND2_X1 U468 ( .A1(G231GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U469 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U470 ( .A(KEYINPUT13), .B(G57GAT), .Z(n438) );
  XOR2_X1 U471 ( .A(n402), .B(n438), .Z(n410) );
  XOR2_X1 U472 ( .A(KEYINPUT86), .B(KEYINPUT14), .Z(n404) );
  XNOR2_X1 U473 ( .A(KEYINPUT15), .B(KEYINPUT87), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U475 ( .A(KEYINPUT85), .B(G155GAT), .Z(n406) );
  XNOR2_X1 U476 ( .A(G183GAT), .B(G127GAT), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U480 ( .A(n412), .B(n411), .Z(n559) );
  OR2_X1 U481 ( .A1(n582), .A2(n559), .ZN(n413) );
  OR2_X1 U482 ( .A1(n482), .A2(n413), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n514) );
  XOR2_X1 U484 ( .A(G15GAT), .B(KEYINPUT68), .Z(n417) );
  XNOR2_X1 U485 ( .A(G169GAT), .B(KEYINPUT29), .ZN(n416) );
  XOR2_X1 U486 ( .A(n417), .B(n416), .Z(n433) );
  XOR2_X1 U487 ( .A(KEYINPUT67), .B(KEYINPUT69), .Z(n419) );
  XNOR2_X1 U488 ( .A(KEYINPUT70), .B(G8GAT), .ZN(n418) );
  XNOR2_X1 U489 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U490 ( .A(G36GAT), .B(G50GAT), .Z(n423) );
  XNOR2_X1 U491 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U492 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U493 ( .A(n425), .B(n424), .Z(n427) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U496 ( .A(n428), .B(G197GAT), .Z(n431) );
  XNOR2_X1 U497 ( .A(n429), .B(KEYINPUT30), .ZN(n430) );
  XNOR2_X1 U498 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n557) );
  XNOR2_X1 U500 ( .A(n435), .B(n434), .ZN(n437) );
  AND2_X1 U501 ( .A1(G230GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U502 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U503 ( .A(n439), .B(n438), .Z(n443) );
  XOR2_X1 U504 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n441) );
  XNOR2_X1 U505 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n440) );
  XNOR2_X1 U506 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n575) );
  NAND2_X1 U508 ( .A1(n557), .A2(n575), .ZN(n483) );
  NOR2_X1 U509 ( .A1(n514), .A2(n483), .ZN(n448) );
  XNOR2_X1 U510 ( .A(KEYINPUT38), .B(n448), .ZN(n501) );
  NAND2_X1 U511 ( .A1(n501), .A2(n527), .ZN(n450) );
  XNOR2_X1 U512 ( .A(KEYINPUT55), .B(KEYINPUT122), .ZN(n471) );
  XOR2_X1 U513 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n456) );
  XOR2_X1 U514 ( .A(n575), .B(KEYINPUT65), .Z(n451) );
  XNOR2_X1 U515 ( .A(n451), .B(KEYINPUT41), .ZN(n547) );
  AND2_X1 U516 ( .A1(n547), .A2(n557), .ZN(n452) );
  XNOR2_X1 U517 ( .A(n452), .B(KEYINPUT46), .ZN(n454) );
  INV_X1 U518 ( .A(n478), .ZN(n562) );
  OR2_X1 U519 ( .A1(n559), .A2(n562), .ZN(n453) );
  XNOR2_X1 U520 ( .A(n456), .B(n455), .ZN(n462) );
  INV_X1 U521 ( .A(n559), .ZN(n579) );
  NOR2_X1 U522 ( .A1(n579), .A2(n582), .ZN(n457) );
  XNOR2_X1 U523 ( .A(KEYINPUT45), .B(n457), .ZN(n458) );
  NAND2_X1 U524 ( .A1(n458), .A2(n575), .ZN(n459) );
  NOR2_X1 U525 ( .A1(n557), .A2(n459), .ZN(n460) );
  XNOR2_X1 U526 ( .A(n460), .B(KEYINPUT112), .ZN(n461) );
  NOR2_X1 U527 ( .A1(n462), .A2(n461), .ZN(n465) );
  INV_X1 U528 ( .A(KEYINPUT48), .ZN(n463) );
  NAND2_X1 U529 ( .A1(n517), .A2(n526), .ZN(n467) );
  XOR2_X1 U530 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n466) );
  XOR2_X1 U531 ( .A(n467), .B(n466), .Z(n567) );
  AND2_X1 U532 ( .A1(n468), .A2(n566), .ZN(n469) );
  NAND2_X1 U533 ( .A1(n567), .A2(n469), .ZN(n470) );
  XNOR2_X1 U534 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n472), .A2(n527), .ZN(n473) );
  NAND2_X1 U536 ( .A1(n563), .A2(n547), .ZN(n477) );
  XOR2_X1 U537 ( .A(G176GAT), .B(KEYINPUT56), .Z(n475) );
  XNOR2_X1 U538 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n474) );
  NAND2_X1 U539 ( .A1(n559), .A2(n478), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n479), .B(KEYINPUT16), .ZN(n480) );
  XNOR2_X1 U541 ( .A(n480), .B(KEYINPUT88), .ZN(n481) );
  NOR2_X1 U542 ( .A1(n483), .A2(n504), .ZN(n493) );
  NAND2_X1 U543 ( .A1(n515), .A2(n493), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n485) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U548 ( .A1(n517), .A2(n493), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT103), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U551 ( .A1(n493), .A2(n527), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U553 ( .A(G15GAT), .B(n491), .Z(G1326GAT) );
  INV_X1 U554 ( .A(n492), .ZN(n520) );
  NAND2_X1 U555 ( .A1(n493), .A2(n520), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(KEYINPUT104), .ZN(n495) );
  XNOR2_X1 U557 ( .A(G22GAT), .B(n495), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n497) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n499) );
  NAND2_X1 U561 ( .A1(n501), .A2(n515), .ZN(n498) );
  XOR2_X1 U562 ( .A(n499), .B(n498), .Z(G1328GAT) );
  NAND2_X1 U563 ( .A1(n501), .A2(n517), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n501), .A2(n520), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U567 ( .A(n557), .ZN(n570) );
  NAND2_X1 U568 ( .A1(n547), .A2(n570), .ZN(n503) );
  XOR2_X1 U569 ( .A(n503), .B(KEYINPUT107), .Z(n513) );
  OR2_X1 U570 ( .A1(n513), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(KEYINPUT42), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G57GAT), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n517), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U575 ( .A1(n510), .A2(n527), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U578 ( .A1(n520), .A2(n510), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n521), .A2(n515), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n521), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n527), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n525) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U589 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n537), .A2(n557), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n533) );
  NAND2_X1 U598 ( .A1(n537), .A2(n547), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  NAND2_X1 U601 ( .A1(n537), .A2(n559), .ZN(n535) );
  XNOR2_X1 U602 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U605 ( .A1(n537), .A2(n562), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT115), .Z(n540) );
  XNOR2_X1 U608 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  XOR2_X1 U609 ( .A(G141GAT), .B(KEYINPUT117), .Z(n546) );
  NAND2_X1 U610 ( .A1(n526), .A2(n542), .ZN(n543) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n555), .A2(n557), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n551) );
  XOR2_X1 U615 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n549) );
  NAND2_X1 U616 ( .A1(n555), .A2(n547), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1345GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n553) );
  NAND2_X1 U620 ( .A1(n555), .A2(n559), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n562), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n563), .A2(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(G183GAT), .B(KEYINPUT125), .Z(n561) );
  NAND2_X1 U628 ( .A1(n563), .A2(n559), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(G1350GAT) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  AND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n581) );
  NOR2_X1 U635 ( .A1(n570), .A2(n581), .ZN(n574) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT60), .ZN(n572) );
  XNOR2_X1 U638 ( .A(KEYINPUT126), .B(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U640 ( .A1(n575), .A2(n581), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT127), .B(KEYINPUT61), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XOR2_X1 U645 ( .A(G211GAT), .B(n580), .Z(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

