//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n603, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AND4_X1   g045(.A1(new_n463), .A2(new_n466), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n462), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n466), .A2(new_n468), .A3(new_n470), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n466), .A2(new_n468), .A3(new_n470), .A4(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(KEYINPUT69), .A3(new_n462), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n464), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  OR2_X1    g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n480), .A2(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n464), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n482), .A2(G112), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n464), .A2(new_n482), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n490), .B1(G136), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT70), .ZN(G162));
  AND2_X1   g069(.A1(KEYINPUT71), .A2(G138), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n468), .A2(new_n470), .A3(new_n495), .A4(new_n482), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n464), .A2(KEYINPUT4), .A3(new_n482), .A4(new_n495), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n468), .A2(new_n470), .A3(G126), .A4(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n502), .A2(new_n504), .A3(G2104), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n500), .A2(new_n506), .ZN(G164));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n514), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n527));
  INV_X1    g102(.A(new_n510), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n514), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n529), .B1(new_n535), .B2(G51), .ZN(G168));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n539), .A2(new_n512), .B1(new_n540), .B2(new_n515), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n535), .A2(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  INV_X1    g119(.A(G56), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n528), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n510), .A2(new_n514), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n546), .A2(G651), .B1(new_n547), .B2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT74), .ZN(G188));
  NAND2_X1  g132(.A1(new_n530), .A2(G53), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n547), .A2(G91), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(new_n512), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT75), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  OR2_X1    g144(.A1(new_n538), .A2(new_n541), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n547), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n530), .A2(G49), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n508), .B2(new_n509), .ZN(new_n577));
  AND2_X1   g152(.A1(G73), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n510), .A2(new_n514), .A3(G86), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G305));
  XNOR2_X1  g157(.A(KEYINPUT76), .B(G47), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n534), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI22_X1  g161(.A1(new_n585), .A2(new_n512), .B1(new_n586), .B2(new_n515), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(new_n535), .A2(G54), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n547), .A2(G92), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT10), .Z(new_n592));
  AOI22_X1  g167(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n512), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n590), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G171), .B2(new_n596), .ZN(G284));
  OAI21_X1  g173(.A(new_n597), .B1(G171), .B2(new_n596), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n568), .B2(G868), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(new_n568), .B2(G868), .ZN(G280));
  INV_X1    g177(.A(new_n595), .ZN(new_n603));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n492), .A2(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  OR2_X1    g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n614), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n615));
  INV_X1    g190(.A(G135), .ZN(new_n616));
  INV_X1    g191(.A(G123), .ZN(new_n617));
  OAI221_X1 g192(.A(new_n615), .B1(new_n491), .B2(new_n616), .C1(new_n617), .C2(new_n485), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT77), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2096), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n613), .A2(new_n620), .ZN(G156));
  XOR2_X1   g196(.A(G1341), .B(G1348), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT79), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT16), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n623), .B(new_n625), .Z(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT78), .B(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n626), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n634), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT80), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT81), .B(KEYINPUT17), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n639), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n643), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n642), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n640), .A3(new_n639), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND2_X1  g225(.A1(new_n641), .A2(new_n639), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n650), .C1(new_n645), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2096), .B(G2100), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(G227));
  XOR2_X1   g229(.A(G1971), .B(G1976), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1956), .B(G2474), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1961), .B(G1966), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n656), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n659), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT20), .Z(new_n663));
  AOI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n656), .C2(new_n660), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT82), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT83), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(G229));
  INV_X1    g249(.A(G29), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G26), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT88), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  AOI22_X1  g253(.A1(G128), .A2(new_n486), .B1(new_n492), .B2(G140), .ZN(new_n679));
  OAI21_X1  g254(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G116), .B2(new_n482), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT87), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n678), .B1(new_n684), .B2(new_n675), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2067), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT25), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n464), .A2(G127), .ZN(new_n689));
  NAND2_X1  g264(.A1(G115), .A2(G2104), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n482), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AOI211_X1 g266(.A(new_n688), .B(new_n691), .C1(G139), .C2(new_n492), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n692), .A2(new_n675), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n675), .B2(G33), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(G2072), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(G2072), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n618), .A2(new_n675), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT30), .B(G28), .ZN(new_n699));
  OR2_X1    g274(.A1(KEYINPUT31), .A2(G11), .ZN(new_n700));
  NAND2_X1  g275(.A1(KEYINPUT31), .A2(G11), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n699), .A2(new_n675), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n696), .A2(new_n697), .A3(new_n698), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G164), .A2(new_n675), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G27), .B2(new_n675), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n686), .B(new_n703), .C1(G2078), .C2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G19), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n550), .B2(G16), .ZN(new_n709));
  OAI22_X1  g284(.A1(new_n709), .A2(G1341), .B1(G2078), .B2(new_n706), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n492), .A2(G141), .B1(G105), .B2(new_n460), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT26), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(new_n486), .B2(G129), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(new_n675), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT92), .B1(G29), .B2(G32), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(new_n716), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n710), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NOR2_X1   g299(.A1(G171), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G5), .B2(new_n724), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n727), .A2(G1961), .B1(new_n721), .B2(new_n720), .ZN(new_n728));
  INV_X1    g303(.A(G1961), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n726), .A2(new_n729), .B1(new_n709), .B2(G1341), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n707), .A2(new_n723), .A3(new_n728), .A4(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G160), .A2(G29), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n675), .B1(new_n733), .B2(G34), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT89), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(new_n733), .B2(G34), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(new_n734), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT90), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT91), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n731), .B1(G2084), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n724), .A2(G23), .ZN(new_n743));
  INV_X1    g318(.A(G288), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n724), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT33), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1976), .ZN(new_n747));
  MUX2_X1   g322(.A(G6), .B(G305), .S(G16), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT85), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT32), .B(G1981), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G22), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G166), .B2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1971), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n747), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT34), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT34), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n724), .A2(G24), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n588), .B2(new_n724), .ZN(new_n760));
  INV_X1    g335(.A(G1986), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n492), .A2(G131), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n486), .A2(G119), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n482), .A2(G107), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT84), .ZN(new_n768));
  MUX2_X1   g343(.A(G25), .B(new_n768), .S(G29), .Z(new_n769));
  XOR2_X1   g344(.A(KEYINPUT35), .B(G1991), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n757), .A2(new_n758), .A3(new_n762), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT36), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n741), .A2(G2084), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT94), .Z(new_n775));
  NOR2_X1   g350(.A1(G29), .A2(G35), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G162), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT29), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2090), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n603), .B2(G16), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT86), .B(G1348), .Z(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(G168), .A2(G16), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n784), .A2(KEYINPUT93), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT93), .B1(G16), .B2(G21), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n785), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n789), .A2(G1966), .B1(new_n781), .B2(new_n782), .ZN(new_n790));
  INV_X1    g365(.A(G1966), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n779), .A2(new_n783), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n724), .A2(G20), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT23), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n568), .B2(new_n724), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n778), .A2(G2090), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n793), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n742), .A2(new_n773), .A3(new_n775), .A4(new_n800), .ZN(G150));
  INV_X1    g376(.A(G150), .ZN(G311));
  NAND2_X1  g377(.A1(new_n603), .A2(G559), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT38), .ZN(new_n804));
  INV_X1    g379(.A(G55), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n534), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n807), .A2(new_n512), .B1(new_n808), .B2(new_n515), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n550), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(new_n549), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n804), .B(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n810), .A2(new_n818), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(G162), .B(new_n618), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G160), .Z(new_n825));
  NAND3_X1  g400(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT96), .ZN(new_n826));
  AOI21_X1  g401(.A(KEYINPUT97), .B1(new_n501), .B2(new_n505), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n501), .A2(KEYINPUT97), .A3(new_n505), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT96), .B1(new_n498), .B2(new_n499), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n684), .ZN(new_n834));
  INV_X1    g409(.A(G130), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT98), .B1(new_n482), .B2(G118), .ZN(new_n836));
  OR2_X1    g411(.A1(G106), .A2(G2105), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(G2104), .A3(new_n837), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n482), .A2(KEYINPUT98), .A3(G118), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n485), .A2(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G142), .B2(new_n492), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n834), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n692), .B(new_n715), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n611), .B(new_n767), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n842), .B(new_n845), .ZN(new_n846));
  AOI21_X1  g421(.A(G37), .B1(new_n825), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n825), .B2(new_n846), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g424(.A1(new_n812), .A2(new_n596), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n814), .B(new_n606), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n568), .A2(KEYINPUT99), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n564), .A2(new_n567), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n595), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n568), .A2(KEYINPUT99), .A3(new_n603), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n855), .A2(new_n856), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n855), .A2(KEYINPUT41), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n858), .B1(new_n851), .B2(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(G305), .B(KEYINPUT100), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n588), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G303), .B(new_n744), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n866), .B(new_n867), .Z(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT42), .Z(new_n869));
  XNOR2_X1  g444(.A(new_n864), .B(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n850), .B1(new_n870), .B2(new_n596), .ZN(G295));
  OAI21_X1  g446(.A(new_n850), .B1(new_n870), .B2(new_n596), .ZN(G331));
  INV_X1    g447(.A(KEYINPUT105), .ZN(new_n873));
  NAND2_X1  g448(.A1(G301), .A2(KEYINPUT101), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n538), .A2(KEYINPUT101), .A3(new_n541), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n874), .A2(G168), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(G168), .B1(new_n874), .B2(new_n875), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n815), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n814), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n862), .A3(new_n861), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g459(.A(KEYINPUT102), .B(new_n814), .C1(new_n876), .C2(new_n877), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n857), .A3(new_n879), .A4(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n868), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n857), .A2(new_n879), .A3(new_n880), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n861), .A2(new_n862), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n879), .A3(new_n885), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n894), .B2(new_n887), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n857), .A2(new_n879), .A3(new_n880), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n884), .A2(new_n879), .A3(new_n885), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n896), .B1(new_n897), .B2(new_n863), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n899), .A3(new_n868), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n890), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n873), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n890), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n893), .A2(new_n862), .A3(new_n861), .ZN(new_n905));
  AOI211_X1 g480(.A(KEYINPUT104), .B(new_n887), .C1(new_n905), .C2(new_n896), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n899), .B1(new_n898), .B2(new_n868), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n868), .A2(KEYINPUT103), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n882), .A2(new_n886), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n882), .B2(new_n886), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n912), .A2(new_n913), .A3(G37), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n910), .B1(new_n914), .B2(new_n902), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n903), .A2(new_n909), .A3(new_n915), .ZN(new_n916));
  AOI211_X1 g491(.A(KEYINPUT43), .B(new_n890), .C1(new_n895), .C2(new_n900), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n914), .A2(new_n902), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(G397));
  AOI21_X1  g495(.A(KEYINPUT69), .B1(new_n478), .B2(new_n462), .ZN(new_n921));
  AOI211_X1 g496(.A(new_n473), .B(new_n461), .C1(new_n476), .C2(new_n477), .ZN(new_n922));
  OAI211_X1 g497(.A(G40), .B(new_n483), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n480), .A2(KEYINPUT106), .A3(G40), .A4(new_n483), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n829), .B2(new_n831), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G2067), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n684), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT108), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n711), .B2(new_n714), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n932), .A2(new_n937), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(new_n715), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT107), .ZN(new_n942));
  INV_X1    g517(.A(new_n770), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n767), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n932), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n939), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n588), .B(new_n761), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n932), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n563), .B(KEYINPUT57), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n928), .B1(new_n500), .B2(new_n506), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n930), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(KEYINPUT45), .B(new_n928), .C1(new_n829), .C2(new_n831), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n950), .A2(KEYINPUT109), .A3(new_n930), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n927), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g532(.A(KEYINPUT56), .B(G2072), .Z(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(KEYINPUT122), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT122), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n950), .A2(KEYINPUT109), .A3(new_n930), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT109), .B1(new_n950), .B2(new_n930), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n964), .A2(new_n925), .A3(new_n926), .A4(new_n954), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n965), .B2(new_n958), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n927), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n950), .A2(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n929), .B2(KEYINPUT50), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  XOR2_X1   g546(.A(KEYINPUT121), .B(G1956), .Z(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n949), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT123), .ZN(new_n975));
  INV_X1    g550(.A(new_n929), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n925), .A2(new_n926), .A3(new_n976), .ZN(new_n977));
  OR2_X1    g552(.A1(new_n977), .A2(G2067), .ZN(new_n978));
  INV_X1    g553(.A(G1348), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n980), .B(new_n928), .C1(new_n829), .C2(new_n831), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n950), .A2(KEYINPUT50), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n979), .B1(new_n927), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n975), .B1(new_n978), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n978), .A2(new_n975), .A3(new_n984), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(new_n595), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n967), .A2(new_n949), .A3(new_n973), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n974), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n974), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(KEYINPUT61), .A3(new_n990), .ZN(new_n993));
  INV_X1    g568(.A(new_n987), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT60), .B1(new_n994), .B2(new_n985), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT60), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n986), .A2(new_n996), .A3(new_n987), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n997), .A3(new_n603), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n988), .A2(KEYINPUT60), .A3(new_n595), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT61), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n967), .A2(new_n949), .A3(new_n973), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n974), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT58), .B(G1341), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n977), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1005), .B1(G1996), .B2(new_n965), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n550), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT124), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT124), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1009), .A3(new_n550), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1008), .A2(KEYINPUT59), .A3(new_n1010), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1003), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n991), .B1(new_n1000), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n729), .B1(new_n927), .B2(new_n983), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n950), .A2(new_n930), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  AOI211_X1 g595(.A(new_n1020), .B(G2078), .C1(new_n929), .C2(new_n930), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n968), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1023), .A2(KEYINPUT110), .A3(new_n925), .A4(new_n926), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT110), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1025), .B1(new_n927), .B2(new_n956), .ZN(new_n1026));
  AOI21_X1  g601(.A(G2078), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1018), .B(new_n1022), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT126), .B1(new_n1030), .B2(G301), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT126), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1032), .A3(G171), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1021), .A2(G40), .A3(G160), .A4(new_n954), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1018), .B(new_n1035), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G171), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1017), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT112), .B(G8), .Z(new_n1039));
  NOR2_X1   g614(.A1(G168), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1040), .A2(KEYINPUT51), .ZN(new_n1041));
  AND4_X1   g616(.A1(new_n925), .A2(new_n926), .A3(new_n981), .A4(new_n982), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT118), .B(G2084), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n925), .A2(new_n931), .A3(new_n926), .A4(new_n1019), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1042), .A2(new_n1043), .B1(new_n1044), .B2(new_n791), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1041), .B1(new_n1045), .B2(new_n1039), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1044), .A2(new_n791), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1040), .B1(new_n1049), .B2(G8), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1049), .A2(new_n1040), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1024), .A2(new_n1026), .A3(new_n754), .ZN(new_n1055));
  INV_X1    g630(.A(G2090), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n968), .A2(new_n1056), .A3(new_n970), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1039), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G303), .A2(G8), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT111), .B(KEYINPUT55), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1042), .A2(new_n1056), .ZN(new_n1065));
  AOI211_X1 g640(.A(new_n1064), .B(new_n1061), .C1(new_n1055), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1039), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G288), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT113), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n977), .A2(new_n1067), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(KEYINPUT49), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G305), .A2(G1981), .ZN(new_n1079));
  INV_X1    g654(.A(G1981), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n579), .A2(new_n1080), .A3(new_n580), .A4(new_n581), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1077), .A2(KEYINPUT49), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1077), .B(KEYINPUT49), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n977), .A3(new_n1067), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n977), .A2(new_n1090), .A3(new_n1067), .A4(new_n1071), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1075), .A2(new_n1076), .A3(new_n1087), .A4(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1066), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1054), .A2(new_n1063), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT54), .B1(new_n1029), .B2(G171), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1036), .A2(KEYINPUT127), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1036), .B2(KEYINPUT127), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1094), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1016), .A2(new_n1038), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1054), .B(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1102), .A2(new_n1063), .A3(new_n1093), .A4(new_n1034), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1087), .A2(new_n1068), .A3(new_n744), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1081), .B(KEYINPUT117), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1067), .A3(new_n977), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1055), .A2(new_n1065), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(G8), .A3(new_n1062), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1109), .B2(new_n1092), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1072), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT114), .B1(new_n1072), .B2(KEYINPUT52), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1091), .A2(new_n1087), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1109), .B(new_n1115), .C1(new_n1058), .C2(new_n1062), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1045), .A2(G286), .A3(new_n1039), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1111), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1093), .A2(new_n1063), .A3(KEYINPUT119), .A4(new_n1117), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1108), .A2(G8), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1061), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1093), .A2(KEYINPUT63), .A3(new_n1117), .A4(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1110), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1100), .B(new_n1103), .C1(new_n1126), .C2(KEYINPUT120), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1128), .B(new_n1110), .C1(new_n1122), .C2(new_n1125), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n948), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n940), .A2(KEYINPUT46), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n940), .A2(KEYINPUT46), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n934), .A2(new_n715), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1131), .A2(new_n1132), .B1(new_n932), .B2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(new_n1134), .B(KEYINPUT47), .Z(new_n1135));
  NAND3_X1  g710(.A1(new_n932), .A2(new_n761), .A3(new_n588), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT48), .Z(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n946), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n768), .A2(new_n943), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n939), .A2(new_n942), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n684), .A2(new_n933), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n932), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1130), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g719(.A(G319), .ZN(new_n1146));
  NOR4_X1   g720(.A1(G229), .A2(new_n1146), .A3(G401), .A4(G227), .ZN(new_n1147));
  OAI211_X1 g721(.A(new_n848), .B(new_n1147), .C1(new_n917), .C2(new_n918), .ZN(G225));
  INV_X1    g722(.A(G225), .ZN(G308));
endmodule


