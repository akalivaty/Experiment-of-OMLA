//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G113), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT2), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G113), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G116), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT2), .B(G113), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n199), .A2(new_n200), .A3(KEYINPUT68), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n202), .B1(new_n191), .B2(new_n192), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n194), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT70), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT68), .B1(new_n199), .B2(new_n200), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n191), .A2(new_n192), .A3(new_n202), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT70), .A3(new_n194), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  AOI22_X1  g027(.A1(KEYINPUT66), .A2(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  OAI22_X1  g028(.A1(KEYINPUT66), .A2(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT11), .A4(G134), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n218), .A2(G134), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n213), .A2(G137), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(KEYINPUT65), .A2(G143), .ZN(new_n224));
  NOR2_X1   g038(.A1(KEYINPUT65), .A2(G143), .ZN(new_n225));
  OAI21_X1  g039(.A(G146), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n226), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n227), .ZN(new_n234));
  INV_X1    g048(.A(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT65), .A2(G143), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n235), .A2(G143), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT67), .B(G128), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT1), .B1(new_n227), .B2(G146), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n237), .A2(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n220), .B(new_n223), .C1(new_n232), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n247), .B1(new_n237), .B2(new_n239), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT0), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n230), .A3(KEYINPUT64), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(KEYINPUT0), .B2(G128), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n234), .A2(new_n236), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n228), .B1(new_n254), .B2(G146), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n248), .A2(new_n253), .B1(new_n255), .B2(new_n247), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G131), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n220), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n240), .A2(new_n241), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n224), .A2(new_n225), .A3(G146), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(new_n238), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n226), .A2(new_n229), .A3(new_n231), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n265), .A2(KEYINPUT69), .A3(new_n220), .A4(new_n223), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n211), .A2(new_n245), .A3(new_n260), .A4(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G237), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G210), .ZN(new_n270));
  INV_X1    g084(.A(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n272), .B(new_n273), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n260), .A2(new_n276), .A3(new_n243), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n245), .A2(new_n266), .A3(new_n260), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(KEYINPUT30), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n204), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n267), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n205), .B(new_n193), .C1(new_n208), .C2(new_n207), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n209), .B2(new_n194), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n258), .A2(new_n220), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n255), .A2(new_n247), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n246), .B(new_n253), .C1(new_n262), .C2(new_n238), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n243), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n282), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n204), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n291), .B(new_n292), .C1(new_n267), .C2(new_n282), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n274), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n281), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT72), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n300), .A3(new_n296), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n291), .B(KEYINPUT73), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n278), .A2(new_n285), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n267), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT28), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n303), .A2(KEYINPUT29), .A3(new_n274), .A4(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT74), .ZN(new_n308));
  OAI21_X1  g122(.A(G472), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n267), .B(new_n274), .C1(new_n279), .C2(new_n280), .ZN(new_n310));
  OAI21_X1  g124(.A(KEYINPUT71), .B1(new_n310), .B2(KEYINPUT31), .ZN(new_n311));
  INV_X1    g125(.A(new_n267), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n278), .A2(KEYINPUT30), .ZN(new_n313));
  INV_X1    g127(.A(new_n277), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n315), .B2(new_n204), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT31), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .A4(new_n274), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n310), .A2(KEYINPUT31), .B1(new_n275), .B2(new_n293), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(G472), .A2(G902), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT32), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(new_n323), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(new_n320), .B2(new_n321), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT32), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n309), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n224), .A2(new_n225), .ZN(new_n331));
  OAI22_X1  g145(.A1(new_n331), .A2(new_n230), .B1(new_n240), .B2(new_n227), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(G134), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n197), .A2(KEYINPUT14), .A3(G122), .ZN(new_n334));
  XNOR2_X1  g148(.A(G116), .B(G122), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(G107), .B(new_n334), .C1(new_n336), .C2(KEYINPUT14), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n333), .B(new_n337), .C1(G107), .C2(new_n336), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT67), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G128), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT13), .B1(new_n343), .B2(G143), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n332), .B1(new_n344), .B2(new_n213), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n254), .A2(G128), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(G143), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT13), .A4(G134), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n335), .B(G107), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n339), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  AOI211_X1 g166(.A(KEYINPUT92), .B(new_n350), .C1(new_n345), .C2(new_n348), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n338), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT9), .B(G234), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n356), .A2(new_n357), .A3(G953), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n338), .B(new_n358), .C1(new_n352), .C2(new_n353), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(KEYINPUT93), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT93), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n354), .A2(new_n363), .A3(new_n359), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(new_n299), .A3(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n365), .A2(KEYINPUT94), .ZN(new_n366));
  INV_X1    g180(.A(G478), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n367), .A2(KEYINPUT15), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n365), .B2(KEYINPUT94), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n366), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n196), .A2(KEYINPUT5), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT85), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n187), .B1(new_n192), .B2(KEYINPUT5), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT3), .B1(new_n377), .B2(G107), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G104), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(G107), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n378), .A2(new_n381), .A3(new_n271), .A4(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n377), .A2(G107), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n380), .A2(G104), .ZN(new_n385));
  OAI21_X1  g199(.A(G101), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT81), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n383), .B2(new_n386), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n376), .B(new_n209), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n378), .A2(new_n381), .A3(new_n382), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(G101), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT4), .A3(new_n383), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n204), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g212(.A(G110), .B(G122), .Z(new_n399));
  OR2_X1    g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n289), .A2(G125), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(G125), .B2(new_n265), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n269), .A2(G224), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n398), .A2(new_n407), .A3(new_n399), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT7), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n404), .A2(new_n410), .A3(new_n405), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n376), .A2(new_n209), .ZN(new_n412));
  INV_X1    g226(.A(new_n387), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n391), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n399), .B(KEYINPUT8), .Z(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n404), .B1(new_n410), .B2(new_n405), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n400), .A2(new_n411), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n409), .A2(new_n299), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  XOR2_X1   g234(.A(new_n420), .B(KEYINPUT86), .Z(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(G234), .A2(G237), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(G952), .A3(new_n269), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT21), .B(G898), .Z(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(G902), .A3(G953), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n409), .A2(new_n299), .A3(new_n421), .A4(new_n418), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n423), .A2(new_n428), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n268), .A2(new_n269), .A3(G214), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n254), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n227), .A2(new_n268), .A3(new_n269), .A4(G214), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n254), .B2(KEYINPUT87), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n216), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n432), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n331), .B2(KEYINPUT87), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n432), .B(new_n227), .C1(KEYINPUT65), .C2(new_n433), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(G131), .A3(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT17), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n437), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT91), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G140), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(G125), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT16), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT79), .B1(new_n446), .B2(G125), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT79), .ZN(new_n451));
  INV_X1    g265(.A(G125), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(G140), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n450), .A2(new_n453), .B1(G125), .B2(new_n446), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n449), .B1(new_n454), .B2(new_n448), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n235), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n441), .A2(new_n442), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT91), .A4(new_n442), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n445), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(G113), .B(G122), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(new_n377), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n452), .A2(G140), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n447), .A2(new_n462), .A3(new_n235), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n454), .B2(new_n235), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n439), .A2(new_n440), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT18), .A2(G131), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n467), .B(KEYINPUT89), .Z(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(KEYINPUT88), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT88), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n439), .A2(new_n471), .A3(new_n440), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n465), .B(new_n469), .C1(new_n473), .C2(new_n467), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n459), .A2(new_n461), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n461), .B1(new_n459), .B2(new_n474), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n299), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G475), .ZN(new_n478));
  INV_X1    g292(.A(G475), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n437), .A2(new_n441), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n455), .A2(G146), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT19), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n447), .A2(new_n462), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n454), .B2(new_n484), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n486), .A2(G146), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n437), .A2(new_n441), .A3(KEYINPUT90), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n482), .A2(new_n483), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n461), .B1(new_n489), .B2(new_n474), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n479), .B(new_n299), .C1(new_n475), .C2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT20), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n474), .ZN(new_n494));
  INV_X1    g308(.A(new_n461), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n459), .A2(new_n461), .A3(new_n474), .ZN(new_n497));
  AOI21_X1  g311(.A(G475), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n493), .B1(new_n498), .B2(new_n299), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n478), .B1(new_n492), .B2(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n372), .A2(new_n431), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n357), .B1(G234), .B2(new_n299), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n195), .A2(G128), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT76), .ZN(new_n504));
  OR3_X1    g318(.A1(new_n240), .A2(KEYINPUT75), .A3(new_n195), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n343), .A2(G119), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT75), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT24), .B(G110), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT77), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT23), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n511), .A2(KEYINPUT78), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(KEYINPUT78), .ZN(new_n513));
  OAI22_X1  g327(.A1(new_n512), .A2(new_n513), .B1(new_n195), .B2(G128), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n514), .B(new_n503), .C1(new_n506), .C2(new_n511), .ZN(new_n515));
  OAI22_X1  g329(.A1(new_n508), .A2(new_n510), .B1(new_n515), .B2(G110), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n464), .A3(new_n483), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n455), .B(G146), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n508), .A2(new_n510), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n515), .A2(G110), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT22), .B(G137), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n523), .B(new_n524), .Z(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n517), .A2(new_n521), .A3(new_n525), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n299), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n502), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G221), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n355), .B2(new_n299), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n527), .A2(new_n528), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n502), .A2(G902), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n533), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT80), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n230), .B1(new_n237), .B2(KEYINPUT1), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n255), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n226), .A2(new_n229), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT1), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n331), .B2(new_n235), .ZN(new_n547));
  OAI211_X1 g361(.A(KEYINPUT80), .B(new_n545), .C1(new_n547), .C2(new_n230), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n548), .A3(new_n264), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n388), .A2(new_n390), .ZN(new_n550));
  INV_X1    g364(.A(new_n265), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n413), .A2(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n541), .B1(new_n552), .B2(new_n286), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n413), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT10), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n265), .B(KEYINPUT10), .C1(new_n388), .C2(new_n390), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n256), .A2(new_n394), .A3(new_n396), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n560), .A2(new_n563), .A3(new_n286), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT83), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  INV_X1    g380(.A(G227), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n566), .B(new_n568), .Z(new_n569));
  AND3_X1   g383(.A1(new_n564), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n565), .B1(new_n564), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n558), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT84), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT10), .B1(new_n549), .B2(new_n413), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n561), .A2(new_n562), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n259), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n564), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n569), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g394(.A(KEYINPUT84), .B(new_n558), .C1(new_n570), .C2(new_n571), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n574), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G469), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n583), .A3(new_n299), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n583), .A2(new_n299), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n564), .A2(new_n577), .A3(new_n569), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n558), .A2(new_n564), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT82), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n569), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n558), .A2(KEYINPUT82), .A3(new_n564), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n585), .B1(new_n591), .B2(G469), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n540), .B1(new_n584), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n330), .A2(new_n501), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  NAND2_X1  g409(.A1(new_n322), .A2(new_n299), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n328), .B1(new_n596), .B2(G472), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n593), .A2(new_n600), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n361), .A2(KEYINPUT97), .ZN(new_n602));
  INV_X1    g416(.A(new_n348), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT13), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n240), .B2(new_n227), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n605), .A2(G134), .B1(new_n347), .B2(new_n346), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n351), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT92), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n349), .A2(new_n339), .A3(new_n351), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n338), .A4(new_n358), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n602), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n360), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n354), .A2(KEYINPUT96), .A3(new_n359), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n613), .A2(KEYINPUT33), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n362), .A2(new_n618), .A3(new_n364), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n367), .A2(G902), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n365), .A2(new_n367), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n500), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n624), .A2(new_n431), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n599), .A2(new_n601), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  INV_X1    g442(.A(new_n500), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n372), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n431), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n599), .A2(new_n601), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  XNOR2_X1  g448(.A(new_n529), .B(new_n530), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n522), .B(new_n636), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n635), .A2(new_n502), .B1(new_n538), .B2(new_n637), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n535), .B(new_n638), .C1(new_n584), .C2(new_n592), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n501), .A3(new_n597), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT98), .B(KEYINPUT37), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G110), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n640), .B(new_n642), .ZN(G12));
  NAND3_X1  g457(.A1(new_n423), .A2(new_n429), .A3(new_n430), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n427), .A2(G900), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n425), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n630), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n639), .A2(new_n330), .A3(new_n645), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  AOI21_X1  g465(.A(new_n535), .B1(new_n584), .B2(new_n592), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n647), .B(KEYINPUT39), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g468(.A(new_n500), .B(new_n372), .C1(new_n654), .C2(KEYINPUT40), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n423), .A2(new_n430), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT38), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n316), .A2(new_n275), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n305), .A2(new_n274), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n299), .B1(new_n662), .B2(KEYINPUT99), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n665), .A2(new_n326), .A3(new_n329), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n659), .A2(new_n429), .A3(new_n638), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n331), .ZN(G45));
  INV_X1    g482(.A(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n491), .A2(KEYINPUT20), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n498), .A2(new_n493), .A3(new_n299), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n478), .A2(new_n672), .B1(new_n621), .B2(new_n622), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n669), .B1(new_n673), .B2(new_n647), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n669), .A2(new_n500), .A3(new_n623), .A4(new_n647), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(new_n639), .A3(new_n645), .A4(new_n330), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  NAND2_X1  g492(.A1(KEYINPUT101), .A2(G469), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n582), .A2(new_n299), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n679), .B1(new_n582), .B2(new_n299), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n680), .A2(new_n681), .A3(new_n535), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n533), .A2(new_n539), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n682), .A2(new_n330), .A3(new_n684), .A4(new_n625), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  AND4_X1   g501(.A1(new_n330), .A2(new_n682), .A3(new_n684), .A4(new_n631), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n197), .ZN(G18));
  INV_X1    g503(.A(new_n638), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n682), .A2(new_n330), .A3(new_n501), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n365), .A2(KEYINPUT94), .A3(new_n368), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n365), .A2(KEYINPUT94), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n369), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n365), .A2(KEYINPUT94), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n693), .B1(new_n698), .B2(new_n629), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n372), .A2(KEYINPUT104), .A3(new_n500), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n431), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n310), .A2(KEYINPUT31), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n303), .A2(new_n306), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n275), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n320), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n323), .B(KEYINPUT102), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n596), .A2(G472), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(KEYINPUT103), .B1(new_n707), .B2(new_n684), .ZN(new_n708));
  AOI21_X1  g522(.A(G902), .B1(new_n320), .B2(new_n321), .ZN(new_n709));
  INV_X1    g523(.A(G472), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n706), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n311), .A2(new_n319), .B1(new_n275), .B2(new_n703), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n712), .B1(new_n713), .B2(new_n702), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n711), .A2(new_n714), .A3(new_n683), .A4(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n682), .B(new_n701), .C1(new_n708), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n705), .A2(new_n706), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n710), .B2(new_n709), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n715), .B1(new_n721), .B2(new_n683), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n707), .A2(KEYINPUT103), .A3(new_n684), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(KEYINPUT105), .A3(new_n682), .A4(new_n701), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(G122), .Z(G24));
  NOR3_X1   g541(.A1(new_n711), .A2(new_n714), .A3(new_n638), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n676), .A2(new_n682), .A3(new_n645), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  INV_X1    g545(.A(new_n674), .ZN(new_n732));
  INV_X1    g546(.A(new_n675), .ZN(new_n733));
  INV_X1    g547(.A(new_n429), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n734), .B1(new_n423), .B2(new_n430), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n330), .A2(new_n593), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n735), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n674), .A2(new_n675), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(KEYINPUT42), .A3(new_n330), .A4(new_n593), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n744), .B1(new_n630), .B2(new_n648), .ZN(new_n745));
  AND4_X1   g559(.A1(new_n330), .A2(new_n745), .A3(new_n684), .A4(new_n735), .ZN(new_n746));
  INV_X1    g560(.A(new_n652), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(KEYINPUT106), .B2(new_n649), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  OR2_X1    g564(.A1(new_n591), .A2(KEYINPUT45), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n591), .A2(KEYINPUT45), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(G469), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n585), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT46), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT107), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n755), .A2(new_n760), .A3(new_n756), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n584), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n762), .A2(new_n536), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n653), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT108), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n766), .A3(new_n653), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT43), .B1(new_n629), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n629), .A2(new_n623), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI211_X1 g585(.A(new_n771), .B(new_n690), .C1(new_n328), .C2(new_n711), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT44), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n735), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n765), .A2(new_n767), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  INV_X1    g590(.A(KEYINPUT47), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n762), .A2(new_n777), .A3(new_n536), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n777), .B1(new_n762), .B2(new_n536), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n778), .A2(new_n779), .A3(new_n736), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n328), .B(new_n325), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n309), .A4(new_n683), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G140), .ZN(G42));
  NOR2_X1   g597(.A1(new_n680), .A2(new_n681), .ZN(new_n784));
  XOR2_X1   g598(.A(new_n784), .B(KEYINPUT49), .Z(new_n785));
  NOR3_X1   g599(.A1(new_n770), .A2(new_n734), .A3(new_n540), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  INV_X1    g601(.A(new_n658), .ZN(new_n788));
  OR4_X1    g602(.A1(new_n666), .A2(new_n785), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n682), .A2(new_n735), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n425), .B1(new_n790), .B2(KEYINPUT115), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n682), .A2(new_n792), .A3(new_n735), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n666), .A2(new_n683), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n673), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(G952), .A3(new_n269), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n798));
  INV_X1    g612(.A(new_n425), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n724), .A2(new_n771), .A3(new_n799), .A4(new_n734), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n682), .A2(new_n658), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(KEYINPUT50), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n500), .A2(new_n623), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n791), .A2(new_n793), .A3(new_n795), .A4(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n794), .A2(new_n771), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n728), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n803), .A2(new_n808), .A3(new_n810), .A4(KEYINPUT117), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT113), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT113), .B1(new_n680), .B2(new_n681), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n535), .ZN(new_n814));
  OAI22_X1  g628(.A1(new_n778), .A2(new_n779), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n724), .A2(new_n771), .A3(new_n799), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n735), .A3(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n811), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n802), .A2(KEYINPUT50), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n820), .A2(new_n821), .B1(new_n806), .B2(new_n807), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT117), .B1(new_n822), .B2(new_n810), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT118), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n811), .A2(KEYINPUT51), .A3(new_n818), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n826), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n797), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT53), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n685), .A2(new_n691), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n688), .B(new_n831), .C1(new_n719), .C2(new_n725), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n644), .B1(new_n699), .B2(new_n700), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n535), .B(new_n648), .C1(new_n584), .C2(new_n592), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n833), .A2(new_n834), .A3(new_n638), .A4(new_n666), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n677), .A3(new_n729), .A4(new_n650), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n644), .B1(new_n781), .B2(new_n309), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n839), .B(new_n639), .C1(new_n649), .C2(new_n676), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(KEYINPUT52), .A3(new_n729), .A4(new_n835), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT111), .ZN(new_n844));
  INV_X1    g658(.A(new_n431), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n844), .B1(new_n845), .B2(new_n673), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n624), .A2(new_n431), .A3(KEYINPUT111), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n599), .A2(new_n601), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n632), .A2(new_n849), .A3(new_n594), .A4(new_n640), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n738), .A2(new_n741), .B1(new_n746), .B2(new_n748), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n330), .A2(new_n629), .A3(new_n698), .A4(new_n647), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n676), .A2(new_n707), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n639), .A3(new_n735), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n851), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n830), .B1(new_n843), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n742), .A2(new_n749), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n855), .A2(new_n639), .A3(new_n735), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n859), .A2(new_n850), .A3(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n832), .A4(new_n842), .ZN(new_n862));
  XOR2_X1   g676(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n858), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n867), .B1(new_n858), .B2(new_n862), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n817), .A2(new_n645), .A3(new_n682), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n818), .A2(new_n810), .A3(new_n822), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n869), .B(new_n870), .C1(KEYINPUT51), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n683), .B1(new_n781), .B2(new_n309), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n809), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n829), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(G952), .A2(G953), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n789), .B1(new_n877), .B2(new_n878), .ZN(G75));
  AOI21_X1  g693(.A(new_n299), .B1(new_n858), .B2(new_n862), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n421), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n402), .A2(new_n408), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(new_n406), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT55), .Z(new_n885));
  AND3_X1   g699(.A1(new_n881), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n881), .B2(new_n882), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n269), .A2(G952), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G51));
  NAND2_X1  g703(.A1(new_n858), .A2(new_n862), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n863), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(KEYINPUT120), .A3(new_n865), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n754), .A2(KEYINPUT57), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n894), .A3(new_n863), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n754), .A2(KEYINPUT57), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n892), .A2(new_n893), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n582), .ZN(new_n898));
  INV_X1    g712(.A(new_n753), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n880), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n888), .B1(new_n898), .B2(new_n900), .ZN(G54));
  NAND3_X1  g715(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n496), .A2(new_n497), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n902), .A2(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n888), .ZN(G60));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT59), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n866), .B2(new_n868), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n617), .A2(new_n619), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n888), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n911), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n892), .A2(new_n913), .A3(new_n895), .A4(new_n909), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(KEYINPUT121), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n912), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(G63));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT122), .Z(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT60), .Z(new_n922));
  NAND2_X1  g736(.A1(new_n890), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n537), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n888), .ZN(new_n926));
  INV_X1    g740(.A(new_n922), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n858), .B2(new_n862), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n637), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n925), .A2(KEYINPUT61), .A3(new_n926), .A4(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n925), .B2(new_n926), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n932), .B(new_n926), .C1(new_n928), .C2(new_n537), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n929), .ZN(new_n935));
  OAI211_X1 g749(.A(KEYINPUT124), .B(new_n931), .C1(new_n933), .C2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n926), .B1(new_n928), .B2(new_n537), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(new_n934), .A3(new_n929), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT124), .B1(new_n940), .B2(new_n931), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n930), .B1(new_n937), .B2(new_n941), .ZN(G66));
  AOI21_X1  g756(.A(new_n269), .B1(new_n426), .B2(G224), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n832), .A2(new_n851), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n944), .B2(new_n269), .ZN(new_n945));
  MUX2_X1   g759(.A(new_n943), .B(new_n945), .S(KEYINPUT125), .Z(new_n946));
  INV_X1    g760(.A(G898), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n883), .B1(new_n947), .B2(G953), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  INV_X1    g763(.A(G900), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n315), .B(new_n486), .ZN(new_n951));
  OAI21_X1  g765(.A(G953), .B1(new_n951), .B2(new_n567), .ZN(new_n952));
  AOI211_X1 g766(.A(new_n950), .B(new_n952), .C1(new_n567), .C2(new_n951), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n840), .A2(new_n729), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n667), .A2(KEYINPUT62), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT62), .B1(new_n667), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n782), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n654), .B1(new_n624), .B2(new_n630), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n873), .A3(new_n735), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n775), .A2(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n961), .B2(new_n951), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n873), .A2(new_n833), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n765), .B(new_n767), .C1(new_n774), .C2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n964), .A2(new_n782), .A3(new_n852), .A4(new_n954), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n965), .A2(new_n951), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n953), .B1(new_n962), .B2(new_n966), .ZN(G72));
  XNOR2_X1  g781(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n710), .A2(new_n299), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n968), .B(new_n969), .Z(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n965), .B2(new_n944), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n281), .B1(new_n972), .B2(KEYINPUT127), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n974), .B(new_n971), .C1(new_n965), .C2(new_n944), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n971), .B1(new_n961), .B2(new_n944), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n660), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n660), .A2(new_n970), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n890), .A2(new_n281), .A3(new_n979), .ZN(new_n980));
  AND4_X1   g794(.A1(new_n926), .A2(new_n976), .A3(new_n978), .A4(new_n980), .ZN(G57));
endmodule


