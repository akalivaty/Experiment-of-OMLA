//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n577, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT65), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n458), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  NOR3_X1   g040(.A1(new_n463), .A2(G2105), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  INV_X1    g042(.A(G113), .ZN(new_n468));
  OR3_X1    g043(.A1(new_n468), .A2(new_n459), .A3(KEYINPUT67), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n468), .B2(new_n459), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n461), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n476), .A2(new_n477), .A3(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n467), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n466), .A2(G136), .ZN(new_n482));
  NOR3_X1   g057(.A1(KEYINPUT69), .A2(G100), .A3(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(KEYINPUT69), .B1(G100), .B2(G2105), .ZN(new_n484));
  INV_X1    g059(.A(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n482), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(G2104), .ZN(new_n488));
  OAI211_X1 g063(.A(G2105), .B(new_n464), .C1(new_n488), .C2(new_n458), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n487), .B1(G124), .B2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT70), .Z(G162));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(new_n485), .A3(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n473), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT3), .B1(new_n476), .B2(new_n477), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n496), .A2(G138), .A3(new_n485), .A4(new_n464), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n495), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n485), .A2(G114), .ZN(new_n500));
  OAI221_X1 g075(.A(G2104), .B1(G102), .B2(G2105), .C1(new_n500), .C2(KEYINPUT71), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n502));
  OAI22_X1  g077(.A1(new_n489), .A2(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n498), .A2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT72), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(new_n509), .B1(KEYINPUT5), .B2(new_n505), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n510), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(G543), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n513), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n518), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT73), .Z(new_n528));
  INV_X1    g103(.A(new_n521), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n529), .A2(G51), .B1(new_n510), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n506), .A2(new_n509), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n541), .B(new_n534), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n540), .A2(G651), .A3(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n518), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G90), .B1(new_n529), .B2(G52), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n543), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n512), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n518), .A2(new_n549), .B1(new_n550), .B2(new_n521), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT75), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n559), .B(KEYINPUT76), .Z(G188));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n537), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n510), .A2(KEYINPUT78), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(G65), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n512), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n514), .A2(new_n516), .A3(G53), .A4(G543), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT9), .Z(new_n569));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n518), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n510), .A2(KEYINPUT77), .A3(new_n517), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n569), .B1(new_n573), .B2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n567), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n577));
  XNOR2_X1  g152(.A(G166), .B(new_n577), .ZN(G303));
  NAND2_X1  g153(.A1(new_n573), .A2(G87), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n510), .A2(G74), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n529), .B2(G49), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(new_n573), .A2(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n537), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n529), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n544), .A2(G85), .B1(new_n529), .B2(G47), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n512), .B2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n573), .A2(G92), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n562), .A2(G66), .A3(new_n563), .ZN(new_n596));
  INV_X1    g171(.A(G79), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n505), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n592), .B1(new_n600), .B2(G868), .ZN(G321));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g178(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n600), .B1(new_n605), .B2(G860), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT81), .Z(G148));
  INV_X1    g182(.A(new_n600), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n608), .A2(G559), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n552), .ZN(new_n611));
  MUX2_X1   g186(.A(new_n610), .B(new_n611), .S(KEYINPUT82), .Z(G323));
  XNOR2_X1  g187(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g188(.A(G323), .B(new_n613), .ZN(G282));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(G111), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G2105), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n466), .B2(G135), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n490), .A2(KEYINPUT85), .A3(G123), .ZN(new_n619));
  INV_X1    g194(.A(KEYINPUT85), .ZN(new_n620));
  INV_X1    g195(.A(G123), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n489), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n478), .A2(new_n464), .A3(new_n472), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT84), .B(G2100), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n626), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n624), .A2(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2443), .B(G2446), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT87), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2067), .B(G2678), .Z(new_n651));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT17), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT89), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n651), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT88), .B(KEYINPUT18), .Z(new_n659));
  AOI22_X1  g234(.A1(new_n656), .A2(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n655), .B(new_n660), .C1(new_n658), .C2(new_n659), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1971), .B(G1976), .Z(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n670), .A2(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(KEYINPUT20), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n666), .A2(new_n673), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n666), .A2(new_n669), .A3(new_n673), .ZN(new_n675));
  NAND4_X1  g250(.A1(new_n671), .A2(new_n672), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT91), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n676), .B(new_n682), .ZN(G229));
  MUX2_X1   g258(.A(G24), .B(G290), .S(G16), .Z(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G1986), .Z(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G25), .ZN(new_n687));
  OR2_X1    g262(.A1(G95), .A2(G2105), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n688), .B(G2104), .C1(G107), .C2(new_n485), .ZN(new_n689));
  INV_X1    g264(.A(new_n466), .ZN(new_n690));
  INV_X1    g265(.A(G131), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g267(.A1(new_n490), .A2(G119), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n687), .B1(new_n694), .B2(new_n686), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT35), .B(G1991), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NOR2_X1   g274(.A1(G166), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(G22), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n700), .A2(G1971), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n699), .A2(G6), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G305), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT32), .B(G1981), .Z(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g281(.A(G1971), .B1(new_n700), .B2(new_n701), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G288), .B(KEYINPUT92), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n699), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n712), .B(new_n715), .C1(new_n713), .C2(new_n699), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n710), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n685), .B(new_n698), .C1(new_n719), .C2(KEYINPUT34), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT93), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(KEYINPUT34), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT36), .ZN(new_n724));
  NOR2_X1   g299(.A1(G29), .A2(G35), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G162), .B2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT29), .ZN(new_n727));
  INV_X1    g302(.A(G2090), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n473), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(new_n485), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT98), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n485), .A2(G103), .A3(G2104), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT97), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT25), .Z(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G139), .B2(new_n466), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n738), .A2(new_n686), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n686), .B2(G33), .ZN(new_n740));
  INV_X1    g315(.A(G2072), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n686), .B1(KEYINPUT24), .B2(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(KEYINPUT24), .B2(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n480), .B2(G29), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n623), .A2(new_n686), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n752), .A2(G28), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n686), .B1(new_n752), .B2(G28), .ZN(new_n754));
  AND2_X1   g329(.A1(KEYINPUT31), .A2(G11), .ZN(new_n755));
  NOR2_X1   g330(.A1(KEYINPUT31), .A2(G11), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n753), .A2(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n745), .B2(new_n746), .ZN(new_n758));
  NAND4_X1  g333(.A1(new_n742), .A2(new_n750), .A3(new_n751), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n552), .A2(new_n699), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n699), .B2(G19), .ZN(new_n761));
  INV_X1    g336(.A(G1341), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n761), .A2(new_n762), .B1(new_n748), .B2(new_n749), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n740), .B2(new_n741), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n699), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n699), .ZN(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n699), .A2(G5), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G171), .B2(new_n699), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI22_X1  g346(.A1(new_n767), .A2(G1966), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NOR4_X1   g347(.A1(new_n759), .A2(new_n763), .A3(new_n765), .A4(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n699), .A2(G4), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n600), .B2(new_n699), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT94), .B(G1348), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT95), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n775), .B(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT23), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n699), .A2(G20), .ZN(new_n781));
  MUX2_X1   g356(.A(new_n779), .B(new_n780), .S(new_n781), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n767), .A2(G1966), .B1(new_n768), .B2(new_n771), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n686), .A2(G26), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT96), .ZN(new_n786));
  OR3_X1    g361(.A1(new_n786), .A2(G104), .A3(G2105), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(G104), .B2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(G116), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n459), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G128), .ZN(new_n792));
  INV_X1    g367(.A(G140), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n791), .B1(new_n792), .B2(new_n489), .C1(new_n690), .C2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n785), .B1(new_n795), .B2(new_n686), .ZN(new_n796));
  MUX2_X1   g371(.A(new_n785), .B(new_n796), .S(KEYINPUT28), .Z(new_n797));
  INV_X1    g372(.A(G2067), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AND4_X1   g374(.A1(new_n778), .A2(new_n783), .A3(new_n784), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n490), .A2(G129), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n466), .A2(G141), .ZN(new_n802));
  NAND3_X1  g377(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT26), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G105), .B2(new_n478), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n801), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G32), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT27), .B(G1996), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(G27), .A2(G29), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G164), .B2(G29), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G2078), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n729), .A2(new_n773), .A3(new_n800), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT100), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n724), .A2(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  AOI22_X1  g392(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n512), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n518), .A2(new_n820), .B1(new_n821), .B2(new_n521), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n600), .A2(G559), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n823), .B(new_n552), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT101), .ZN(new_n832));
  INV_X1    g407(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(G860), .B1(new_n829), .B2(new_n830), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n831), .B2(KEYINPUT101), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n825), .B1(new_n833), .B2(new_n835), .ZN(G145));
  INV_X1    g411(.A(KEYINPUT102), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n738), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G164), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n794), .B(new_n806), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n694), .B(new_n626), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n466), .A2(G142), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n485), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n490), .A2(G130), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n847), .B2(new_n848), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n842), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n841), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(KEYINPUT104), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n841), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G162), .B(new_n480), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n623), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(G37), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n856), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g437(.A(new_n713), .B(G290), .Z(new_n863));
  XNOR2_X1  g438(.A(G305), .B(G166), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n609), .B(new_n828), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n600), .B(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(KEYINPUT41), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n870), .B1(new_n871), .B2(new_n868), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n867), .A2(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(KEYINPUT105), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n874), .A2(KEYINPUT105), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n823), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(G868), .B2(new_n878), .ZN(G295));
  OAI21_X1  g454(.A(new_n877), .B1(G868), .B2(new_n878), .ZN(G331));
  NAND2_X1  g455(.A1(new_n871), .A2(KEYINPUT109), .ZN(new_n881));
  NOR2_X1   g456(.A1(G171), .A2(KEYINPUT108), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n828), .B(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(G286), .B1(KEYINPUT108), .B2(G171), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n869), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n869), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n865), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n891), .B(new_n865), .C1(new_n871), .C2(new_n885), .ZN(new_n893));
  INV_X1    g468(.A(G37), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n891), .B1(new_n871), .B2(new_n885), .ZN(new_n898));
  INV_X1    g473(.A(new_n865), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n897), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(new_n903), .A3(KEYINPUT44), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n892), .A2(new_n895), .A3(new_n901), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n902), .B1(new_n897), .B2(new_n900), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n904), .B1(new_n907), .B2(new_n908), .ZN(G397));
  INV_X1    g484(.A(G1384), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n910), .B1(new_n498), .B2(new_n503), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n467), .A2(new_n475), .A3(G40), .A4(new_n479), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n794), .B(new_n798), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(KEYINPUT110), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n919), .A2(KEYINPUT110), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n806), .B(G1996), .ZN(new_n922));
  AOI211_X1 g497(.A(new_n920), .B(new_n921), .C1(new_n915), .C2(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n694), .A2(new_n697), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n692), .A2(new_n693), .A3(new_n696), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(G1986), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n915), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT113), .ZN(new_n930));
  NAND4_X1  g505(.A1(G303), .A2(new_n930), .A3(KEYINPUT55), .A4(G8), .ZN(new_n931));
  NOR2_X1   g506(.A1(G166), .A2(new_n577), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n513), .A2(new_n522), .A3(KEYINPUT79), .ZN(new_n933));
  OAI211_X1 g508(.A(KEYINPUT55), .B(G8), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT113), .ZN(new_n935));
  OAI21_X1  g510(.A(G8), .B1(new_n932), .B2(new_n933), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n931), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1971), .ZN(new_n941));
  INV_X1    g516(.A(new_n914), .ZN(new_n942));
  OAI211_X1 g517(.A(KEYINPUT45), .B(new_n910), .C1(new_n498), .C2(new_n503), .ZN(new_n943));
  AND4_X1   g518(.A1(KEYINPUT111), .A2(new_n913), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n914), .B1(new_n911), .B2(new_n912), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT111), .B1(new_n945), .B2(new_n943), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n941), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n911), .A2(new_n948), .ZN(new_n949));
  OAI211_X1 g524(.A(KEYINPUT112), .B(new_n910), .C1(new_n498), .C2(new_n503), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT50), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(new_n910), .C1(new_n498), .C2(new_n503), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n953), .A2(new_n942), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n728), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n947), .A2(KEYINPUT116), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(G8), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT116), .B1(new_n947), .B2(new_n955), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n940), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT117), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT117), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n961), .B(new_n940), .C1(new_n957), .C2(new_n958), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n913), .A2(new_n942), .A3(new_n943), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n945), .A2(KEYINPUT111), .A3(new_n943), .ZN(new_n966));
  AOI21_X1  g541(.A(G1971), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT50), .B1(new_n949), .B2(new_n950), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n914), .B1(new_n911), .B2(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n968), .A2(new_n970), .A3(G2090), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n939), .B(G8), .C1(new_n967), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n914), .B1(new_n949), .B2(new_n950), .ZN(new_n973));
  INV_X1    g548(.A(G8), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1976), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(G288), .B2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n975), .B(new_n977), .C1(new_n976), .C2(new_n713), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n975), .B1(new_n713), .B2(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT52), .ZN(new_n980));
  INV_X1    g555(.A(G1981), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n583), .A2(new_n981), .A3(new_n587), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n544), .A2(G86), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n587), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n982), .B1(new_n984), .B2(new_n981), .ZN(new_n985));
  NOR2_X1   g560(.A1(KEYINPUT114), .A2(KEYINPUT49), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n975), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n972), .A2(new_n978), .A3(new_n980), .A4(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n960), .A2(new_n962), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2078), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n965), .A2(new_n993), .A3(new_n966), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n949), .A2(new_n950), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n952), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n969), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n768), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n913), .A2(new_n942), .A3(new_n943), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n995), .A2(G2078), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n996), .A2(G301), .A3(new_n1000), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n949), .A2(new_n912), .A3(new_n950), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n942), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(KEYINPUT118), .A3(new_n942), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n943), .A4(new_n1002), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1010), .A2(new_n996), .A3(new_n1000), .ZN(new_n1011));
  AOI22_X1  g586(.A1(KEYINPUT125), .A2(new_n1004), .B1(new_n1011), .B2(G171), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n994), .A2(new_n995), .B1(new_n999), .B2(new_n768), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT125), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n1014), .A3(G301), .A4(new_n1003), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT54), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n992), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT124), .B1(G286), .B2(G8), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(KEYINPUT51), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT119), .B(G2084), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n998), .A2(new_n969), .A3(new_n1020), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1005), .A2(KEYINPUT118), .A3(new_n942), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT118), .B1(new_n1005), .B2(new_n942), .ZN(new_n1023));
  INV_X1    g598(.A(new_n943), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(G1966), .ZN(new_n1026));
  OAI211_X1 g601(.A(G8), .B(new_n1019), .C1(new_n1026), .C2(G286), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G286), .A2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1019), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1021), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1008), .A2(new_n1009), .A3(new_n943), .ZN(new_n1031));
  INV_X1    g606(.A(G1966), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1028), .B(new_n1029), .C1(new_n1033), .C2(new_n974), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1026), .A2(G8), .A3(G286), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1027), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1013), .A2(new_n1003), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1037), .B1(new_n1038), .B2(G171), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G171), .B2(new_n1011), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT126), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1017), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1011), .A2(G171), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1004), .A2(KEYINPUT125), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1045), .A3(new_n1015), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n1037), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n990), .B1(KEYINPUT117), .B2(new_n959), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n962), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT126), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n951), .A2(new_n954), .ZN(new_n1053));
  INV_X1    g628(.A(G1956), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1053), .A2(new_n1054), .B1(new_n1001), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n567), .A2(new_n574), .A3(KEYINPUT57), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n1058));
  INV_X1    g633(.A(new_n572), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT77), .B1(new_n510), .B2(new_n517), .ZN(new_n1060));
  OAI21_X1  g635(.A(G91), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n569), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1058), .B1(new_n1063), .B2(new_n566), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1057), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1052), .B1(new_n1056), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1956), .B1(new_n951), .B2(new_n954), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n945), .A2(new_n943), .A3(new_n1055), .ZN(new_n1069));
  NOR4_X1   g644(.A1(new_n1068), .A2(new_n1065), .A3(new_n1069), .A4(KEYINPUT120), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1065), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT61), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1056), .A2(new_n1066), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1072), .ZN(new_n1075));
  INV_X1    g650(.A(new_n973), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT58), .B(G1341), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(KEYINPUT121), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1996), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1001), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n973), .B2(new_n1077), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n552), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n1084), .B2(new_n552), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1075), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT122), .B1(new_n1073), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1074), .A2(KEYINPUT120), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1056), .A2(new_n1052), .A3(new_n1066), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(new_n1072), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT61), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1084), .A2(new_n552), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT59), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1084), .A2(new_n1085), .A3(new_n552), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1094), .A2(new_n1095), .A3(new_n1075), .A4(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n1101));
  INV_X1    g676(.A(G1348), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n968), .B2(new_n970), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n973), .A2(new_n798), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1101), .B(new_n600), .C1(new_n1105), .C2(KEYINPUT60), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1105), .A2(KEYINPUT60), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT60), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT123), .B1(new_n1108), .B2(new_n608), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1106), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1089), .A2(new_n1100), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1072), .B1(new_n1105), .B2(new_n608), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1071), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1043), .A2(new_n1051), .A3(new_n1116), .ZN(new_n1117));
  AND4_X1   g692(.A1(new_n976), .A2(new_n989), .A3(new_n579), .A4(new_n581), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n982), .B(KEYINPUT115), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n975), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n980), .A2(new_n978), .A3(new_n989), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(new_n972), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1033), .A2(new_n974), .A3(G286), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1121), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n967), .A2(new_n971), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n940), .B1(new_n1125), .B2(new_n974), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1123), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1122), .B1(new_n1127), .B2(KEYINPUT63), .ZN(new_n1128));
  NOR4_X1   g703(.A1(new_n1033), .A2(KEYINPUT63), .A3(new_n974), .A4(G286), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1044), .B1(new_n1036), .B2(KEYINPUT62), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1027), .A2(new_n1034), .A3(new_n1035), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1128), .B1(new_n1133), .B2(new_n992), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n929), .B1(new_n1117), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n923), .A2(new_n925), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n795), .A2(new_n798), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n916), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n917), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n915), .B1(new_n1139), .B2(new_n806), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT46), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n916), .B2(G1996), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n915), .A2(KEYINPUT46), .A3(new_n1080), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(new_n1144), .B(KEYINPUT127), .Z(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT47), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n916), .A2(G1986), .A3(G290), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1147), .B(KEYINPUT48), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n927), .A2(new_n1148), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1138), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1135), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g726(.A(G319), .ZN(new_n1153));
  NOR3_X1   g727(.A1(G227), .A2(new_n1153), .A3(G229), .ZN(new_n1154));
  NAND3_X1  g728(.A1(new_n861), .A2(new_n646), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g729(.A1(new_n907), .A2(new_n1155), .ZN(G308));
  OR2_X1    g730(.A1(new_n907), .A2(new_n1155), .ZN(G225));
endmodule


