//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT86), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT86), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  AOI21_X1  g005(.A(G50gat), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT87), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT87), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G50gat), .ZN(new_n211));
  AOI21_X1  g010(.A(G43gat), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(new_n207), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n202), .B1(G43gat), .B2(new_n208), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(G50gat), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT85), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT15), .B1(new_n203), .B2(G50gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n208), .A2(G43gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT85), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(G36gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT14), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT14), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G29gat), .B2(G36gat), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT88), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT88), .B1(new_n225), .B2(new_n227), .ZN(new_n229));
  OAI22_X1  g028(.A1(new_n218), .A2(new_n222), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT84), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n225), .A2(new_n227), .A3(new_n214), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n219), .A2(new_n220), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n232), .A2(new_n233), .A3(new_n231), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n215), .A2(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G22gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G15gat), .ZN(new_n240));
  INV_X1    g039(.A(G15gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G22gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT89), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n240), .B2(new_n242), .ZN(new_n245));
  INV_X1    g044(.A(G1gat), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n246), .A2(KEYINPUT16), .ZN(new_n247));
  NOR3_X1   g046(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n241), .A2(G22gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n239), .A2(G15gat), .ZN(new_n250));
  OAI21_X1  g049(.A(KEYINPUT89), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n252));
  AOI21_X1  g051(.A(G1gat), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(G8gat), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n246), .B1(new_n244), .B2(new_n245), .ZN(new_n255));
  INV_X1    g054(.A(G8gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(new_n252), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n255), .B(new_n256), .C1(new_n247), .C2(new_n257), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  OAI221_X1 g058(.A(KEYINPUT17), .B1(new_n234), .B2(new_n235), .C1(new_n215), .C2(new_n230), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n238), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G229gat), .A2(G233gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n254), .A2(new_n258), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT90), .ZN(new_n264));
  AND3_X1   g063(.A1(new_n263), .A2(new_n236), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n264), .B1(new_n263), .B2(new_n236), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n261), .B(new_n262), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT18), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n267), .A2(KEYINPUT92), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT92), .B1(new_n267), .B2(new_n268), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n266), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n263), .A2(new_n236), .A3(new_n264), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n274), .A2(KEYINPUT18), .A3(new_n262), .A4(new_n261), .ZN(new_n275));
  OAI22_X1  g074(.A1(new_n265), .A2(new_n266), .B1(new_n236), .B2(new_n263), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n262), .B(KEYINPUT13), .Z(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G141gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G169gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(G197gat), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n281), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G197gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n283), .A2(new_n287), .A3(KEYINPUT12), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT12), .B1(new_n283), .B2(new_n287), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n278), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT93), .B1(new_n271), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n267), .A2(new_n268), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n267), .A2(KEYINPUT92), .A3(new_n268), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n275), .A2(new_n278), .A3(new_n290), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT93), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n293), .A2(new_n275), .A3(new_n278), .ZN(new_n302));
  INV_X1    g101(.A(new_n290), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT91), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(KEYINPUT91), .A3(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT94), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n292), .A2(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT94), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT36), .ZN(new_n315));
  XNOR2_X1  g114(.A(G15gat), .B(G43gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G71gat), .B(G99gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n322), .B(new_n323), .C1(new_n320), .C2(new_n321), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n320), .A2(new_n321), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(G113gat), .B2(G120gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT67), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n319), .B1(new_n324), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n328), .A2(new_n319), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n332));
  INV_X1    g131(.A(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G183gat), .A2(G190gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(KEYINPUT24), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n284), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OR2_X1    g140(.A1(new_n336), .A2(KEYINPUT24), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n337), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G169gat), .A2(G176gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n339), .B2(new_n340), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n332), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT64), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT64), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n348), .B(new_n332), .C1(new_n343), .C2(new_n345), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n343), .A2(new_n332), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(KEYINPUT65), .B(new_n344), .C1(new_n339), .C2(new_n340), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n347), .A2(new_n349), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356));
  NOR2_X1   g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n357), .A2(KEYINPUT66), .A3(new_n356), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT66), .B1(new_n357), .B2(new_n356), .ZN(new_n359));
  OAI221_X1 g158(.A(new_n344), .B1(new_n356), .B2(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT27), .B(G183gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n334), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n362), .A2(KEYINPUT28), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n362), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n360), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n331), .B1(new_n355), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n354), .A2(new_n350), .ZN(new_n368));
  INV_X1    g167(.A(new_n345), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n369), .A2(new_n337), .A3(new_n341), .A4(new_n342), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n348), .B1(new_n370), .B2(new_n332), .ZN(new_n371));
  INV_X1    g170(.A(new_n349), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n368), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n331), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(new_n365), .ZN(new_n375));
  INV_X1    g174(.A(G227gat), .ZN(new_n376));
  INV_X1    g175(.A(G233gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n367), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT33), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n318), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(KEYINPUT32), .ZN(new_n382));
  OR2_X1    g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n382), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n375), .ZN(new_n386));
  INV_X1    g185(.A(new_n378), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n388), .A2(KEYINPUT34), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(KEYINPUT34), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n385), .A2(new_n391), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n315), .B1(new_n394), .B2(KEYINPUT68), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT68), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(KEYINPUT36), .C1(new_n392), .C2(new_n393), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n400), .B1(new_n355), .B2(new_n366), .ZN(new_n401));
  INV_X1    g200(.A(G226gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(new_n377), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT73), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G197gat), .B(G204gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT22), .ZN(new_n408));
  INV_X1    g207(.A(G211gat), .ZN(new_n409));
  INV_X1    g208(.A(G218gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G211gat), .B(G218gat), .Z(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT70), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n413), .A2(KEYINPUT69), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(KEYINPUT69), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n415), .A2(KEYINPUT71), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT71), .B1(new_n415), .B2(new_n418), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n404), .B1(new_n373), .B2(new_n365), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n401), .B2(new_n404), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT73), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n406), .B(new_n422), .C1(new_n424), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT72), .ZN(new_n427));
  NOR3_X1   g226(.A1(new_n424), .A2(new_n427), .A3(new_n422), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n401), .A2(new_n404), .ZN(new_n429));
  INV_X1    g228(.A(new_n423), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n422), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT72), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n426), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT74), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n427), .B1(new_n424), .B2(new_n422), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n431), .A2(KEYINPUT72), .A3(new_n432), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n439), .A2(KEYINPUT74), .A3(new_n426), .ZN(new_n440));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G64gat), .ZN(new_n442));
  INV_X1    g241(.A(G92gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n436), .A2(new_n440), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT5), .ZN(new_n447));
  XOR2_X1   g246(.A(G155gat), .B(G162gat), .Z(new_n448));
  XNOR2_X1  g247(.A(G141gat), .B(G148gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(KEYINPUT2), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n448), .A2(new_n449), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT75), .B(G162gat), .ZN(new_n453));
  INV_X1    g252(.A(G155gat), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT2), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n452), .B1(new_n451), .B2(new_n455), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n450), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n374), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n331), .B(new_n450), .C1(new_n457), .C2(new_n458), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n447), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n466), .A3(KEYINPUT4), .ZN(new_n467));
  INV_X1    g266(.A(new_n450), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n455), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT76), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n470), .B2(new_n456), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT3), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n374), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n467), .B(new_n463), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n461), .A2(KEYINPUT4), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n471), .A2(new_n477), .A3(new_n331), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n476), .A2(KEYINPUT77), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n465), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n473), .A2(new_n474), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n476), .A2(new_n478), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(new_n482), .A3(new_n447), .A4(new_n463), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G1gat), .B(G29gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n485), .B(KEYINPUT0), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(G57gat), .ZN(new_n487));
  INV_X1    g286(.A(G85gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n480), .A2(new_n483), .A3(new_n489), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n484), .A2(KEYINPUT6), .A3(new_n490), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n439), .A2(new_n426), .A3(new_n444), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n405), .B1(new_n431), .B2(KEYINPUT73), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n422), .A2(new_n500), .B1(new_n437), .B2(new_n438), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n444), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n446), .A2(new_n496), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT78), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n502), .A2(new_n499), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT78), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n496), .A4(new_n446), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n432), .B1(KEYINPUT29), .B2(new_n474), .ZN(new_n509));
  NAND2_X1  g308(.A1(G228gat), .A2(G233gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n415), .A2(new_n418), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT3), .B1(new_n512), .B2(new_n400), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n509), .B(new_n511), .C1(new_n471), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n412), .A2(new_n413), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT29), .B1(new_n415), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n459), .B1(new_n516), .B2(KEYINPUT3), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n517), .A2(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(KEYINPUT80), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n509), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n510), .B(KEYINPUT79), .Z(new_n521));
  OAI21_X1  g320(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT31), .B(G50gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(new_n239), .ZN(new_n526));
  NAND2_X1  g325(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(new_n525), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n522), .B(new_n528), .Z(new_n529));
  OAI211_X1 g328(.A(KEYINPUT82), .B(new_n399), .C1(new_n508), .C2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT40), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n463), .B1(new_n481), .B2(new_n482), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT39), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n489), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT39), .B1(new_n462), .B2(new_n464), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n531), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n490), .B1(new_n532), .B2(new_n533), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n539), .B(KEYINPUT40), .C1(new_n532), .C2(new_n536), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n538), .A2(new_n491), .A3(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n436), .A2(new_n440), .A3(new_n445), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n502), .A2(new_n499), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n444), .B1(new_n501), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n500), .A2(new_n432), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT37), .B1(new_n424), .B2(new_n432), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n425), .B1(new_n429), .B2(new_n430), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n552), .A2(new_n422), .A3(new_n405), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT83), .B1(new_n553), .B2(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT38), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n496), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n497), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n436), .A2(KEYINPUT37), .A3(new_n440), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n556), .B1(new_n560), .B2(new_n546), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n544), .B(new_n529), .C1(new_n559), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT82), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n529), .B1(new_n504), .B2(new_n507), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n398), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n530), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n394), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n522), .B(new_n528), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n569), .A2(new_n504), .A3(new_n507), .ZN(new_n570));
  INV_X1    g369(.A(new_n503), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT35), .ZN(new_n572));
  AOI22_X1  g371(.A1(new_n570), .A2(KEYINPUT35), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n314), .B1(new_n566), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G71gat), .B(G78gat), .Z(new_n577));
  INV_X1    g376(.A(G57gat), .ZN(new_n578));
  INV_X1    g377(.A(G64gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G78gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT9), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592));
  OAI21_X1  g391(.A(G64gat), .B1(new_n592), .B2(new_n578), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n579), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n585), .A2(KEYINPUT96), .A3(new_n586), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n589), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT97), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n577), .A2(KEYINPUT96), .B1(new_n593), .B2(new_n594), .ZN(new_n600));
  AOI22_X1  g399(.A1(new_n587), .A2(new_n588), .B1(new_n590), .B2(new_n586), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n599), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n582), .B1(new_n598), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n263), .B1(new_n604), .B2(KEYINPUT21), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G183gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n604), .A2(KEYINPUT21), .ZN(new_n611));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(new_n409), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT7), .ZN(new_n619));
  OR2_X1    g418(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n488), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G99gat), .A2(G106gat), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT8), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G99gat), .B(G106gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n236), .A2(new_n628), .B1(KEYINPUT41), .B2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n625), .B(new_n626), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n238), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n260), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT98), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n636), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n630), .B(new_n638), .C1(new_n632), .C2(new_n633), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G190gat), .B(G218gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n640), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G176gat), .ZN(new_n648));
  INV_X1    g447(.A(G204gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n603), .A2(new_n631), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n597), .A2(KEYINPUT97), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n600), .A2(new_n599), .A3(new_n601), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n628), .A2(new_n654), .A3(new_n582), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G230gat), .A2(G233gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(new_n660), .A3(new_n655), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n657), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n650), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n657), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n661), .B2(new_n662), .ZN(new_n667));
  INV_X1    g466(.A(new_n650), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n658), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n617), .A2(new_n646), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n576), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n496), .B(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT101), .B(G1gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n505), .A2(new_n446), .ZN(new_n679));
  INV_X1    g478(.A(new_n671), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT16), .B(G8gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n575), .A2(new_n679), .A3(new_n680), .A4(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684));
  AND3_X1   g483(.A1(new_n683), .A2(KEYINPUT102), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT102), .B1(new_n683), .B2(new_n684), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n575), .A2(new_n679), .A3(new_n680), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(G8gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n684), .B2(new_n683), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT103), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n683), .ZN(new_n692));
  AOI22_X1  g491(.A1(new_n692), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n688), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n693), .B(new_n694), .C1(new_n686), .C2(new_n685), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(G1325gat));
  AOI21_X1  g495(.A(G15gat), .B1(new_n672), .B2(new_n394), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT104), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(KEYINPUT104), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n399), .A2(new_n241), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n698), .A2(new_n699), .B1(new_n672), .B2(new_n700), .ZN(G1326gat));
  NAND2_X1  g500(.A1(new_n672), .A2(new_n568), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  NAND2_X1  g503(.A1(new_n566), .A2(new_n574), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n646), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n562), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n564), .A3(new_n398), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n573), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n706), .B1(new_n711), .B2(new_n646), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n670), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n617), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n309), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G29gat), .B1(new_n719), .B2(new_n674), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n645), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n223), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n674), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n575), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n721), .B1(new_n575), .B2(new_n725), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n720), .A2(KEYINPUT105), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n713), .A2(new_n717), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n223), .B1(new_n732), .B2(new_n675), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(new_n728), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(G1328gat));
  INV_X1    g534(.A(new_n679), .ZN(new_n736));
  OAI21_X1  g535(.A(G36gat), .B1(new_n719), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n575), .A2(new_n224), .A3(new_n679), .A4(new_n723), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT46), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1329gat));
  NAND4_X1  g539(.A1(new_n708), .A2(new_n712), .A3(new_n398), .A4(new_n718), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n204), .A2(new_n206), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT47), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n575), .A2(new_n742), .A3(new_n394), .A4(new_n723), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n746), .B(new_n748), .ZN(G1330gat));
  NAND4_X1  g548(.A1(new_n708), .A2(new_n712), .A3(new_n568), .A4(new_n718), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n209), .A2(new_n211), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n722), .A2(new_n752), .A3(new_n529), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n575), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1331gat));
  OAI211_X1 g558(.A(new_n399), .B(new_n562), .C1(new_n508), .C2(new_n529), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n574), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n617), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n762), .A2(new_n309), .A3(new_n645), .A4(new_n670), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n674), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(new_n578), .ZN(G1332gat));
  INV_X1    g565(.A(new_n764), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n679), .B1(new_n768), .B2(new_n579), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT108), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n579), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n764), .B2(new_n399), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n394), .A2(new_n583), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n764), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g576(.A1(new_n764), .A2(new_n529), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(new_n584), .ZN(G1335gat));
  NOR3_X1   g578(.A1(new_n617), .A2(new_n309), .A3(new_n670), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n714), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(G85gat), .B1(new_n781), .B2(new_n674), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n617), .A2(new_n309), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n645), .A4(new_n783), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n645), .B(new_n783), .C1(new_n710), .C2(new_n573), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n715), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n675), .A2(new_n488), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n782), .B1(new_n789), .B2(new_n790), .ZN(G1336gat));
  NAND4_X1  g590(.A1(new_n708), .A2(new_n712), .A3(new_n679), .A4(new_n780), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n620), .A2(new_n621), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  INV_X1    g594(.A(new_n788), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n679), .A2(new_n443), .A3(new_n715), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n794), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(KEYINPUT109), .ZN(new_n800));
  OR2_X1    g599(.A1(new_n797), .A2(KEYINPUT109), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n788), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n794), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n803), .B2(KEYINPUT52), .ZN(new_n804));
  AOI211_X1 g603(.A(KEYINPUT110), .B(new_n795), .C1(new_n794), .C2(new_n802), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n798), .B1(new_n804), .B2(new_n805), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n781), .B2(new_n399), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n567), .A2(G99gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n789), .B2(new_n808), .ZN(G1338gat));
  NOR3_X1   g608(.A1(new_n529), .A2(G106gat), .A3(new_n670), .ZN(new_n810));
  XOR2_X1   g609(.A(new_n810), .B(KEYINPUT111), .Z(new_n811));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(KEYINPUT53), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n708), .A2(new_n712), .A3(new_n568), .A4(new_n780), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT112), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n815), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(G106gat), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n813), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n814), .A2(G106gat), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT53), .B1(new_n820), .B2(new_n812), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1339gat));
  NOR2_X1   g621(.A1(new_n671), .A2(new_n309), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n262), .B1(new_n274), .B2(new_n261), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n276), .A2(new_n277), .ZN(new_n826));
  INV_X1    g625(.A(new_n283), .ZN(new_n827));
  INV_X1    g626(.A(new_n287), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n825), .A2(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n271), .A2(KEYINPUT93), .A3(new_n291), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n299), .B1(new_n297), .B2(new_n298), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n715), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n650), .B1(new_n667), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n669), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT113), .A4(KEYINPUT55), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n834), .A2(KEYINPUT55), .A3(new_n836), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n839), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n832), .B1(new_n312), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n839), .A2(new_n843), .A3(new_n645), .A4(new_n840), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n847), .B2(KEYINPUT114), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n301), .A2(new_n849), .A3(new_n829), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n646), .A2(new_n845), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n762), .B1(new_n851), .B2(KEYINPUT115), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n646), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n850), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT115), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n824), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT116), .B1(new_n857), .B2(new_n568), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n859), .A3(new_n529), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n674), .A2(new_n679), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n394), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n314), .A2(new_n320), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n857), .A2(new_n568), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n864), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n320), .B1(new_n868), .B2(new_n312), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT117), .ZN(G1340gat));
  NAND4_X1  g670(.A1(new_n861), .A2(G120gat), .A3(new_n715), .A4(new_n864), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n321), .B1(new_n868), .B2(new_n670), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT118), .ZN(G1341gat));
  NAND4_X1  g674(.A1(new_n861), .A2(G127gat), .A3(new_n617), .A4(new_n864), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n868), .A2(new_n762), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(G127gat), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(G1342gat));
  NOR3_X1   g681(.A1(new_n868), .A2(G134gat), .A3(new_n646), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT56), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n646), .B(new_n863), .C1(new_n858), .C2(new_n860), .ZN(new_n885));
  INV_X1    g684(.A(G134gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(G1343gat));
  NOR2_X1   g686(.A1(new_n857), .A2(new_n529), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n399), .A2(new_n862), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(G141gat), .A3(new_n314), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(KEYINPUT58), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n309), .A2(new_n310), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n312), .A2(KEYINPUT94), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n844), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n832), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n646), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n617), .B1(new_n898), .B2(new_n854), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n568), .B1(new_n899), .B2(new_n823), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT57), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n856), .A2(new_n902), .A3(new_n568), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n890), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(G141gat), .B1(new_n904), .B2(new_n314), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n893), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n901), .A2(new_n309), .A3(new_n890), .A4(new_n903), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n907), .A2(KEYINPUT120), .A3(G141gat), .ZN(new_n908));
  AOI21_X1  g707(.A(KEYINPUT120), .B1(new_n907), .B2(G141gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n892), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT58), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(G1344gat));
  INV_X1    g711(.A(new_n891), .ZN(new_n913));
  INV_X1    g712(.A(G148gat), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(new_n914), .A3(new_n715), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n904), .A2(new_n670), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n916), .A2(KEYINPUT59), .A3(new_n914), .ZN(new_n917));
  XNOR2_X1  g716(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n902), .B1(new_n856), .B2(new_n568), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n568), .A2(new_n902), .ZN(new_n920));
  INV_X1    g719(.A(new_n844), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n921), .B1(new_n311), .B2(new_n313), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n645), .B1(new_n922), .B2(new_n832), .ZN(new_n923));
  INV_X1    g722(.A(new_n854), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n762), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n314), .A2(new_n680), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT122), .B1(new_n919), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n902), .A2(KEYINPUT122), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n856), .A2(new_n568), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n928), .A2(new_n715), .A3(new_n890), .A4(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n918), .B1(new_n931), .B2(G148gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n915), .B1(new_n917), .B2(new_n932), .ZN(G1345gat));
  OAI21_X1  g732(.A(G155gat), .B1(new_n904), .B2(new_n762), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n617), .A2(new_n454), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n891), .B2(new_n935), .ZN(G1346gat));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n453), .A3(new_n645), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n904), .A2(new_n646), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n453), .ZN(G1347gat));
  OAI21_X1  g738(.A(KEYINPUT123), .B1(new_n857), .B2(new_n675), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n856), .A2(new_n941), .A3(new_n674), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n569), .A2(new_n679), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n309), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n674), .A2(new_n679), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n394), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n949), .B1(new_n858), .B2(new_n860), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n314), .A2(new_n284), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n946), .A2(new_n284), .B1(new_n950), .B2(new_n951), .ZN(G1348gat));
  AND2_X1   g751(.A1(new_n950), .A2(new_n715), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n943), .A2(new_n945), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n715), .A2(new_n338), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n953), .A2(new_n338), .B1(new_n954), .B2(new_n955), .ZN(G1349gat));
  NAND2_X1  g755(.A1(new_n617), .A2(new_n361), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n333), .B1(new_n950), .B2(new_n617), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(KEYINPUT60), .B1(new_n958), .B2(new_n959), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1350gat));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n645), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(G190gat), .ZN(new_n967));
  AOI211_X1 g766(.A(KEYINPUT61), .B(new_n334), .C1(new_n950), .C2(new_n645), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n645), .A2(new_n334), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n954), .B2(new_n969), .ZN(G1351gat));
  NAND2_X1  g769(.A1(new_n948), .A2(new_n399), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n971), .B(new_n972), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n928), .A2(new_n930), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n314), .A2(new_n286), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n398), .A2(new_n736), .A3(new_n529), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n943), .A2(new_n309), .A3(new_n976), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n974), .A2(new_n975), .B1(new_n977), .B2(new_n286), .ZN(G1352gat));
  NAND4_X1  g777(.A1(new_n943), .A2(new_n649), .A3(new_n715), .A4(new_n976), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n981));
  AND4_X1   g780(.A1(new_n715), .A2(new_n928), .A3(new_n930), .A4(new_n973), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n980), .B(new_n981), .C1(new_n649), .C2(new_n982), .ZN(G1353gat));
  NAND4_X1  g782(.A1(new_n928), .A2(new_n617), .A3(new_n930), .A4(new_n973), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G211gat), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT63), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n984), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(KEYINPUT126), .A3(new_n988), .ZN(new_n989));
  AND4_X1   g788(.A1(new_n409), .A2(new_n943), .A3(new_n617), .A4(new_n976), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n984), .B2(G211gat), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n989), .A2(new_n993), .ZN(G1354gat));
  NOR2_X1   g793(.A1(new_n646), .A2(new_n410), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n943), .A2(new_n645), .A3(new_n976), .ZN(new_n996));
  AOI22_X1  g795(.A1(new_n974), .A2(new_n995), .B1(new_n996), .B2(new_n410), .ZN(G1355gat));
endmodule


