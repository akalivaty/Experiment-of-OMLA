

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756;

  XNOR2_X1 U372 ( .A(n400), .B(KEYINPUT104), .ZN(n753) );
  XNOR2_X1 U373 ( .A(n379), .B(KEYINPUT35), .ZN(n752) );
  AND2_X1 U374 ( .A1(n520), .A2(n396), .ZN(n521) );
  XNOR2_X1 U375 ( .A(n399), .B(KEYINPUT102), .ZN(n520) );
  XNOR2_X1 U376 ( .A(n505), .B(n504), .ZN(n645) );
  NOR2_X1 U377 ( .A1(n752), .A2(n628), .ZN(n578) );
  XNOR2_X1 U378 ( .A(n459), .B(n458), .ZN(n525) );
  NOR2_X2 U379 ( .A1(n669), .A2(n412), .ZN(n542) );
  XNOR2_X2 U380 ( .A(n460), .B(KEYINPUT41), .ZN(n712) );
  OR2_X2 U381 ( .A1(n534), .A2(n533), .ZN(n536) );
  XNOR2_X2 U382 ( .A(n577), .B(KEYINPUT98), .ZN(n627) );
  XNOR2_X2 U383 ( .A(G143), .B(G128), .ZN(n360) );
  NOR2_X2 U384 ( .A1(n568), .A2(n691), .ZN(n582) );
  INV_X1 U385 ( .A(KEYINPUT85), .ZN(n392) );
  INV_X1 U386 ( .A(KEYINPUT4), .ZN(n416) );
  NOR2_X1 U387 ( .A1(n609), .A2(n606), .ZN(n603) );
  AND2_X1 U388 ( .A1(n544), .A2(n754), .ZN(n394) );
  XNOR2_X1 U389 ( .A(n378), .B(n567), .ZN(n628) );
  AND2_X1 U390 ( .A1(n538), .A2(KEYINPUT47), .ZN(n412) );
  XNOR2_X1 U391 ( .A(n572), .B(n571), .ZN(n713) );
  NOR2_X1 U392 ( .A1(n403), .A2(n408), .ZN(n375) );
  XOR2_X1 U393 ( .A(n531), .B(n530), .Z(n367) );
  INV_X1 U394 ( .A(n517), .ZN(n697) );
  XNOR2_X1 U395 ( .A(n469), .B(n468), .ZN(n619) );
  NAND2_X1 U396 ( .A1(n358), .A2(n359), .ZN(n462) );
  XNOR2_X1 U397 ( .A(n391), .B(n390), .ZN(n731) );
  XNOR2_X1 U398 ( .A(n392), .B(KEYINPUT3), .ZN(n391) );
  INV_X1 U399 ( .A(n416), .ZN(n357) );
  INV_X2 U400 ( .A(G953), .ZN(n743) );
  XNOR2_X1 U401 ( .A(G113), .B(G119), .ZN(n390) );
  XNOR2_X1 U402 ( .A(G143), .B(G128), .ZN(n453) );
  INV_X1 U403 ( .A(n704), .ZN(n352) );
  NAND2_X1 U404 ( .A1(n356), .A2(n357), .ZN(n359) );
  AND2_X1 U405 ( .A1(n506), .A2(n523), .ZN(n532) );
  AND2_X2 U406 ( .A1(n532), .A2(n367), .ZN(n672) );
  AND2_X1 U407 ( .A1(n386), .A2(n385), .ZN(n384) );
  AND2_X2 U408 ( .A1(n618), .A2(n718), .ZN(n353) );
  AND2_X2 U409 ( .A1(n618), .A2(n718), .ZN(n649) );
  NAND2_X1 U410 ( .A1(n372), .A2(n608), .ZN(n618) );
  XNOR2_X1 U411 ( .A(n477), .B(n354), .ZN(n355) );
  XOR2_X1 U412 ( .A(G119), .B(G128), .Z(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n480), .ZN(n366) );
  NAND2_X1 U414 ( .A1(n375), .A2(n511), .ZN(n527) );
  NAND2_X1 U415 ( .A1(n360), .A2(n416), .ZN(n358) );
  INV_X1 U416 ( .A(n453), .ZN(n356) );
  BUF_X1 U417 ( .A(n629), .Z(n361) );
  XNOR2_X1 U418 ( .A(n529), .B(n365), .ZN(n684) );
  NOR2_X2 U419 ( .A1(n570), .A2(n569), .ZN(n572) );
  NAND2_X1 U420 ( .A1(n697), .A2(n407), .ZN(n406) );
  AND2_X1 U421 ( .A1(n410), .A2(n528), .ZN(n407) );
  NAND2_X1 U422 ( .A1(n405), .A2(KEYINPUT30), .ZN(n404) );
  INV_X1 U423 ( .A(n509), .ZN(n409) );
  NOR2_X1 U424 ( .A1(n697), .A2(n410), .ZN(n408) );
  NAND2_X1 U425 ( .A1(n367), .A2(n362), .ZN(n558) );
  NAND2_X2 U426 ( .A1(n384), .A2(n381), .ZN(n523) );
  NAND2_X1 U427 ( .A1(G902), .A2(G469), .ZN(n385) );
  NOR2_X1 U428 ( .A1(G237), .A2(G953), .ZN(n442) );
  XOR2_X1 U429 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n433) );
  XNOR2_X1 U430 ( .A(G113), .B(G143), .ZN(n440) );
  INV_X1 U431 ( .A(KEYINPUT33), .ZN(n571) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n550) );
  INV_X1 U433 ( .A(KEYINPUT39), .ZN(n373) );
  NOR2_X1 U434 ( .A1(n527), .A2(n684), .ZN(n374) );
  NAND2_X1 U435 ( .A1(n383), .A2(n484), .ZN(n382) );
  INV_X1 U436 ( .A(G469), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U438 ( .A(n505), .B(n464), .ZN(n469) );
  INV_X1 U439 ( .A(KEYINPUT83), .ZN(n602) );
  NAND2_X1 U440 ( .A1(n683), .A2(n685), .ZN(n460) );
  NOR2_X1 U441 ( .A1(n549), .A2(n405), .ZN(n396) );
  NAND2_X1 U442 ( .A1(n406), .A2(n370), .ZN(n403) );
  BUF_X1 U443 ( .A(G953), .Z(n371) );
  XNOR2_X1 U444 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U445 ( .A(n499), .B(n498), .ZN(n503) );
  NOR2_X1 U446 ( .A1(n743), .A2(G952), .ZN(n655) );
  XNOR2_X1 U447 ( .A(n402), .B(KEYINPUT43), .ZN(n401) );
  XNOR2_X1 U448 ( .A(n388), .B(n363), .ZN(n513) );
  NAND2_X1 U449 ( .A1(n550), .A2(n518), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n574), .B(n380), .ZN(n376) );
  NAND2_X1 U451 ( .A1(n593), .A2(n377), .ZN(n378) );
  AND2_X1 U452 ( .A1(n566), .A2(n565), .ZN(n377) );
  XOR2_X1 U453 ( .A(n556), .B(KEYINPUT87), .Z(n362) );
  XOR2_X1 U454 ( .A(n512), .B(KEYINPUT40), .Z(n363) );
  XOR2_X1 U455 ( .A(n428), .B(KEYINPUT80), .Z(n364) );
  XOR2_X1 U456 ( .A(KEYINPUT75), .B(KEYINPUT38), .Z(n365) );
  AND2_X1 U457 ( .A1(n593), .A2(n565), .ZN(n368) );
  INV_X1 U458 ( .A(KEYINPUT30), .ZN(n410) );
  NOR2_X1 U459 ( .A1(n534), .A2(n525), .ZN(n369) );
  AND2_X1 U460 ( .A1(n409), .A2(n404), .ZN(n370) );
  INV_X1 U461 ( .A(n528), .ZN(n405) );
  NAND2_X1 U462 ( .A1(n604), .A2(n605), .ZN(n372) );
  NAND2_X1 U463 ( .A1(n376), .A2(n369), .ZN(n379) );
  INV_X1 U464 ( .A(KEYINPUT34), .ZN(n380) );
  NAND2_X1 U465 ( .A1(n645), .A2(G469), .ZN(n386) );
  XNOR2_X2 U466 ( .A(n523), .B(n522), .ZN(n568) );
  OR2_X1 U467 ( .A1(n645), .A2(n382), .ZN(n381) );
  INV_X1 U468 ( .A(n529), .ZN(n549) );
  XNOR2_X2 U469 ( .A(n429), .B(n364), .ZN(n529) );
  XNOR2_X1 U470 ( .A(n387), .B(n515), .ZN(n393) );
  NAND2_X1 U471 ( .A1(n389), .A2(n513), .ZN(n387) );
  INV_X1 U472 ( .A(n625), .ZN(n389) );
  XNOR2_X2 U473 ( .A(n508), .B(n507), .ZN(n625) );
  XNOR2_X2 U474 ( .A(n431), .B(KEYINPUT107), .ZN(n683) );
  NAND2_X1 U475 ( .A1(n394), .A2(n393), .ZN(n547) );
  XNOR2_X2 U476 ( .A(n395), .B(KEYINPUT108), .ZN(n754) );
  NAND2_X1 U477 ( .A1(n524), .A2(n575), .ZN(n395) );
  NAND2_X1 U478 ( .A1(n520), .A2(n528), .ZN(n397) );
  XNOR2_X1 U479 ( .A(n397), .B(KEYINPUT103), .ZN(n548) );
  XNOR2_X1 U480 ( .A(n603), .B(n602), .ZN(n604) );
  AND2_X1 U481 ( .A1(n398), .A2(n671), .ZN(n399) );
  XNOR2_X2 U482 ( .A(n518), .B(KEYINPUT100), .ZN(n671) );
  NOR2_X1 U483 ( .A1(n569), .A2(n519), .ZN(n398) );
  INV_X1 U484 ( .A(n569), .ZN(n592) );
  NAND2_X1 U485 ( .A1(n401), .A2(n549), .ZN(n400) );
  NAND2_X1 U486 ( .A1(n548), .A2(n568), .ZN(n402) );
  INV_X1 U487 ( .A(n513), .ZN(n751) );
  XNOR2_X2 U488 ( .A(n471), .B(n470), .ZN(n517) );
  AND2_X1 U489 ( .A1(G221), .A2(n481), .ZN(n411) );
  INV_X1 U490 ( .A(G107), .ZN(n496) );
  XNOR2_X1 U491 ( .A(n463), .B(G137), .ZN(n464) );
  XNOR2_X1 U492 ( .A(n497), .B(n496), .ZN(n499) );
  INV_X1 U493 ( .A(KEYINPUT63), .ZN(n623) );
  NAND2_X1 U494 ( .A1(n743), .A2(G224), .ZN(n414) );
  XNOR2_X2 U495 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n413) );
  XNOR2_X1 U496 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X2 U497 ( .A(G125), .B(G146), .ZN(n436) );
  XNOR2_X1 U498 ( .A(n415), .B(n436), .ZN(n418) );
  INV_X1 U499 ( .A(n462), .ZN(n417) );
  XNOR2_X1 U500 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U501 ( .A(G101), .B(KEYINPUT66), .ZN(n419) );
  XNOR2_X1 U502 ( .A(n419), .B(KEYINPUT67), .ZN(n501) );
  XNOR2_X1 U503 ( .A(n731), .B(n501), .ZN(n467) );
  XNOR2_X1 U504 ( .A(n420), .B(n467), .ZN(n426) );
  XNOR2_X1 U505 ( .A(KEYINPUT76), .B(G110), .ZN(n422) );
  INV_X1 U506 ( .A(G104), .ZN(n421) );
  XNOR2_X1 U507 ( .A(n422), .B(n421), .ZN(n500) );
  INV_X1 U508 ( .A(n500), .ZN(n423) );
  XNOR2_X1 U509 ( .A(n423), .B(KEYINPUT16), .ZN(n425) );
  XNOR2_X1 U510 ( .A(G122), .B(G116), .ZN(n424) );
  XNOR2_X1 U511 ( .A(n424), .B(G107), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n425), .B(n452), .ZN(n732) );
  XNOR2_X1 U513 ( .A(n426), .B(n732), .ZN(n650) );
  XNOR2_X1 U514 ( .A(G902), .B(KEYINPUT15), .ZN(n606) );
  NAND2_X1 U515 ( .A1(n650), .A2(n606), .ZN(n429) );
  INV_X1 U516 ( .A(G902), .ZN(n484) );
  INV_X1 U517 ( .A(G237), .ZN(n427) );
  NAND2_X1 U518 ( .A1(n484), .A2(n427), .ZN(n430) );
  NAND2_X1 U519 ( .A1(n430), .A2(G210), .ZN(n428) );
  NAND2_X1 U520 ( .A1(n430), .A2(G214), .ZN(n528) );
  OR2_X2 U521 ( .A1(n684), .A2(n405), .ZN(n431) );
  XNOR2_X1 U522 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n432) );
  XNOR2_X1 U523 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U524 ( .A(G104), .B(n434), .ZN(n439) );
  XNOR2_X1 U525 ( .A(G122), .B(G140), .ZN(n437) );
  INV_X1 U526 ( .A(KEYINPUT10), .ZN(n435) );
  XNOR2_X1 U527 ( .A(n436), .B(n435), .ZN(n482) );
  XNOR2_X1 U528 ( .A(n437), .B(n482), .ZN(n438) );
  XNOR2_X1 U529 ( .A(n439), .B(n438), .ZN(n446) );
  XOR2_X1 U530 ( .A(KEYINPUT11), .B(G131), .Z(n441) );
  XOR2_X1 U531 ( .A(n441), .B(n440), .Z(n444) );
  XNOR2_X1 U532 ( .A(n442), .B(KEYINPUT78), .ZN(n465) );
  NAND2_X1 U533 ( .A1(n465), .A2(G214), .ZN(n443) );
  XNOR2_X1 U534 ( .A(n446), .B(n445), .ZN(n639) );
  NAND2_X1 U535 ( .A1(n639), .A2(n484), .ZN(n448) );
  XNOR2_X1 U536 ( .A(KEYINPUT13), .B(G475), .ZN(n447) );
  XNOR2_X1 U537 ( .A(n448), .B(n447), .ZN(n534) );
  NAND2_X1 U538 ( .A1(G234), .A2(n743), .ZN(n449) );
  XOR2_X1 U539 ( .A(KEYINPUT8), .B(n449), .Z(n481) );
  NAND2_X1 U540 ( .A1(G217), .A2(n481), .ZN(n451) );
  XNOR2_X1 U541 ( .A(G134), .B(KEYINPUT9), .ZN(n450) );
  XNOR2_X1 U542 ( .A(n451), .B(n450), .ZN(n457) );
  INV_X1 U543 ( .A(n452), .ZN(n455) );
  XNOR2_X1 U544 ( .A(n360), .B(KEYINPUT7), .ZN(n454) );
  XNOR2_X1 U545 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U546 ( .A(n457), .B(n456), .ZN(n634) );
  NAND2_X1 U547 ( .A1(n634), .A2(n484), .ZN(n459) );
  INV_X1 U548 ( .A(G478), .ZN(n458) );
  AND2_X1 U549 ( .A1(n534), .A2(n525), .ZN(n685) );
  XNOR2_X1 U550 ( .A(G131), .B(G134), .ZN(n461) );
  XNOR2_X2 U551 ( .A(n462), .B(n461), .ZN(n739) );
  XNOR2_X2 U552 ( .A(n739), .B(G146), .ZN(n505) );
  XOR2_X1 U553 ( .A(KEYINPUT5), .B(G116), .Z(n463) );
  NAND2_X1 U554 ( .A1(n465), .A2(G210), .ZN(n466) );
  NAND2_X1 U555 ( .A1(n619), .A2(n484), .ZN(n471) );
  XNOR2_X1 U556 ( .A(G472), .B(KEYINPUT71), .ZN(n470) );
  NAND2_X1 U557 ( .A1(G234), .A2(G237), .ZN(n472) );
  XNOR2_X1 U558 ( .A(n472), .B(KEYINPUT14), .ZN(n473) );
  NAND2_X1 U559 ( .A1(G952), .A2(n473), .ZN(n711) );
  NOR2_X1 U560 ( .A1(n371), .A2(n711), .ZN(n555) );
  NAND2_X1 U561 ( .A1(G902), .A2(n473), .ZN(n553) );
  OR2_X1 U562 ( .A1(n743), .A2(n553), .ZN(n474) );
  XOR2_X1 U563 ( .A(KEYINPUT101), .B(n474), .Z(n475) );
  NOR2_X1 U564 ( .A1(G900), .A2(n475), .ZN(n476) );
  NOR2_X1 U565 ( .A1(n555), .A2(n476), .ZN(n509) );
  XOR2_X1 U566 ( .A(KEYINPUT88), .B(G110), .Z(n477) );
  XOR2_X1 U567 ( .A(KEYINPUT23), .B(KEYINPUT82), .Z(n479) );
  XNOR2_X1 U568 ( .A(KEYINPUT69), .B(KEYINPUT24), .ZN(n478) );
  XNOR2_X1 U569 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U570 ( .A(n366), .B(n411), .ZN(n483) );
  XOR2_X1 U571 ( .A(G137), .B(G140), .Z(n498) );
  XNOR2_X1 U572 ( .A(n482), .B(n498), .ZN(n742) );
  XNOR2_X1 U573 ( .A(n483), .B(n742), .ZN(n629) );
  NAND2_X1 U574 ( .A1(n629), .A2(n484), .ZN(n489) );
  NAND2_X1 U575 ( .A1(n606), .A2(G234), .ZN(n485) );
  XNOR2_X1 U576 ( .A(n485), .B(KEYINPUT20), .ZN(n490) );
  NAND2_X1 U577 ( .A1(n490), .A2(G217), .ZN(n487) );
  XNOR2_X1 U578 ( .A(KEYINPUT25), .B(KEYINPUT89), .ZN(n486) );
  XNOR2_X1 U579 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X2 U580 ( .A(n489), .B(n488), .ZN(n694) );
  NOR2_X1 U581 ( .A1(n509), .A2(n694), .ZN(n493) );
  XOR2_X1 U582 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n492) );
  NAND2_X1 U583 ( .A1(n490), .A2(G221), .ZN(n491) );
  XNOR2_X1 U584 ( .A(n492), .B(n491), .ZN(n693) );
  NAND2_X1 U585 ( .A1(n493), .A2(n693), .ZN(n519) );
  OR2_X1 U586 ( .A1(n517), .A2(n519), .ZN(n495) );
  INV_X1 U587 ( .A(KEYINPUT28), .ZN(n494) );
  XNOR2_X1 U588 ( .A(n495), .B(n494), .ZN(n506) );
  NAND2_X1 U589 ( .A1(G227), .A2(n743), .ZN(n497) );
  XNOR2_X1 U590 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U591 ( .A(n503), .B(n502), .ZN(n504) );
  NAND2_X1 U592 ( .A1(n712), .A2(n532), .ZN(n508) );
  INV_X1 U593 ( .A(KEYINPUT42), .ZN(n507) );
  XOR2_X1 U594 ( .A(n693), .B(KEYINPUT91), .Z(n559) );
  NAND2_X1 U595 ( .A1(n694), .A2(n559), .ZN(n691) );
  INV_X1 U596 ( .A(n691), .ZN(n510) );
  NAND2_X1 U597 ( .A1(n523), .A2(n510), .ZN(n585) );
  XNOR2_X1 U598 ( .A(KEYINPUT105), .B(n585), .ZN(n511) );
  INV_X1 U599 ( .A(n525), .ZN(n533) );
  INV_X2 U600 ( .A(n536), .ZN(n518) );
  INV_X1 U601 ( .A(KEYINPUT106), .ZN(n512) );
  INV_X1 U602 ( .A(KEYINPUT64), .ZN(n514) );
  XNOR2_X1 U603 ( .A(n514), .B(KEYINPUT46), .ZN(n515) );
  INV_X1 U604 ( .A(KEYINPUT6), .ZN(n516) );
  XNOR2_X1 U605 ( .A(n517), .B(n516), .ZN(n569) );
  XNOR2_X1 U606 ( .A(n521), .B(KEYINPUT36), .ZN(n524) );
  XNOR2_X1 U607 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n522) );
  INV_X1 U608 ( .A(n568), .ZN(n575) );
  NAND2_X1 U609 ( .A1(n369), .A2(n529), .ZN(n526) );
  NOR2_X1 U610 ( .A1(n527), .A2(n526), .ZN(n669) );
  NAND2_X1 U611 ( .A1(n529), .A2(n528), .ZN(n531) );
  INV_X1 U612 ( .A(KEYINPUT19), .ZN(n530) );
  NAND2_X1 U613 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U614 ( .A(n535), .B(KEYINPUT96), .ZN(n678) );
  NAND2_X1 U615 ( .A1(n678), .A2(n536), .ZN(n682) );
  AND2_X1 U616 ( .A1(n682), .A2(KEYINPUT74), .ZN(n537) );
  NAND2_X1 U617 ( .A1(n672), .A2(n537), .ZN(n538) );
  XOR2_X1 U618 ( .A(KEYINPUT74), .B(n682), .Z(n539) );
  NOR2_X1 U619 ( .A1(KEYINPUT47), .A2(n539), .ZN(n540) );
  NAND2_X1 U620 ( .A1(n672), .A2(n540), .ZN(n541) );
  NAND2_X1 U621 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U622 ( .A(n543), .B(KEYINPUT73), .ZN(n544) );
  INV_X1 U623 ( .A(KEYINPUT68), .ZN(n545) );
  XNOR2_X1 U624 ( .A(n545), .B(KEYINPUT48), .ZN(n546) );
  XNOR2_X1 U625 ( .A(n547), .B(n546), .ZN(n610) );
  INV_X1 U626 ( .A(n678), .ZN(n664) );
  AND2_X1 U627 ( .A1(n550), .A2(n664), .ZN(n681) );
  INV_X1 U628 ( .A(n681), .ZN(n611) );
  AND2_X1 U629 ( .A1(n753), .A2(n611), .ZN(n551) );
  NAND2_X1 U630 ( .A1(n610), .A2(n551), .ZN(n552) );
  XNOR2_X2 U631 ( .A(n552), .B(KEYINPUT84), .ZN(n716) );
  XNOR2_X1 U632 ( .A(n716), .B(KEYINPUT77), .ZN(n605) );
  XOR2_X1 U633 ( .A(G898), .B(KEYINPUT86), .Z(n728) );
  NAND2_X1 U634 ( .A1(n371), .A2(n728), .ZN(n734) );
  NOR2_X1 U635 ( .A1(n553), .A2(n734), .ZN(n554) );
  OR2_X1 U636 ( .A1(n555), .A2(n554), .ZN(n556) );
  INV_X1 U637 ( .A(KEYINPUT0), .ZN(n557) );
  XNOR2_X2 U638 ( .A(n558), .B(n557), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n685), .A2(n559), .ZN(n560) );
  XNOR2_X1 U640 ( .A(n560), .B(KEYINPUT97), .ZN(n561) );
  NAND2_X1 U641 ( .A1(n573), .A2(n561), .ZN(n564) );
  INV_X1 U642 ( .A(KEYINPUT72), .ZN(n562) );
  XNOR2_X1 U643 ( .A(n562), .B(KEYINPUT22), .ZN(n563) );
  XNOR2_X2 U644 ( .A(n564), .B(n563), .ZN(n593) );
  INV_X1 U645 ( .A(n694), .ZN(n565) );
  NOR2_X1 U646 ( .A1(n592), .A2(n568), .ZN(n566) );
  XNOR2_X1 U647 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n567) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT99), .ZN(n570) );
  NAND2_X1 U649 ( .A1(n713), .A2(n573), .ZN(n574) );
  NOR2_X1 U650 ( .A1(n697), .A2(n575), .ZN(n576) );
  NAND2_X1 U651 ( .A1(n368), .A2(n576), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n627), .ZN(n581) );
  INV_X1 U653 ( .A(KEYINPUT44), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n579), .A2(KEYINPUT70), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n581), .B(n580), .ZN(n600) );
  INV_X1 U656 ( .A(n573), .ZN(n586) );
  INV_X1 U657 ( .A(n697), .ZN(n588) );
  INV_X1 U658 ( .A(n582), .ZN(n583) );
  OR2_X1 U659 ( .A1(n588), .A2(n583), .ZN(n701) );
  NOR2_X1 U660 ( .A1(n586), .A2(n701), .ZN(n584) );
  XNOR2_X1 U661 ( .A(n584), .B(KEYINPUT31), .ZN(n677) );
  NOR2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U663 ( .A(KEYINPUT92), .B(n587), .ZN(n589) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n660) );
  NAND2_X1 U665 ( .A1(n677), .A2(n660), .ZN(n590) );
  NAND2_X1 U666 ( .A1(n590), .A2(n682), .ZN(n598) );
  NAND2_X1 U667 ( .A1(n568), .A2(n694), .ZN(n591) );
  NOR2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n594) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n658) );
  INV_X1 U670 ( .A(KEYINPUT70), .ZN(n595) );
  NAND2_X1 U671 ( .A1(n595), .A2(KEYINPUT44), .ZN(n596) );
  AND2_X1 U672 ( .A1(n658), .A2(n596), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X2 U674 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X2 U675 ( .A(n601), .B(KEYINPUT45), .ZN(n609) );
  INV_X1 U676 ( .A(n606), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n607), .A2(KEYINPUT2), .ZN(n608) );
  INV_X1 U678 ( .A(n609), .ZN(n617) );
  INV_X1 U679 ( .A(n610), .ZN(n615) );
  NAND2_X1 U680 ( .A1(n611), .A2(KEYINPUT2), .ZN(n612) );
  XNOR2_X1 U681 ( .A(n612), .B(KEYINPUT81), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n753), .A2(n613), .ZN(n614) );
  NOR2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n718) );
  NAND2_X1 U685 ( .A1(n353), .A2(G472), .ZN(n621) );
  XOR2_X1 U686 ( .A(KEYINPUT62), .B(n619), .Z(n620) );
  XNOR2_X1 U687 ( .A(n621), .B(n620), .ZN(n622) );
  NOR2_X2 U688 ( .A1(n622), .A2(n655), .ZN(n624) );
  XNOR2_X1 U689 ( .A(n624), .B(n623), .ZN(G57) );
  XOR2_X1 U690 ( .A(n625), .B(G137), .Z(G39) );
  XOR2_X1 U691 ( .A(G110), .B(KEYINPUT109), .Z(n626) );
  XNOR2_X1 U692 ( .A(n627), .B(n626), .ZN(G12) );
  XOR2_X1 U693 ( .A(n628), .B(G119), .Z(G21) );
  NAND2_X1 U694 ( .A1(n353), .A2(G217), .ZN(n631) );
  XNOR2_X1 U695 ( .A(n361), .B(KEYINPUT123), .ZN(n630) );
  XNOR2_X1 U696 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X2 U697 ( .A1(n632), .A2(n655), .ZN(n633) );
  XNOR2_X1 U698 ( .A(n633), .B(KEYINPUT124), .ZN(G66) );
  NAND2_X1 U699 ( .A1(n649), .A2(G478), .ZN(n636) );
  XNOR2_X1 U700 ( .A(n634), .B(KEYINPUT121), .ZN(n635) );
  XNOR2_X1 U701 ( .A(n636), .B(n635), .ZN(n637) );
  NOR2_X2 U702 ( .A1(n637), .A2(n655), .ZN(n638) );
  XNOR2_X1 U703 ( .A(n638), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U704 ( .A1(n649), .A2(G475), .ZN(n641) );
  XNOR2_X1 U705 ( .A(n639), .B(KEYINPUT59), .ZN(n640) );
  XNOR2_X1 U706 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X2 U707 ( .A1(n642), .A2(n655), .ZN(n643) );
  XNOR2_X1 U708 ( .A(n643), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U709 ( .A1(n649), .A2(G469), .ZN(n647) );
  XOR2_X1 U710 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X1 U713 ( .A1(n648), .A2(n655), .ZN(G54) );
  NAND2_X1 U714 ( .A1(n353), .A2(G210), .ZN(n654) );
  XNOR2_X1 U715 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n651) );
  XNOR2_X1 U716 ( .A(n651), .B(KEYINPUT55), .ZN(n652) );
  XNOR2_X1 U717 ( .A(n650), .B(n652), .ZN(n653) );
  XNOR2_X1 U718 ( .A(n654), .B(n653), .ZN(n656) );
  NOR2_X2 U719 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U720 ( .A(n657), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U721 ( .A(G101), .B(n658), .ZN(G3) );
  INV_X1 U722 ( .A(n671), .ZN(n675) );
  NOR2_X1 U723 ( .A1(n675), .A2(n660), .ZN(n659) );
  XOR2_X1 U724 ( .A(G104), .B(n659), .Z(G6) );
  NOR2_X1 U725 ( .A1(n678), .A2(n660), .ZN(n662) );
  XNOR2_X1 U726 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n661) );
  XNOR2_X1 U727 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U728 ( .A(G107), .B(n663), .ZN(G9) );
  XOR2_X1 U729 ( .A(KEYINPUT29), .B(KEYINPUT111), .Z(n666) );
  NAND2_X1 U730 ( .A1(n672), .A2(n664), .ZN(n665) );
  XNOR2_X1 U731 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U732 ( .A(G128), .B(KEYINPUT110), .Z(n667) );
  XNOR2_X1 U733 ( .A(n668), .B(n667), .ZN(G30) );
  XOR2_X1 U734 ( .A(G143), .B(n669), .Z(n670) );
  XNOR2_X1 U735 ( .A(KEYINPUT112), .B(n670), .ZN(G45) );
  XOR2_X1 U736 ( .A(G146), .B(KEYINPUT113), .Z(n674) );
  NAND2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n674), .B(n673), .ZN(G48) );
  NOR2_X1 U739 ( .A1(n675), .A2(n677), .ZN(n676) );
  XOR2_X1 U740 ( .A(G113), .B(n676), .Z(G15) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U742 ( .A(KEYINPUT114), .B(n679), .Z(n680) );
  XNOR2_X1 U743 ( .A(G116), .B(n680), .ZN(G18) );
  XOR2_X1 U744 ( .A(G134), .B(n681), .Z(G36) );
  NAND2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n688) );
  NAND2_X1 U746 ( .A1(n684), .A2(n405), .ZN(n686) );
  NAND2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U749 ( .A1(n713), .A2(n689), .ZN(n690) );
  XNOR2_X1 U750 ( .A(n690), .B(KEYINPUT117), .ZN(n707) );
  NAND2_X1 U751 ( .A1(n568), .A2(n691), .ZN(n692) );
  XNOR2_X1 U752 ( .A(KEYINPUT50), .B(n692), .ZN(n699) );
  NOR2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U754 ( .A(KEYINPUT49), .B(n695), .Z(n696) );
  NOR2_X1 U755 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U756 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U757 ( .A(n700), .B(KEYINPUT116), .ZN(n702) );
  NAND2_X1 U758 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U759 ( .A(KEYINPUT51), .B(n703), .ZN(n705) );
  INV_X1 U760 ( .A(n712), .ZN(n704) );
  NOR2_X1 U761 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U762 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n708), .B(KEYINPUT52), .ZN(n709) );
  XNOR2_X1 U764 ( .A(KEYINPUT118), .B(n709), .ZN(n710) );
  NOR2_X1 U765 ( .A1(n711), .A2(n710), .ZN(n715) );
  AND2_X1 U766 ( .A1(n713), .A2(n352), .ZN(n714) );
  NOR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(n723) );
  NOR2_X1 U768 ( .A1(n609), .A2(n716), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n717), .A2(KEYINPUT2), .ZN(n720) );
  INV_X1 U770 ( .A(n718), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n721), .A2(n371), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U774 ( .A(KEYINPUT119), .B(n724), .ZN(n725) );
  XNOR2_X1 U775 ( .A(KEYINPUT53), .B(n725), .ZN(G75) );
  NOR2_X1 U776 ( .A1(n609), .A2(n371), .ZN(n730) );
  NAND2_X1 U777 ( .A1(n371), .A2(G224), .ZN(n726) );
  XOR2_X1 U778 ( .A(KEYINPUT61), .B(n726), .Z(n727) );
  NOR2_X1 U779 ( .A1(n728), .A2(n727), .ZN(n729) );
  NOR2_X1 U780 ( .A1(n730), .A2(n729), .ZN(n737) );
  XOR2_X1 U781 ( .A(G101), .B(n731), .Z(n733) );
  XNOR2_X1 U782 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U784 ( .A(n737), .B(n736), .ZN(n738) );
  XOR2_X1 U785 ( .A(KEYINPUT125), .B(n738), .Z(G69) );
  BUF_X1 U786 ( .A(n739), .Z(n740) );
  XNOR2_X1 U787 ( .A(n740), .B(KEYINPUT126), .ZN(n741) );
  XOR2_X1 U788 ( .A(n742), .B(n741), .Z(n745) );
  XOR2_X1 U789 ( .A(n745), .B(n716), .Z(n744) );
  NAND2_X1 U790 ( .A1(n744), .A2(n743), .ZN(n750) );
  XOR2_X1 U791 ( .A(G227), .B(n745), .Z(n746) );
  NAND2_X1 U792 ( .A1(n746), .A2(G900), .ZN(n747) );
  NAND2_X1 U793 ( .A1(n371), .A2(n747), .ZN(n748) );
  XOR2_X1 U794 ( .A(KEYINPUT127), .B(n748), .Z(n749) );
  NAND2_X1 U795 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U796 ( .A(G131), .B(n751), .Z(G33) );
  XOR2_X1 U797 ( .A(G122), .B(n752), .Z(G24) );
  XNOR2_X1 U798 ( .A(G140), .B(n753), .ZN(G42) );
  XNOR2_X1 U799 ( .A(n754), .B(KEYINPUT37), .ZN(n755) );
  XNOR2_X1 U800 ( .A(n755), .B(KEYINPUT115), .ZN(n756) );
  XNOR2_X1 U801 ( .A(G125), .B(n756), .ZN(G27) );
endmodule

