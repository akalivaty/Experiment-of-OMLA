//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT65), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n220), .B(new_n221), .C1(G107), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G87), .ZN(new_n228));
  INV_X1    g0028(.A(G250), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n203), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n206), .B(new_n212), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G264), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n217), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  AND2_X1   g0049(.A1(G1), .A2(G13), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n224), .A2(G1698), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(G226), .B2(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G97), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n253), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(KEYINPUT67), .A3(new_n209), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n250), .B2(new_n251), .ZN(new_n268));
  OAI211_X1 g0068(.A(G274), .B(new_n264), .C1(new_n266), .C2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT67), .B1(new_n265), .B2(new_n209), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n250), .A2(new_n267), .A3(new_n251), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n262), .A2(new_n263), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(G1), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n273), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n272), .A2(G238), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n261), .A2(new_n269), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n281), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n261), .A2(new_n279), .A3(new_n269), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT14), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n293), .A3(G169), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n287), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n276), .A2(KEYINPUT68), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n274), .A2(G1), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(G13), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G68), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT12), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT69), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n304), .A2(new_n305), .A3(new_n209), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n304), .B2(new_n209), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n298), .A2(G20), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G68), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT77), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G20), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G50), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT76), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n301), .A2(G20), .ZN(new_n316));
  INV_X1    g0116(.A(G77), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n210), .A2(G33), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT11), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n306), .A2(new_n307), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n320), .B1(new_n319), .B2(new_n321), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n303), .B(new_n311), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n295), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n210), .A2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT8), .B(G58), .Z(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(KEYINPUT72), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT15), .B(G87), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n331), .B1(new_n210), .B2(new_n317), .C1(new_n318), .C2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n321), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n300), .A2(new_n317), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n308), .A2(G77), .A3(new_n309), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n278), .B(G244), .C1(new_n268), .C2(new_n266), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n269), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT70), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT70), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n341), .A3(new_n269), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n326), .ZN(new_n344));
  NAND2_X1  g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G1698), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G232), .ZN(new_n348));
  INV_X1    g0148(.A(G238), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n346), .B(new_n348), .C1(new_n349), .C2(new_n347), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n350), .B(new_n253), .C1(G107), .C2(new_n346), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n340), .A2(new_n342), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G169), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT71), .A4(new_n351), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n338), .A2(new_n341), .A3(new_n269), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n341), .B1(new_n338), .B2(new_n269), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT71), .B1(new_n360), .B2(new_n351), .ZN(new_n361));
  INV_X1    g0161(.A(new_n356), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n337), .B(new_n357), .C1(new_n363), .C2(G179), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n325), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT17), .ZN(new_n366));
  INV_X1    g0166(.A(G223), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n347), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n215), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(new_n255), .C2(new_n256), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n253), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n272), .A2(G232), .A3(new_n278), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n269), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT80), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n375), .A2(new_n376), .A3(G190), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT80), .ZN(new_n380));
  AND2_X1   g0180(.A1(new_n374), .A2(new_n269), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(new_n373), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n377), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n299), .A2(new_n329), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n308), .A2(new_n309), .ZN(new_n387));
  INV_X1    g0187(.A(new_n329), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n344), .A2(new_n210), .A3(new_n345), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT7), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n344), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n345), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(KEYINPUT79), .A3(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(G68), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n223), .A2(new_n301), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n312), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n392), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n255), .A2(new_n256), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT7), .B1(new_n407), .B2(new_n210), .ZN(new_n408));
  INV_X1    g0208(.A(new_n396), .ZN(new_n409));
  OAI21_X1  g0209(.A(G68), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n321), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n390), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n366), .B1(new_n384), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n399), .A2(new_n405), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n391), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n301), .B1(new_n395), .B2(new_n396), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n404), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n308), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n389), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n381), .A2(KEYINPUT80), .A3(new_n382), .A4(new_n373), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n376), .B1(new_n375), .B2(new_n378), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n375), .A2(G190), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n420), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n375), .A2(G169), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n290), .B2(new_n375), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n413), .A2(KEYINPUT18), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT18), .B1(new_n413), .B2(new_n427), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n414), .B(new_n425), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n365), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n347), .A2(G222), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n346), .B(new_n433), .C1(new_n367), .C2(new_n347), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n434), .B(new_n253), .C1(G77), .C2(new_n346), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n272), .A2(G226), .A3(new_n278), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(new_n269), .A3(new_n436), .ZN(new_n437));
  OR2_X1    g0237(.A1(new_n437), .A2(new_n382), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT73), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(G200), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT74), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n388), .A2(new_n318), .ZN(new_n445));
  NOR3_X1   g0245(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n446));
  INV_X1    g0246(.A(G150), .ZN(new_n447));
  OAI22_X1  g0247(.A1(new_n446), .A2(new_n210), .B1(new_n327), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n321), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n300), .A2(new_n214), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n449), .B(new_n450), .C1(new_n214), .C2(new_n387), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT9), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT10), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n444), .A2(KEYINPUT10), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n444), .A2(KEYINPUT10), .ZN(new_n455));
  INV_X1    g0255(.A(new_n452), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n455), .C1(new_n442), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n437), .A2(new_n355), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n451), .C1(G179), .C2(new_n437), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n453), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n289), .A2(new_n382), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n378), .B1(new_n282), .B2(new_n284), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n461), .A2(new_n324), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(G190), .B1(new_n361), .B2(new_n362), .ZN(new_n464));
  INV_X1    g0264(.A(new_n337), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n354), .A2(G200), .A3(new_n356), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NOR4_X1   g0268(.A1(new_n432), .A2(new_n460), .A3(new_n463), .A4(new_n468), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n210), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT22), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT22), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n346), .A2(new_n472), .A3(new_n210), .A4(G87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G116), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n471), .A2(new_n473), .B1(new_n210), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n210), .A2(G107), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT23), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n476), .A2(KEYINPUT24), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT24), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n298), .A2(G33), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n308), .A2(G107), .A3(new_n299), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G107), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n298), .A2(G13), .A3(G20), .A4(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT25), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(new_n486), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT85), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n483), .B(KEYINPUT85), .C1(new_n487), .C2(new_n488), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n481), .A2(new_n321), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g0293(.A(KEYINPUT5), .B(G41), .ZN(new_n494));
  AND3_X1   g0294(.A1(new_n298), .A2(new_n494), .A3(G45), .ZN(new_n495));
  INV_X1    g0295(.A(G274), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n270), .B2(new_n271), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n298), .A2(new_n494), .A3(G45), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(new_n272), .A3(G264), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n229), .A2(new_n347), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n226), .A2(G1698), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n502), .C1(new_n255), .C2(new_n256), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G294), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n253), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n498), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT86), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n498), .A2(new_n500), .A3(new_n506), .A4(KEYINPUT86), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n355), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n507), .A2(new_n290), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n493), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n509), .A2(new_n382), .A3(new_n510), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n507), .A2(new_n378), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT87), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT87), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n507), .A2(new_n518), .A3(new_n378), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n515), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n491), .A2(new_n492), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n476), .A2(new_n478), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT24), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n476), .A2(KEYINPUT24), .A3(new_n478), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n321), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT88), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n515), .A2(new_n517), .A3(new_n519), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT88), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n493), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n514), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n499), .A2(new_n272), .A3(G270), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G264), .A2(G1698), .ZN(new_n534));
  OAI221_X1 g0334(.A(new_n534), .B1(new_n226), .B2(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n535));
  INV_X1    g0335(.A(G303), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n407), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n537), .A3(new_n253), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n498), .A2(new_n533), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n498), .A2(new_n533), .A3(KEYINPUT83), .A4(new_n538), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(G200), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT84), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n300), .A2(new_n216), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n308), .A2(G116), .A3(new_n299), .A4(new_n482), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n304), .A2(new_n209), .B1(G20), .B2(new_n216), .ZN(new_n547));
  INV_X1    g0347(.A(G283), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n326), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n210), .B1(new_n225), .B2(G33), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT20), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n551), .A2(new_n552), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n545), .B(new_n546), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n543), .A2(new_n544), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n544), .B1(new_n543), .B2(new_n556), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n382), .B1(new_n541), .B2(new_n542), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n556), .A2(new_n290), .A3(new_n539), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n541), .A2(new_n555), .A3(G169), .A4(new_n542), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(KEYINPUT21), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(KEYINPUT21), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n346), .A2(G250), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n347), .B1(new_n568), .B2(KEYINPUT4), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT4), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n570), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n571), .B(G244), .C1(new_n256), .C2(new_n255), .ZN(new_n572));
  INV_X1    g0372(.A(new_n549), .ZN(new_n573));
  INV_X1    g0373(.A(G244), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n344), .B2(new_n345), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n572), .B(new_n573), .C1(new_n575), .C2(KEYINPUT4), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n253), .B1(new_n569), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n263), .B1(new_n296), .B2(new_n297), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(new_n494), .B1(new_n270), .B2(new_n271), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n579), .A2(G257), .B1(new_n495), .B2(new_n497), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G169), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n580), .A3(G179), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n397), .A2(G107), .A3(new_n398), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n484), .A2(KEYINPUT6), .A3(G97), .ZN(new_n586));
  XOR2_X1   g0386(.A(G97), .B(G107), .Z(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(KEYINPUT6), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT81), .B1(new_n327), .B2(new_n317), .ZN(new_n589));
  OR3_X1    g0389(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n317), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n588), .A2(G20), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n321), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n300), .A2(new_n225), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n308), .A2(new_n299), .A3(new_n482), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n225), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n308), .B1(new_n585), .B2(new_n591), .ZN(new_n600));
  OAI21_X1  g0400(.A(KEYINPUT82), .B1(new_n600), .B2(new_n597), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n584), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n597), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n581), .A2(G200), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n603), .B(new_n604), .C1(new_n382), .C2(new_n581), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n228), .A2(new_n225), .A3(new_n484), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(KEYINPUT19), .C1(G20), .C2(new_n260), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n210), .B(G68), .C1(new_n255), .C2(new_n256), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n259), .B2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n321), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n308), .A2(G87), .A3(new_n299), .A4(new_n482), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n300), .A2(new_n332), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n349), .A2(new_n347), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n574), .A2(G1698), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n617), .B(new_n618), .C1(new_n255), .C2(new_n256), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n252), .B1(new_n619), .B2(new_n474), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n578), .A2(new_n496), .B1(new_n270), .B2(new_n271), .ZN(new_n621));
  XNOR2_X1  g0421(.A(KEYINPUT68), .B(G1), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n229), .B1(new_n622), .B2(new_n263), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G190), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n616), .B(new_n625), .C1(new_n378), .C2(new_n624), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n623), .ZN(new_n627));
  INV_X1    g0427(.A(new_n620), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n355), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n624), .A2(new_n290), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n613), .B(new_n615), .C1(new_n332), .C2(new_n596), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n606), .A2(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n469), .A2(new_n532), .A3(new_n567), .A4(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n453), .A2(new_n457), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n365), .A2(new_n463), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n639), .A2(new_n414), .A3(new_n425), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n428), .A2(new_n429), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n642), .A2(new_n459), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n528), .A2(new_n531), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n541), .A2(new_n542), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT21), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n646), .A3(G169), .A4(new_n555), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n563), .A2(KEYINPUT21), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n561), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n527), .B1(new_n511), .B2(new_n512), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n606), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT89), .B1(new_n624), .B2(new_n378), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT89), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n298), .A2(G45), .A3(new_n496), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n623), .A2(new_n272), .A3(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n654), .B(G200), .C1(new_n656), .C2(new_n620), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n653), .A2(new_n616), .A3(new_n625), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n633), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n644), .A2(new_n651), .A3(new_n652), .A4(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n584), .A2(new_n599), .A3(new_n601), .ZN(new_n663));
  INV_X1    g0463(.A(new_n634), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n593), .A2(new_n598), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n584), .A2(new_n658), .A3(new_n633), .A4(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n633), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n665), .A2(new_n668), .A3(KEYINPUT90), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT90), .ZN(new_n670));
  INV_X1    g0470(.A(new_n633), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n577), .A2(G179), .A3(new_n580), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n355), .B1(new_n577), .B2(new_n580), .ZN(new_n673));
  OAI22_X1  g0473(.A1(new_n672), .A2(new_n673), .B1(new_n600), .B2(new_n597), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n659), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n675), .B2(new_n662), .ZN(new_n676));
  OAI21_X1  g0476(.A(KEYINPUT26), .B1(new_n602), .B2(new_n634), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n670), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n661), .B1(new_n669), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n469), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n643), .A2(new_n680), .ZN(G369));
  NAND2_X1  g0481(.A1(new_n210), .A2(G13), .ZN(new_n682));
  OR3_X1    g0482(.A1(new_n622), .A2(KEYINPUT27), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT27), .B1(new_n622), .B2(new_n682), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n683), .A2(new_n684), .A3(G213), .ZN(new_n685));
  INV_X1    g0485(.A(G343), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n532), .B1(new_n493), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n514), .A2(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n567), .A2(KEYINPUT91), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n555), .A2(new_n687), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT91), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n560), .B2(new_n566), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n649), .A2(new_n555), .A3(new_n687), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n691), .A2(new_n696), .A3(G330), .A4(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n650), .A2(new_n687), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n649), .A2(new_n687), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n699), .B1(new_n532), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n204), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n607), .A2(G116), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(G1), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n208), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n708), .B2(new_n705), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n606), .A2(KEYINPUT94), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n602), .A2(new_n712), .A3(new_n605), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n644), .A3(new_n651), .A4(new_n660), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n633), .B1(new_n675), .B2(new_n662), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n602), .A2(KEYINPUT26), .A3(new_n634), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n687), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n679), .A2(new_n688), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT93), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT90), .B1(new_n665), .B2(new_n668), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n675), .A2(new_n662), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(new_n677), .A3(new_n670), .A4(new_n633), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n687), .B1(new_n728), .B2(new_n661), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n721), .B1(new_n731), .B2(new_n720), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n532), .A2(new_n567), .A3(new_n635), .A4(new_n688), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n581), .A2(new_n541), .A3(new_n290), .A4(new_n542), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT92), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n629), .A2(new_n507), .ZN(new_n736));
  OR3_X1    g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n734), .B2(new_n736), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n583), .A2(new_n629), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n500), .A2(new_n506), .ZN(new_n741));
  INV_X1    g0541(.A(new_n539), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n741), .A4(new_n742), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n687), .B1(new_n739), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n734), .A2(new_n736), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT31), .B(new_n687), .C1(new_n747), .C2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n733), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n732), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n710), .B1(new_n756), .B2(G1), .ZN(G364));
  NAND3_X1  g0557(.A1(new_n696), .A2(G330), .A3(new_n697), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(KEYINPUT95), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n696), .A2(new_n697), .ZN(new_n760));
  INV_X1    g0560(.A(G330), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n759), .B(new_n762), .Z(new_n763));
  INV_X1    g0563(.A(new_n682), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G45), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n705), .A2(G1), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n210), .A2(new_n290), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT96), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(KEYINPUT96), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n768), .A2(new_n382), .A3(G200), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n772), .A2(new_n317), .B1(new_n301), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n382), .A2(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n769), .A2(new_n775), .A3(new_n770), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n774), .B1(G58), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n210), .A2(G179), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n382), .A3(G200), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n780), .A2(KEYINPUT97), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(KEYINPUT97), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n775), .A2(new_n290), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n784), .A2(G107), .B1(G97), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n382), .A2(new_n378), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n779), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n346), .B1(new_n789), .B2(new_n228), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n768), .A2(new_n788), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G50), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n779), .A2(new_n771), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT32), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n778), .A2(new_n787), .A3(new_n793), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(G326), .ZN(new_n799));
  XOR2_X1   g0599(.A(KEYINPUT33), .B(G317), .Z(new_n800));
  OAI221_X1 g0600(.A(new_n407), .B1(new_n791), .B2(new_n799), .C1(new_n773), .C2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n794), .B(KEYINPUT98), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n784), .A2(G283), .B1(new_n803), .B2(G329), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT99), .Z(new_n805));
  INV_X1    g0605(.A(new_n772), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n801), .B(new_n805), .C1(G311), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(G294), .ZN(new_n808));
  INV_X1    g0608(.A(new_n786), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(new_n808), .B2(new_n809), .C1(new_n536), .C2(new_n789), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n776), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n798), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n209), .B1(G20), .B2(new_n355), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n346), .A2(G355), .A3(new_n204), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n248), .A2(G45), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n703), .A2(new_n346), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n708), .B2(G45), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n816), .B1(G116), .B2(new_n204), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(G13), .A2(G33), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(G20), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n814), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n766), .B1(new_n760), .B2(new_n823), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n815), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n767), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G396));
  NAND2_X1  g0629(.A1(new_n337), .A2(new_n687), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n466), .A2(new_n465), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n382), .B1(new_n354), .B2(new_n356), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n364), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT102), .ZN(new_n835));
  AOI21_X1  g0635(.A(G179), .B1(new_n354), .B2(new_n356), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n355), .B2(new_n363), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n837), .A2(new_n337), .A3(new_n688), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n835), .B1(new_n834), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n724), .A2(new_n730), .A3(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n337), .A2(new_n837), .B1(new_n467), .B2(new_n830), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n364), .A2(new_n687), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT102), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n729), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n842), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n754), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n842), .A2(new_n754), .A3(new_n848), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n766), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n766), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n847), .A2(new_n822), .ZN(new_n855));
  INV_X1    g0655(.A(new_n789), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n784), .A2(G87), .B1(G107), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n225), .B2(new_n809), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n346), .B(new_n858), .C1(G303), .C2(new_n792), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n803), .A2(G311), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n777), .A2(G294), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n772), .A2(new_n216), .B1(new_n548), .B2(new_n773), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT100), .Z(new_n863));
  NAND4_X1  g0663(.A1(new_n859), .A2(new_n860), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n809), .A2(new_n223), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G143), .A2(new_n777), .B1(new_n806), .B2(G159), .ZN(new_n866));
  INV_X1    g0666(.A(new_n773), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n867), .A2(G150), .B1(new_n792), .B2(G137), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT34), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n783), .A2(new_n301), .B1(new_n802), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G50), .B2(new_n856), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n872), .A2(new_n346), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n864), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n814), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n814), .A2(new_n821), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n878), .B1(G77), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n854), .B1(new_n855), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n853), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT103), .ZN(G384));
  OAI21_X1  g0684(.A(new_n838), .B1(new_n722), .B2(new_n841), .ZN(new_n885));
  OR3_X1    g0685(.A1(new_n461), .A2(new_n324), .A3(new_n462), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n324), .A2(new_n687), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n293), .B1(new_n285), .B2(G169), .ZN(new_n888));
  AOI211_X1 g0688(.A(KEYINPUT14), .B(new_n355), .C1(new_n282), .C2(new_n284), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n888), .A2(new_n889), .A3(new_n291), .ZN(new_n890));
  INV_X1    g0690(.A(new_n324), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n886), .B(new_n887), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n324), .B(new_n687), .C1(new_n295), .C2(new_n463), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n685), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n391), .B1(new_n417), .B2(new_n404), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n411), .A3(new_n321), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n390), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n430), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n426), .B(new_n685), .C1(new_n290), .C2(new_n375), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n420), .A2(new_n424), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT37), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT105), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n898), .A2(new_n900), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n384), .B2(new_n413), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT37), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n420), .A2(new_n424), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n413), .A2(new_n427), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n413), .A2(new_n895), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n908), .A2(new_n909), .A3(new_n910), .A4(new_n902), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n903), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n899), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n899), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n885), .B(new_n894), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n899), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n916));
  XOR2_X1   g0716(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n917));
  INV_X1    g0717(.A(KEYINPUT107), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n911), .B(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n908), .A2(KEYINPUT106), .A3(new_n909), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n910), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT106), .B1(new_n908), .B2(new_n909), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT37), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n910), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n919), .A2(new_n923), .B1(new_n430), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n916), .B(new_n917), .C1(new_n925), .C2(KEYINPUT38), .ZN(new_n926));
  OAI21_X1  g0726(.A(KEYINPUT39), .B1(new_n914), .B2(new_n913), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n325), .A2(new_n687), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n641), .A2(new_n685), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n915), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n642), .A2(new_n459), .ZN(new_n934));
  INV_X1    g0734(.A(new_n721), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n723), .B(new_n687), .C1(new_n728), .C2(new_n661), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n935), .B1(new_n938), .B2(KEYINPUT29), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n934), .B1(new_n939), .B2(new_n469), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n933), .B(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  OAI211_X1 g0742(.A(KEYINPUT31), .B(new_n687), .C1(new_n739), .C2(new_n747), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n733), .A2(new_n750), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n847), .A2(new_n944), .A3(new_n894), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n914), .A2(new_n913), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n916), .B1(new_n925), .B2(KEYINPUT38), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n892), .A2(new_n893), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(new_n846), .B2(new_n845), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT40), .A4(new_n944), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n469), .A2(new_n944), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n952), .B(new_n953), .Z(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(new_n761), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n941), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n298), .B2(new_n764), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n588), .B(KEYINPUT104), .Z(new_n958));
  AOI21_X1  g0758(.A(new_n216), .B1(new_n958), .B2(KEYINPUT35), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n959), .B(new_n211), .C1(KEYINPUT35), .C2(new_n958), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT36), .ZN(new_n961));
  INV_X1    g0761(.A(G13), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n708), .A2(new_n317), .A3(new_n400), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n301), .A2(G50), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n962), .B(new_n622), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n957), .A2(new_n961), .A3(new_n965), .ZN(G367));
  NAND2_X1  g0766(.A1(new_n666), .A2(new_n687), .ZN(new_n967));
  AND3_X1   g0767(.A1(new_n602), .A2(new_n712), .A3(new_n605), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n712), .B1(new_n602), .B2(new_n605), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n674), .A2(new_n688), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n493), .A2(new_n530), .A3(new_n529), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n530), .B1(new_n493), .B2(new_n529), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n650), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n566), .A2(new_n688), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT42), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n688), .A2(new_n616), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n660), .A2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n633), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n971), .B1(new_n714), .B2(new_n967), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n602), .B1(new_n987), .B2(new_n650), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n688), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n981), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n986), .B1(new_n981), .B2(new_n989), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n698), .A2(new_n987), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n996), .B(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n704), .B(KEYINPUT41), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT44), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n973), .A2(new_n701), .A3(KEYINPUT110), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT110), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n699), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n976), .B2(new_n977), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1003), .B1(new_n987), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1001), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT45), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n987), .B2(new_n1005), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n973), .A2(new_n701), .A3(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT110), .B1(new_n973), .B2(new_n701), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n987), .A2(new_n1005), .A3(new_n1003), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(KEYINPUT44), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1007), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(KEYINPUT111), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n698), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT111), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1007), .A2(new_n1018), .A3(new_n1011), .A4(new_n1014), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT112), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n691), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n758), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n698), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n700), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n698), .A3(new_n977), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1027), .A2(new_n754), .A3(new_n732), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT112), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1016), .A2(new_n1030), .A3(new_n1017), .A4(new_n1019), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1021), .A2(new_n1029), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1000), .B1(new_n1033), .B2(new_n756), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n765), .A2(G1), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n998), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n794), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n777), .A2(G150), .B1(G137), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(G143), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1038), .B1(new_n223), .B2(new_n789), .C1(new_n1039), .C2(new_n791), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G50), .B2(new_n806), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n407), .B1(new_n867), .B2(G159), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n784), .A2(G77), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n809), .A2(new_n301), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n784), .A2(G97), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n484), .B2(new_n809), .C1(new_n548), .C2(new_n772), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n346), .B(new_n1048), .C1(G294), .C2(new_n867), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n856), .A2(G116), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT46), .ZN(new_n1051));
  INV_X1    g0851(.A(G311), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n776), .A2(new_n536), .B1(new_n1052), .B2(new_n791), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT113), .Z(new_n1054));
  NAND3_X1  g0854(.A1(new_n1049), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(G317), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n794), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1046), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT47), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n814), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n818), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n824), .B1(new_n204), .B2(new_n332), .C1(new_n240), .C2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n854), .A3(new_n1062), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n985), .A2(G20), .A3(new_n822), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1036), .A2(new_n1066), .ZN(G387));
  NAND2_X1  g0867(.A1(new_n1027), .A2(new_n1035), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n789), .A2(new_n317), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n346), .B1(new_n388), .B2(new_n773), .C1(new_n776), .C2(new_n214), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G150), .C2(new_n1037), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n806), .A2(G68), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n332), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G159), .A2(new_n792), .B1(new_n786), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1071), .A2(new_n1047), .A3(new_n1072), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n777), .A2(G317), .B1(G311), .B2(new_n867), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n536), .B2(new_n772), .C1(new_n811), .C2(new_n791), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT48), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n548), .B2(new_n809), .C1(new_n808), .C2(new_n789), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT49), .Z(new_n1080));
  OAI221_X1 g0880(.A(new_n407), .B1(new_n799), .B2(new_n794), .C1(new_n783), .C2(new_n216), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT115), .Z(new_n1082));
  OAI21_X1  g0882(.A(new_n1075), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n814), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n818), .B1(new_n237), .B2(new_n263), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n706), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1086), .A2(new_n204), .A3(new_n346), .ZN(new_n1087));
  AOI211_X1 g0887(.A(G45), .B(new_n1086), .C1(G68), .C2(G77), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n329), .A2(new_n214), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1090));
  XNOR2_X1  g0890(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1085), .A2(new_n1087), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n204), .A2(G107), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n824), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n766), .B1(new_n1022), .B2(new_n823), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1084), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n704), .B1(new_n756), .B2(new_n1027), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1068), .B(new_n1096), .C1(new_n1097), .C2(new_n1029), .ZN(G393));
  NAND2_X1  g0898(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1032), .A2(new_n1035), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n987), .A2(new_n823), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n346), .B1(new_n1037), .B2(G322), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n1102), .B1(new_n548), .B2(new_n789), .C1(new_n783), .C2(new_n484), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n786), .A2(G116), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n776), .A2(new_n1052), .B1(new_n1056), .B2(new_n791), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n806), .A2(G294), .B1(G303), .B2(new_n867), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n776), .A2(new_n795), .B1(new_n447), .B2(new_n791), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT51), .Z(new_n1111));
  OAI22_X1  g0911(.A1(new_n789), .A2(new_n301), .B1(new_n794), .B2(new_n1039), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(KEYINPUT116), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n784), .B2(G87), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(KEYINPUT116), .B2(new_n1112), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n772), .A2(new_n388), .B1(new_n809), .B2(new_n317), .ZN(new_n1116));
  OR4_X1    g0916(.A1(new_n407), .A2(new_n1111), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n773), .A2(new_n214), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1109), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n814), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n244), .A2(new_n818), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n824), .C1(new_n225), .C2(new_n204), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1101), .A2(new_n854), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1100), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n698), .B1(new_n1015), .B2(KEYINPUT111), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1030), .B1(new_n1127), .B2(new_n1019), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(new_n1028), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1032), .A2(new_n1099), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1126), .A2(new_n1129), .B1(new_n1028), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1124), .B1(new_n1131), .B2(new_n704), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G390));
  AOI22_X1  g0933(.A1(new_n784), .A2(G68), .B1(new_n803), .B2(G294), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n806), .A2(G97), .B1(G77), .B2(new_n786), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1134), .B(new_n1135), .C1(new_n484), .C2(new_n773), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n776), .A2(new_n216), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n791), .A2(new_n548), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n407), .B1(new_n789), .B2(new_n228), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT118), .Z(new_n1140));
  NOR4_X1   g0940(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n803), .A2(G125), .B1(G159), .B2(new_n786), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n784), .A2(G50), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n789), .A2(new_n447), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n792), .A2(G128), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT54), .B(G143), .Z(new_n1148));
  AND2_X1   g0948(.A1(new_n806), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n867), .A2(G137), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n346), .B1(new_n776), .B2(new_n873), .ZN(new_n1151));
  NOR4_X1   g0951(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n814), .B1(new_n1141), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1153), .B(new_n854), .C1(new_n329), .C2(new_n880), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n928), .C2(new_n822), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n953), .A2(G330), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n469), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n643), .B(new_n1160), .C1(new_n1161), .C2(new_n732), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n949), .B1(new_n754), .B2(new_n841), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n847), .A2(new_n944), .A3(G330), .A4(new_n894), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n885), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n850), .A2(new_n847), .A3(new_n894), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n844), .B1(new_n719), .B2(new_n847), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n847), .A2(G330), .A3(new_n944), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n949), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n929), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n948), .B(new_n1174), .C1(new_n1168), .C2(new_n949), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1167), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n929), .B1(new_n885), .B2(new_n894), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1175), .B(new_n1176), .C1(new_n1177), .C2(new_n928), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT39), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n899), .A2(new_n912), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT38), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1179), .B1(new_n1182), .B2(new_n916), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n430), .A2(new_n924), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n920), .A2(new_n910), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n922), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n902), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n911), .B(KEYINPUT107), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1184), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n914), .B1(new_n1189), .B2(new_n1181), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1183), .B1(new_n1190), .B2(new_n917), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n844), .B1(new_n729), .B2(new_n847), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1174), .B1(new_n1192), .B2(new_n949), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n719), .A2(new_n847), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n838), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n894), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1190), .A2(new_n929), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1191), .A2(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1164), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1178), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n705), .B1(new_n1173), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n949), .B1(new_n848), .B2(new_n838), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1191), .B1(new_n1202), .B2(new_n929), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n1203), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1199), .B1(new_n1203), .B2(new_n1175), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1166), .A2(new_n1171), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n940), .A2(new_n1207), .A3(new_n1160), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1159), .B1(new_n1201), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1035), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n1206), .ZN(G378));
  XOR2_X1   g1012(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n460), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n451), .A2(new_n895), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1213), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n453), .A2(new_n457), .A3(new_n459), .A4(new_n1217), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1214), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n821), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n880), .A2(G50), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n783), .A2(new_n223), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n407), .B1(new_n317), .B2(new_n789), .C1(new_n772), .C2(new_n332), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(G283), .C2(new_n803), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n262), .B1(new_n773), .B2(new_n225), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1228), .B(new_n1044), .C1(G116), .C2(new_n792), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1227), .B(new_n1229), .C1(new_n484), .C2(new_n776), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT120), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(new_n1231), .B(KEYINPUT58), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n214), .B1(new_n255), .B2(G41), .ZN(new_n1233));
  INV_X1    g1033(.A(G124), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n326), .B1(new_n794), .B2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n777), .A2(G128), .B1(new_n856), .B2(new_n1148), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n806), .A2(G137), .B1(G125), .B2(new_n792), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1238), .B1(new_n873), .B2(new_n773), .C1(new_n447), .C2(new_n809), .ZN(new_n1239));
  AOI211_X1 g1039(.A(G41), .B(new_n1235), .C1(new_n1239), .C2(KEYINPUT59), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(KEYINPUT59), .B2(new_n1239), .C1(new_n795), .C2(new_n783), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1232), .A2(new_n1233), .A3(new_n1241), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n766), .B(new_n1224), .C1(new_n1242), .C2(new_n814), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1223), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT121), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n947), .A2(new_n951), .A3(G330), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1222), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1221), .A2(new_n947), .A3(G330), .A4(new_n951), .ZN(new_n1248));
  AND4_X1   g1048(.A1(new_n1245), .A2(new_n1247), .A3(new_n932), .A4(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1248), .A2(new_n1247), .B1(new_n932), .B2(new_n1245), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1244), .B1(new_n1251), .B2(new_n1035), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1162), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1254), .B2(new_n1251), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n933), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1247), .A2(new_n932), .A3(new_n1248), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(KEYINPUT57), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1162), .B1(new_n1200), .B2(new_n1207), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n704), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1252), .B1(new_n1255), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT122), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT122), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(new_n1252), .C1(new_n1255), .C2(new_n1261), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1263), .A2(new_n1265), .ZN(G375));
  NAND2_X1  g1066(.A1(new_n1162), .A2(new_n1172), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1208), .A3(new_n999), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n407), .B1(new_n803), .B2(G128), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n806), .A2(G150), .B1(G159), .B2(new_n856), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(new_n223), .C2(new_n783), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n777), .A2(G137), .B1(new_n867), .B2(new_n1148), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n873), .B2(new_n791), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(KEYINPUT123), .Z(new_n1274));
  AOI211_X1 g1074(.A(new_n1271), .B(new_n1274), .C1(G50), .C2(new_n786), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n803), .A2(G303), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n346), .B1(new_n806), .B2(G107), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n867), .A2(G116), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1043), .A2(new_n1276), .A3(new_n1277), .A4(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n789), .A2(new_n225), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n776), .A2(new_n548), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n809), .A2(new_n332), .B1(new_n791), .B2(new_n808), .ZN(new_n1282));
  NOR4_X1   g1082(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .A4(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n814), .B1(new_n1275), .B2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1284), .B(new_n854), .C1(new_n822), .C2(new_n894), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n301), .B2(new_n879), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1207), .B2(new_n1035), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1268), .A2(new_n1287), .ZN(G381));
  AND3_X1   g1088(.A1(new_n1036), .A2(new_n1066), .A3(new_n1132), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(G384), .A2(G381), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1206), .A2(new_n1211), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n1159), .B(new_n1293), .C1(new_n1201), .C2(new_n1209), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1263), .A2(new_n1294), .A3(new_n1265), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1292), .A2(new_n1295), .ZN(G407));
  AND2_X1   g1096(.A1(new_n1292), .A2(G343), .ZN(new_n1297));
  OAI21_X1  g1097(.A(G213), .B1(new_n1297), .B2(new_n1295), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT124), .ZN(G409));
  AOI21_X1  g1099(.A(new_n1132), .B1(new_n1036), .B2(new_n1066), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(G393), .B(new_n828), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1289), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1301), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n997), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n996), .B(new_n1304), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1125), .A2(new_n1028), .A3(new_n1128), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n999), .B1(new_n1306), .B2(new_n755), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1305), .B1(new_n1307), .B2(new_n1211), .ZN(new_n1308));
  OAI21_X1  g1108(.A(G390), .B1(new_n1308), .B2(new_n1065), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1036), .A2(new_n1066), .A3(new_n1132), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1303), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  OR2_X1    g1111(.A1(new_n1302), .A2(new_n1311), .ZN(new_n1312));
  AOI22_X1  g1112(.A1(new_n1262), .A2(G378), .B1(G213), .B2(new_n686), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1162), .A2(new_n1172), .A3(KEYINPUT60), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n704), .A3(new_n1208), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1172), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1287), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  OR2_X1    g1117(.A1(new_n1317), .A2(G384), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(G384), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1244), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1254), .A2(new_n1251), .A3(new_n999), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1257), .A2(new_n1035), .A3(new_n1258), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1294), .A2(new_n1321), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1313), .A2(new_n1320), .A3(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT63), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1312), .A2(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n686), .A2(G213), .A3(G2897), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1318), .A2(new_n1319), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1313), .A2(KEYINPUT125), .A3(new_n1324), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT125), .B1(new_n1313), .B2(new_n1324), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT61), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1328), .A2(new_n1335), .A3(new_n1336), .A4(new_n1337), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1313), .A2(new_n1324), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT61), .B1(new_n1332), .B2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1325), .A2(KEYINPUT62), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1339), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1312), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1338), .A2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(new_n1262), .A2(G378), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1295), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1320), .A2(KEYINPUT126), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1302), .A2(new_n1311), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1295), .A2(new_n1348), .A3(new_n1346), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1350), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT127), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1350), .A2(new_n1352), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1312), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1350), .A2(new_n1351), .A3(KEYINPUT127), .A4(new_n1352), .ZN(new_n1358));
  AND3_X1   g1158(.A1(new_n1355), .A2(new_n1357), .A3(new_n1358), .ZN(G402));
endmodule


