//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT11), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n188), .A3(G134), .ZN(new_n193));
  AOI211_X1 g007(.A(G131), .B(new_n189), .C1(new_n191), .C2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n193), .ZN(new_n196));
  INV_X1    g010(.A(new_n189), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT3), .B1(new_n200), .B2(G107), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  INV_X1    g016(.A(G107), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G104), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(G107), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n201), .A2(new_n204), .A3(new_n205), .A4(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT83), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n206), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n200), .A2(G107), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n217), .B2(G146), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(KEYINPUT84), .ZN(new_n221));
  OAI21_X1  g035(.A(G128), .B1(new_n220), .B2(KEYINPUT84), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n226));
  AND4_X1   g040(.A1(new_n224), .A2(new_n226), .A3(new_n216), .A4(new_n218), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n224), .B1(new_n228), .B2(new_n226), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n223), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n214), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n216), .A3(new_n218), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n224), .A3(new_n226), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n225), .A2(KEYINPUT66), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G128), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n233), .A2(new_n234), .B1(new_n219), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n213), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n199), .B1(new_n231), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n187), .B1(new_n241), .B2(KEYINPUT12), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OR2_X1    g057(.A1(new_n241), .A2(KEYINPUT12), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n187), .A3(KEYINPUT12), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n238), .A2(new_n219), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n247), .B1(new_n229), .B2(new_n227), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n214), .A2(KEYINPUT10), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n231), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n201), .A2(new_n204), .A3(new_n206), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G101), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n209), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT4), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT0), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n225), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n219), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n228), .B1(new_n260), .B2(new_n225), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI211_X1 g079(.A(new_n249), .B(new_n251), .C1(new_n259), .C2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(new_n195), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n246), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(G110), .B(G140), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n272), .A2(G227), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n271), .B(new_n273), .Z(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n268), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n269), .A2(new_n277), .A3(new_n274), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(G469), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G469), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n274), .B1(new_n266), .B2(new_n268), .ZN(new_n282));
  INV_X1    g096(.A(new_n245), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(new_n242), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n284), .B2(new_n244), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n274), .B1(new_n269), .B2(new_n277), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n280), .B(new_n281), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n280), .A2(new_n281), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(KEYINPUT9), .B(G234), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G221), .B1(new_n292), .B2(G902), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT20), .ZN(new_n295));
  INV_X1    g109(.A(G125), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n296), .A2(KEYINPUT16), .A3(G140), .ZN(new_n297));
  XNOR2_X1  g111(.A(G125), .B(G140), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(KEYINPUT16), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(new_n215), .ZN(new_n300));
  INV_X1    g114(.A(G237), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(new_n272), .A3(G214), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT91), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n302), .A2(new_n303), .A3(G143), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n217), .A2(KEYINPUT91), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n305), .A2(new_n306), .A3(G214), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n195), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT95), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT17), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n310), .B(KEYINPUT95), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n309), .A2(new_n195), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT94), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n300), .B(new_n313), .C1(new_n317), .C2(KEYINPUT17), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n298), .B(new_n215), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n309), .A2(KEYINPUT93), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT18), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n320), .B1(new_n321), .B2(new_n195), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT92), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n322), .B1(new_n323), .B2(new_n309), .ZN(new_n324));
  NOR4_X1   g138(.A1(new_n320), .A2(KEYINPUT92), .A3(new_n321), .A4(new_n195), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n319), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G113), .B(G122), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(new_n200), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n299), .A2(G146), .ZN(new_n332));
  XOR2_X1   g146(.A(new_n298), .B(KEYINPUT19), .Z(new_n333));
  OAI211_X1 g147(.A(new_n317), .B(new_n332), .C1(G146), .C2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT96), .B1(new_n334), .B2(new_n326), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(new_n329), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(KEYINPUT96), .A3(new_n326), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n295), .B1(new_n338), .B2(KEYINPUT97), .ZN(new_n339));
  INV_X1    g153(.A(G475), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n334), .A2(KEYINPUT96), .A3(new_n326), .ZN(new_n341));
  NOR3_X1   g155(.A1(new_n341), .A2(new_n335), .A3(new_n329), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n340), .B(new_n281), .C1(new_n342), .C2(new_n331), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT97), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n342), .B2(new_n331), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n334), .A2(new_n326), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT96), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n330), .A3(new_n337), .ZN(new_n350));
  INV_X1    g164(.A(new_n331), .ZN(new_n351));
  AOI21_X1  g165(.A(G475), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n346), .A2(new_n352), .A3(new_n295), .A4(new_n281), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n344), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(G234), .A2(G237), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(G952), .A3(new_n272), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  XOR2_X1   g171(.A(KEYINPUT21), .B(G898), .Z(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(G902), .A3(G953), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT98), .ZN(new_n364));
  OR2_X1    g178(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT66), .B(G128), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n365), .B(new_n366), .C1(new_n367), .C2(new_n217), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G134), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n217), .A2(G128), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n370), .B1(new_n367), .B2(new_n217), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n369), .B(new_n371), .ZN(new_n372));
  AND2_X1   g186(.A1(KEYINPUT67), .A2(G116), .ZN(new_n373));
  NOR2_X1   g187(.A1(KEYINPUT67), .A2(G116), .ZN(new_n374));
  OAI21_X1  g188(.A(G122), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G116), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(G122), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(G107), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n372), .A2(new_n378), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n371), .B(G134), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT14), .B(G122), .C1(new_n373), .C2(new_n374), .ZN(new_n381));
  OAI211_X1 g195(.A(G107), .B(new_n381), .C1(new_n377), .C2(KEYINPUT14), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n380), .B(new_n382), .C1(G107), .C2(new_n377), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G217), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n292), .A2(new_n385), .A3(G953), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT99), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n379), .A2(new_n383), .A3(new_n386), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n384), .A2(KEYINPUT99), .A3(new_n387), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(new_n281), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT15), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n394), .A2(KEYINPUT100), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(KEYINPUT100), .ZN(new_n396));
  OAI21_X1  g210(.A(G478), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n393), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n327), .B(new_n330), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n340), .B1(new_n399), .B2(new_n281), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n354), .A2(new_n363), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT101), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G214), .B1(G237), .B2(G902), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT68), .ZN(new_n407));
  OAI21_X1  g221(.A(G119), .B1(new_n373), .B2(new_n374), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n376), .A2(G119), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G113), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT2), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT2), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G113), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n408), .A2(new_n410), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n408), .B2(new_n410), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n407), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n415), .ZN(new_n419));
  INV_X1    g233(.A(G119), .ZN(new_n420));
  OR2_X1    g234(.A1(KEYINPUT67), .A2(G116), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT67), .A2(G116), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n419), .B1(new_n423), .B2(new_n409), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n408), .A2(new_n410), .A3(new_n415), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT68), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n408), .A2(KEYINPUT5), .A3(new_n410), .ZN(new_n428));
  OAI21_X1  g242(.A(G113), .B1(new_n410), .B2(KEYINPUT5), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n416), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n258), .A2(new_n427), .B1(new_n214), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(G110), .B(G122), .Z(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n434), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n263), .A2(new_n264), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G125), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n440), .B1(new_n239), .B2(G125), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT87), .B(G224), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n272), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n432), .A2(new_n436), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT6), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR4_X1   g262(.A1(new_n432), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n436), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n438), .B(new_n444), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT88), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n433), .A2(new_n447), .A3(new_n434), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT86), .ZN(new_n453));
  INV_X1    g267(.A(new_n449), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n444), .A4(new_n438), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n441), .B(new_n458), .Z(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n432), .B2(new_n436), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n434), .B(KEYINPUT8), .Z(new_n461));
  NAND2_X1  g275(.A1(new_n213), .A2(new_n431), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n428), .B(KEYINPUT89), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n429), .B(KEYINPUT90), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n416), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n461), .B(new_n462), .C1(new_n465), .C2(new_n213), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n451), .A2(new_n457), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n451), .A2(new_n457), .A3(new_n469), .A4(new_n467), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n406), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n404), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n235), .A2(new_n237), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(G119), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT23), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n420), .B2(G128), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n420), .A2(G128), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n476), .A2(KEYINPUT78), .A3(KEYINPUT23), .A4(G119), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n300), .B1(new_n484), .B2(G110), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT77), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n477), .A2(new_n486), .A3(new_n481), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n486), .B1(new_n477), .B2(new_n481), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT24), .B(G110), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n298), .A2(new_n215), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n332), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n490), .B1(new_n487), .B2(new_n488), .ZN(new_n494));
  INV_X1    g308(.A(G110), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n479), .A2(new_n495), .A3(new_n482), .A4(new_n483), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(KEYINPUT79), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT79), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n499), .B(new_n493), .C1(new_n494), .C2(new_n496), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n491), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT80), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT22), .Z(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(G137), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n504), .B(new_n188), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(new_n491), .C1(new_n498), .C2(new_n500), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n281), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(KEYINPUT25), .A3(new_n281), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n385), .B1(G234), .B2(new_n281), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT81), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n509), .A2(new_n514), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(G101), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n307), .A2(G210), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT69), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT64), .B1(new_n188), .B2(G134), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT64), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(new_n190), .A3(G137), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n188), .A2(G134), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G131), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n192), .B1(G134), .B2(new_n188), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n190), .A2(KEYINPUT11), .A3(G137), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n195), .B(new_n197), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  AND2_X1   g349(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n268), .A2(new_n439), .B1(new_n536), .B2(new_n248), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n416), .A2(new_n417), .A3(new_n407), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT68), .B1(new_n424), .B2(new_n425), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n526), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n532), .A2(new_n535), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n199), .A2(new_n265), .B1(new_n239), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n543), .A2(new_n427), .A3(KEYINPUT69), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n525), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT70), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n543), .B(KEYINPUT30), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n427), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n537), .A2(new_n526), .A3(new_n540), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT69), .B1(new_n543), .B2(new_n427), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT70), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n525), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n546), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n546), .A2(new_n556), .A3(new_n548), .A4(new_n553), .ZN(new_n557));
  INV_X1    g371(.A(new_n525), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT72), .B1(new_n537), .B2(new_n540), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n543), .A2(new_n562), .A3(new_n427), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n564), .B2(new_n551), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT28), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n543), .B2(new_n427), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n558), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n555), .A2(new_n557), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(G472), .A2(G902), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n570), .A2(KEYINPUT32), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT32), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n571), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT32), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n576), .A2(KEYINPUT75), .A3(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n541), .A2(new_n544), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n561), .A2(new_n563), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n559), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n525), .A3(new_n567), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT29), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n548), .A2(new_n551), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n558), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT73), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n582), .A2(KEYINPUT73), .A3(new_n585), .A4(new_n583), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n549), .A2(new_n550), .B1(new_n427), .B2(new_n543), .ZN(new_n590));
  OAI211_X1 g404(.A(KEYINPUT29), .B(new_n567), .C1(new_n590), .C2(new_n566), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(G902), .B1(new_n592), .B2(new_n525), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n588), .A2(new_n589), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n594), .A2(KEYINPUT74), .A3(G472), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT74), .B1(new_n594), .B2(G472), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n575), .A2(new_n578), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT76), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(G472), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT74), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(KEYINPUT74), .A3(G472), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n576), .A2(new_n577), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n570), .A2(KEYINPUT32), .A3(new_n571), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(KEYINPUT75), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n576), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n574), .A3(KEYINPUT32), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT76), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n603), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n521), .B1(new_n598), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(KEYINPUT82), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT82), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n614), .B(new_n521), .C1(new_n598), .C2(new_n611), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n294), .B(new_n474), .C1(new_n613), .C2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G101), .ZN(G3));
  INV_X1    g431(.A(new_n521), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n293), .ZN(new_n619));
  INV_X1    g433(.A(new_n290), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n570), .A2(new_n281), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n607), .B1(G472), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT102), .Z(new_n625));
  AOI21_X1  g439(.A(new_n400), .B1(new_n344), .B2(new_n353), .ZN(new_n626));
  INV_X1    g440(.A(G478), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n393), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n388), .A2(KEYINPUT33), .A3(new_n390), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n391), .A2(new_n392), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n629), .B1(new_n633), .B2(KEYINPUT33), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n632), .B1(new_n634), .B2(KEYINPUT104), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(G478), .A3(new_n281), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n626), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n472), .A2(KEYINPUT103), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n406), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n471), .A2(KEYINPUT103), .A3(new_n472), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n637), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n625), .A2(new_n363), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND2_X1  g458(.A1(new_n343), .A2(KEYINPUT20), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n352), .A2(new_n295), .A3(new_n281), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n401), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n398), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n639), .A2(new_n649), .A3(new_n640), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n625), .A2(new_n363), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT105), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT35), .B(G107), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n505), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n501), .ZN(new_n657));
  INV_X1    g471(.A(new_n514), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n281), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n519), .A2(new_n655), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n516), .A3(new_n518), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT107), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n474), .A2(new_n294), .A3(new_n622), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT109), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT108), .B(KEYINPUT37), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  NAND2_X1  g484(.A1(new_n598), .A2(new_n611), .ZN(new_n671));
  INV_X1    g485(.A(G900), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n357), .B1(new_n361), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n639), .A2(new_n649), .A3(new_n640), .A4(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n671), .A2(new_n675), .A3(new_n294), .A4(new_n665), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  XNOR2_X1  g491(.A(new_n673), .B(KEYINPUT39), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n294), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT110), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n398), .B(new_n626), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n681), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n406), .B1(new_n684), .B2(KEYINPUT40), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n662), .A2(new_n664), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n471), .A2(new_n472), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT38), .Z(new_n688));
  INV_X1    g502(.A(G472), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n554), .B1(new_n525), .B2(new_n590), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n689), .B1(new_n690), .B2(new_n281), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n609), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n688), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n683), .A2(new_n685), .A3(new_n686), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  AND3_X1   g511(.A1(new_n639), .A2(new_n294), .A3(new_n640), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n637), .A2(new_n674), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n671), .A2(new_n665), .A3(new_n698), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G146), .ZN(G48));
  NOR2_X1   g515(.A1(new_n285), .A2(new_n286), .ZN(new_n702));
  OAI21_X1  g516(.A(G469), .B1(new_n702), .B2(G902), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n287), .ZN(new_n704));
  INV_X1    g518(.A(new_n293), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n704), .A2(new_n705), .A3(new_n362), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n612), .A2(new_n641), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT41), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G113), .ZN(G15));
  NAND4_X1  g523(.A1(new_n671), .A2(new_n618), .A3(new_n650), .A4(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NOR2_X1   g525(.A1(new_n704), .A2(new_n705), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n639), .A2(new_n640), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n671), .A2(new_n404), .A3(new_n665), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  OAI21_X1  g529(.A(new_n567), .B1(new_n590), .B2(new_n566), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n554), .A2(KEYINPUT31), .B1(new_n558), .B2(new_n716), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n717), .A2(KEYINPUT111), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(KEYINPUT111), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n557), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT112), .B(G472), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n720), .A2(new_n571), .B1(new_n621), .B2(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n618), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n626), .A2(new_n398), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n639), .A2(new_n724), .A3(new_n640), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n725), .A3(new_n706), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND4_X1  g541(.A1(new_n699), .A2(new_n713), .A3(new_n665), .A4(new_n722), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G125), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n290), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n279), .A2(new_n287), .A3(KEYINPUT113), .A4(new_n289), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n471), .A2(new_n293), .A3(new_n405), .A4(new_n472), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n603), .A2(new_n610), .A3(new_n609), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n610), .B1(new_n603), .B2(new_n609), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n618), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n699), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT114), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n612), .A2(new_n742), .A3(new_n699), .A4(new_n735), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n572), .B1(new_n601), .B2(new_n602), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n521), .B1(new_n745), .B2(new_n604), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n699), .A2(KEYINPUT42), .A3(new_n746), .A4(new_n735), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  NAND4_X1  g563(.A1(new_n612), .A2(new_n649), .A3(new_n674), .A4(new_n735), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  AND2_X1   g565(.A1(new_n276), .A2(new_n278), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(KEYINPUT45), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(G469), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n289), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT115), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(KEYINPUT46), .A3(new_n289), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n287), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n756), .A2(new_n762), .A3(new_n757), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n764), .A2(new_n705), .A3(new_n678), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n626), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n636), .A2(new_n628), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n626), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n767), .B(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n623), .A3(new_n665), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n406), .B(new_n687), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n765), .B(new_n773), .C1(new_n772), .C2(new_n771), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G137), .ZN(G39));
  INV_X1    g589(.A(KEYINPUT47), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n764), .B2(new_n705), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(KEYINPUT47), .A3(new_n293), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n687), .A2(new_n406), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n671), .A2(new_n618), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n699), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G140), .ZN(G42));
  INV_X1    g598(.A(new_n704), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n619), .A2(new_n787), .A3(new_n406), .A4(new_n769), .ZN(new_n788));
  XOR2_X1   g602(.A(new_n788), .B(KEYINPUT117), .Z(new_n789));
  AOI21_X1  g603(.A(new_n693), .B1(new_n786), .B2(new_n785), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(new_n688), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n705), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n777), .A2(new_n779), .A3(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n770), .A2(new_n357), .A3(new_n723), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n781), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n734), .A2(new_n356), .A3(new_n704), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n796), .A2(new_n618), .A3(new_n694), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n626), .A3(new_n628), .A4(new_n636), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT121), .Z(new_n799));
  NAND4_X1  g613(.A1(new_n794), .A2(new_n406), .A3(new_n688), .A4(new_n712), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n770), .A2(new_n796), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n665), .A2(new_n722), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n795), .A2(new_n799), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n803), .A2(new_n746), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT122), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT122), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(KEYINPUT48), .A3(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(G952), .A3(new_n272), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n808), .A2(new_n809), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n794), .A2(new_n713), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n733), .A2(new_n663), .A3(new_n673), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n725), .A2(new_n817), .A3(new_n293), .A4(new_n693), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n676), .A2(new_n700), .A3(new_n728), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(KEYINPUT119), .B(KEYINPUT52), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n804), .A2(new_n699), .A3(new_n735), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n686), .B1(new_n598), .B2(new_n611), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n398), .A2(new_n674), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n294), .A3(new_n781), .A4(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n750), .B(new_n822), .C1(new_n825), .C2(new_n648), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n748), .A2(new_n827), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n707), .A2(new_n714), .A3(new_n710), .A4(new_n726), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n626), .A2(new_n768), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n398), .B2(new_n626), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n624), .A2(new_n363), .A3(new_n473), .A4(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n616), .A3(new_n666), .A4(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n821), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n828), .A2(new_n833), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n819), .A2(KEYINPUT118), .A3(KEYINPUT52), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(new_n819), .B2(KEYINPUT118), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n837), .A2(new_n835), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n842), .ZN(new_n843));
  AND4_X1   g657(.A1(KEYINPUT53), .A2(new_n616), .A3(new_n666), .A4(new_n832), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n826), .B1(new_n744), .B2(new_n747), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n707), .A2(new_n714), .A3(new_n710), .A4(new_n726), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT120), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n841), .A2(new_n844), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n848), .B(new_n849), .C1(new_n834), .C2(KEYINPUT53), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n815), .A2(new_n816), .A3(new_n843), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n811), .A2(KEYINPUT48), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n797), .A2(new_n637), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(G952), .A2(G953), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT123), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n791), .B1(new_n854), .B2(new_n856), .ZN(G75));
  INV_X1    g671(.A(new_n821), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n837), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n616), .A2(new_n666), .A3(new_n832), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n819), .A2(KEYINPUT118), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n860), .A2(new_n863), .A3(KEYINPUT53), .A4(new_n838), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n846), .A2(KEYINPUT120), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n846), .A2(KEYINPUT120), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n748), .B(new_n827), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n281), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(G210), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n455), .A2(new_n438), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(new_n444), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n871), .B2(new_n872), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n272), .A2(G952), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT124), .Z(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n876), .A2(new_n877), .A3(new_n880), .ZN(G51));
  OAI21_X1  g695(.A(KEYINPUT54), .B1(new_n859), .B2(new_n868), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n882), .A2(new_n883), .A3(new_n850), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n869), .A2(KEYINPUT125), .A3(new_n849), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n288), .B(KEYINPUT57), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n702), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT126), .A4(new_n886), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n869), .A2(new_n281), .A3(new_n755), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n880), .B1(new_n892), .B2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n331), .B2(new_n342), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .A4(new_n338), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n880), .B1(new_n896), .B2(new_n897), .ZN(G60));
  NAND2_X1  g712(.A1(G478), .A2(G902), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT59), .Z(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n843), .B2(new_n850), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n879), .B1(new_n901), .B2(new_n635), .ZN(new_n902));
  INV_X1    g716(.A(new_n900), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n635), .A2(new_n884), .A3(new_n885), .A4(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n869), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n657), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n506), .A2(new_n508), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n909), .B(new_n879), .C1(new_n911), .C2(new_n908), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G66));
  AOI21_X1  g728(.A(new_n272), .B1(new_n358), .B2(new_n442), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n833), .B2(new_n272), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n873), .B1(G898), .B2(new_n272), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n916), .B(new_n917), .Z(G69));
  AND2_X1   g732(.A1(new_n783), .A2(new_n774), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n676), .A2(new_n700), .A3(new_n728), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n696), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT62), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n613), .A2(new_n615), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n924), .A2(new_n681), .A3(new_n781), .A4(new_n831), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n919), .A2(new_n922), .A3(new_n923), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n272), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n547), .B(new_n333), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n272), .A2(G900), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT127), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n765), .A2(new_n725), .A3(new_n746), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n933), .A2(new_n748), .A3(new_n920), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n919), .A2(new_n750), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n932), .B1(new_n935), .B2(new_n272), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(G72));
  NAND2_X1  g753(.A1(G472), .A2(G902), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT63), .Z(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n926), .B2(new_n833), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n584), .A3(new_n525), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n935), .B2(new_n833), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n551), .A3(new_n548), .A4(new_n558), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n554), .A2(new_n585), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n836), .A2(new_n842), .A3(new_n941), .A4(new_n946), .ZN(new_n947));
  AND4_X1   g761(.A1(new_n879), .A2(new_n943), .A3(new_n945), .A4(new_n947), .ZN(G57));
endmodule


