//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR3_X1   g0018(.A1(new_n217), .A2(new_n210), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT65), .B(G238), .Z(new_n221));
  XOR2_X1   g0021(.A(KEYINPUT66), .B(G244), .Z(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n212), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  NOR4_X1   g0031(.A1(new_n216), .A2(new_n219), .A3(new_n230), .A4(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G50), .B(G68), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XOR2_X1   g0042(.A(G58), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  OR2_X1    g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(new_n210), .A3(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT7), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n250), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n220), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G58), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n220), .ZN(new_n257));
  OAI21_X1  g0057(.A(G20), .B1(new_n257), .B2(new_n201), .ZN(new_n258));
  INV_X1    g0058(.A(G159), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT76), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT16), .ZN(new_n264));
  NAND3_X1  g0064(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(new_n218), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT16), .ZN(new_n267));
  OAI211_X1 g0067(.A(KEYINPUT76), .B(new_n267), .C1(new_n255), .C2(new_n262), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  OAI211_X1 g0072(.A(G223), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(G226), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G87), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(new_n218), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT77), .ZN(new_n280));
  INV_X1    g0080(.A(G190), .ZN(new_n281));
  OAI21_X1  g0081(.A(G274), .B1(new_n277), .B2(new_n218), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT68), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  AND2_X1   g0085(.A1(G1), .A2(G13), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  INV_X1    g0089(.A(new_n283), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n287), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n283), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n284), .A2(new_n291), .B1(new_n294), .B2(G232), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT77), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n276), .A2(new_n296), .A3(new_n278), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n280), .A2(new_n281), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n284), .A2(new_n291), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n294), .A2(G232), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n276), .A2(new_n278), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n256), .A2(KEYINPUT8), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT8), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G58), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n209), .A2(G20), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n314), .A2(new_n266), .ZN(new_n315));
  INV_X1    g0115(.A(new_n309), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n312), .A2(new_n315), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n269), .A2(new_n305), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT17), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n269), .A2(new_n317), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT18), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n280), .A2(new_n323), .A3(new_n295), .A4(new_n297), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n302), .B2(new_n303), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n321), .A2(new_n322), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n317), .ZN(new_n330));
  INV_X1    g0130(.A(new_n266), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n263), .B2(KEYINPUT16), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n332), .B2(new_n268), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT18), .B1(new_n333), .B2(new_n327), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(KEYINPUT17), .A3(new_n305), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n320), .A2(new_n329), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n314), .A2(new_n220), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT12), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n210), .A2(G33), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n223), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT11), .A3(new_n266), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n315), .A2(G68), .A3(new_n310), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT11), .B1(new_n342), .B2(new_n266), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  AND3_X1   g0150(.A1(new_n284), .A2(new_n350), .A3(new_n291), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n284), .B2(new_n291), .ZN(new_n352));
  INV_X1    g0152(.A(G238), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(new_n293), .ZN(new_n354));
  OAI211_X1 g0154(.A(G232), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n355));
  OAI211_X1 g0155(.A(G226), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G33), .A2(G97), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT74), .A4(new_n357), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n292), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n354), .A2(KEYINPUT13), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  NOR3_X1   g0164(.A1(new_n282), .A2(KEYINPUT68), .A3(new_n283), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT75), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n284), .A2(new_n350), .A3(new_n291), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n367), .A2(new_n368), .B1(G238), .B2(new_n294), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n360), .A2(new_n361), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n278), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n364), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n349), .B(G169), .C1(new_n363), .C2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT13), .B1(new_n354), .B2(new_n362), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n371), .A3(new_n364), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(G179), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n349), .B1(new_n378), .B2(G169), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n348), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(G200), .B1(new_n363), .B2(new_n372), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n374), .A2(new_n375), .A3(G190), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n347), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n337), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n249), .A2(new_n250), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(G222), .A3(new_n270), .ZN(new_n386));
  INV_X1    g0186(.A(G223), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(G1698), .ZN(new_n388));
  OAI221_X1 g0188(.A(new_n386), .B1(new_n223), .B2(new_n385), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT69), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n292), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n390), .B2(new_n389), .ZN(new_n392));
  INV_X1    g0192(.A(new_n300), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(G226), .B2(new_n294), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G190), .ZN(new_n397));
  INV_X1    g0197(.A(new_n341), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n309), .A2(new_n398), .B1(G150), .B2(new_n260), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(KEYINPUT70), .B1(G20), .B2(new_n203), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(KEYINPUT70), .B2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n266), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n315), .A2(new_n403), .B1(new_n202), .B2(new_n314), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT9), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n395), .A2(G200), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n397), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT10), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT10), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n397), .A2(new_n406), .A3(new_n410), .A4(new_n407), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n396), .A2(new_n323), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n405), .B1(new_n396), .B2(G169), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XOR2_X1   g0216(.A(KEYINPUT15), .B(G87), .Z(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n341), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n316), .A2(new_n261), .B1(new_n210), .B2(new_n223), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n266), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n223), .B1(new_n209), .B2(G20), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n315), .A2(new_n422), .B1(new_n223), .B2(new_n314), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n385), .A2(G232), .A3(new_n270), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n426), .B1(new_n206), .B2(new_n385), .C1(new_n388), .C2(new_n221), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(KEYINPUT71), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n292), .B1(new_n427), .B2(KEYINPUT71), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n300), .B1(new_n222), .B2(new_n293), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n425), .B1(new_n433), .B2(new_n325), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n431), .B1(new_n428), .B2(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n323), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n424), .A2(KEYINPUT72), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n424), .A2(KEYINPUT72), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n439), .B(new_n440), .C1(new_n435), .C2(new_n299), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n433), .A2(new_n281), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n412), .A2(new_n416), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT73), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT73), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n412), .A2(new_n447), .A3(new_n416), .A4(new_n444), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n384), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n417), .A2(new_n313), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT19), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n210), .B1(new_n357), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n452), .B1(G87), .B2(new_n207), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n210), .B(G68), .C1(new_n271), .C2(new_n272), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n451), .B1(new_n341), .B2(new_n205), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n331), .B1(new_n456), .B2(KEYINPUT83), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT83), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n453), .A2(new_n458), .A3(new_n454), .A4(new_n455), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n450), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n209), .A2(G33), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n313), .A2(new_n461), .A3(new_n218), .A4(new_n265), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n417), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n209), .A2(G45), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G250), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT82), .B1(new_n278), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n288), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n292), .A2(new_n471), .A3(G250), .A4(new_n465), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n353), .A2(new_n270), .ZN(new_n474));
  INV_X1    g0274(.A(G244), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G1698), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n476), .C1(new_n271), .C2(new_n272), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n292), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n460), .A2(new_n464), .B1(new_n323), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n325), .B1(new_n473), .B2(new_n479), .ZN(new_n482));
  INV_X1    g0282(.A(G87), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n462), .A2(new_n483), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n450), .B(new_n484), .C1(new_n457), .C2(new_n459), .ZN(new_n485));
  AND3_X1   g0285(.A1(new_n467), .A2(new_n470), .A3(new_n472), .ZN(new_n486));
  INV_X1    g0286(.A(new_n479), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n486), .A2(G190), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(G200), .B1(new_n473), .B2(new_n479), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n481), .A2(new_n482), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  OR3_X1    g0291(.A1(new_n478), .A2(KEYINPUT87), .A3(G20), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT23), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n210), .B2(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT87), .B1(new_n478), .B2(G20), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n492), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n210), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT24), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n498), .B(new_n504), .C1(new_n500), .C2(new_n501), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n331), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n314), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT25), .B1(new_n314), .B2(new_n206), .ZN(new_n508));
  OAI22_X1  g0308(.A1(new_n507), .A2(new_n508), .B1(new_n206), .B2(new_n462), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n469), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND3_X1   g0313(.A1(new_n513), .A2(G264), .A3(new_n292), .ZN(new_n514));
  OAI211_X1 g0314(.A(G257), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT88), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n385), .A2(KEYINPUT88), .A3(G257), .A4(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G294), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n385), .A2(G250), .A3(new_n270), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n514), .B1(new_n521), .B2(new_n278), .ZN(new_n522));
  XNOR2_X1  g0322(.A(KEYINPUT5), .B(G41), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n288), .A2(new_n469), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(new_n281), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n524), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n526), .B(new_n514), .C1(new_n521), .C2(new_n278), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n525), .B1(new_n527), .B2(G200), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n510), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n522), .A2(new_n524), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n325), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n323), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(new_n506), .C2(new_n509), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n491), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n513), .A2(new_n292), .ZN(new_n535));
  INV_X1    g0335(.A(G257), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n524), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT80), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n524), .B(KEYINPUT80), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(G250), .A2(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(KEYINPUT4), .A2(G244), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(G1698), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n385), .A2(new_n544), .B1(G33), .B2(G283), .ZN(new_n545));
  OAI211_X1 g0345(.A(G244), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT4), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT79), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n545), .A2(new_n548), .A3(KEYINPUT79), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n278), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n541), .A2(new_n553), .A3(G179), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n292), .B1(new_n549), .B2(new_n550), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n552), .A2(new_n555), .B1(new_n539), .B2(new_n540), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n556), .B2(new_n325), .ZN(new_n557));
  XNOR2_X1  g0357(.A(G97), .B(G107), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT6), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n559), .A2(new_n205), .A3(G107), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n563), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n253), .A2(new_n254), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G107), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n331), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n313), .A2(G97), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n463), .B2(G97), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(KEYINPUT81), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n561), .B1(new_n559), .B2(new_n558), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n572), .A2(new_n210), .B1(new_n223), .B2(new_n261), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n206), .B1(new_n253), .B2(new_n254), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n266), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT81), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n569), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n557), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT78), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n575), .B2(new_n569), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n575), .A2(new_n580), .A3(new_n569), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n541), .A2(new_n553), .A3(new_n281), .ZN(new_n584));
  AOI21_X1  g0384(.A(G200), .B1(new_n541), .B2(new_n553), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n271), .A2(new_n272), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n292), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  MUX2_X1   g0390(.A(G257), .B(G264), .S(G1698), .Z(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n513), .A2(G270), .A3(new_n292), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n593), .A2(new_n524), .A3(KEYINPUT84), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT84), .B1(new_n593), .B2(new_n524), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(G33), .A2(G283), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n597), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n598));
  INV_X1    g0398(.A(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G20), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n266), .A3(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n598), .A2(KEYINPUT20), .A3(new_n266), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n313), .A2(G116), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n463), .B2(G116), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n325), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n596), .A2(KEYINPUT21), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n593), .A2(new_n524), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT84), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n593), .A2(new_n524), .A3(KEYINPUT84), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n323), .B1(new_n605), .B2(new_n607), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n592), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n596), .A2(G200), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n605), .A2(new_n607), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(new_n281), .C2(new_n596), .ZN(new_n620));
  XNOR2_X1  g0420(.A(KEYINPUT85), .B(KEYINPUT21), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n596), .B2(new_n608), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n622), .A2(KEYINPUT86), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT86), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n624), .B(new_n621), .C1(new_n596), .C2(new_n608), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n617), .B(new_n620), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n534), .A2(new_n587), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n449), .A2(new_n627), .ZN(G372));
  OAI211_X1 g0428(.A(new_n533), .B(new_n617), .C1(new_n623), .C2(new_n625), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n556), .A2(new_n281), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(G200), .B2(new_n556), .ZN(new_n631));
  INV_X1    g0431(.A(new_n583), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n632), .A2(new_n581), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n631), .A2(new_n633), .B1(new_n557), .B2(new_n578), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n479), .A2(KEYINPUT89), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT89), .ZN(new_n636));
  AOI211_X1 g0436(.A(new_n636), .B(new_n292), .C1(new_n477), .C2(new_n478), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n486), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G200), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(new_n488), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n510), .A2(new_n528), .B1(new_n640), .B2(new_n485), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n629), .A2(new_n634), .A3(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  INV_X1    g0443(.A(new_n554), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n325), .B1(new_n541), .B2(new_n553), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n644), .A2(new_n645), .B1(new_n632), .B2(new_n581), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n485), .A2(new_n488), .A3(new_n639), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n638), .A2(new_n325), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n649), .A2(new_n266), .A3(new_n459), .ZN(new_n650));
  INV_X1    g0450(.A(new_n450), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n464), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n480), .A2(new_n323), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n643), .B1(new_n646), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n541), .A2(new_n553), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G169), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n658), .A2(new_n554), .B1(new_n571), .B2(new_n577), .ZN(new_n659));
  XOR2_X1   g0459(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n491), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n642), .A2(new_n662), .A3(new_n654), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n449), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n416), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n329), .A2(new_n334), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(G169), .B1(new_n363), .B2(new_n372), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT14), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n376), .A3(new_n373), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n348), .A2(new_n670), .B1(new_n438), .B2(new_n383), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n320), .A2(new_n335), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n667), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n665), .B1(new_n673), .B2(new_n412), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n664), .A2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n506), .B2(new_n509), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n529), .A2(new_n533), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n531), .A2(new_n532), .ZN(new_n684));
  OAI211_X1 g0484(.A(new_n683), .B(KEYINPUT91), .C1(new_n684), .C2(new_n682), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n684), .A2(new_n682), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT91), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n686), .B1(new_n685), .B2(new_n689), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n617), .B1(new_n623), .B2(new_n625), .ZN(new_n694));
  INV_X1    g0494(.A(new_n681), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n533), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n697), .B1(new_n698), .B2(new_n695), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n619), .A2(new_n695), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n626), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n693), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n213), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n217), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  AOI21_X1  g0513(.A(KEYINPUT29), .B1(new_n663), .B2(new_n695), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n642), .A2(new_n654), .ZN(new_n716));
  OR3_X1    g0516(.A1(new_n646), .A2(new_n655), .A3(new_n643), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n659), .A2(new_n491), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n717), .B1(new_n718), .B2(new_n660), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n681), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n715), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n592), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n614), .A2(new_n522), .A3(new_n480), .A4(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n725), .B1(new_n727), .B2(new_n657), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n486), .A2(new_n592), .A3(new_n487), .A4(G179), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n594), .A2(new_n595), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(new_n556), .A3(KEYINPUT30), .A4(new_n522), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G238), .A2(G1698), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n475), .B2(G1698), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n734), .A2(new_n385), .B1(G33), .B2(G116), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n636), .B1(new_n735), .B2(new_n292), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n479), .A2(KEYINPUT89), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(G179), .B1(new_n738), .B2(new_n486), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n657), .A2(new_n739), .A3(new_n596), .A4(new_n530), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n728), .A2(new_n732), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(KEYINPUT31), .B1(new_n741), .B2(new_n681), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n724), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n744), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(KEYINPUT93), .A3(new_n742), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n491), .A2(new_n529), .A3(new_n533), .ZN(new_n748));
  INV_X1    g0548(.A(new_n626), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n748), .A2(new_n749), .A3(new_n634), .A4(new_n695), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n745), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n723), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n713), .B1(new_n754), .B2(G1), .ZN(G364));
  INV_X1    g0555(.A(new_n703), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n210), .A2(G13), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n209), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n708), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G330), .B2(new_n702), .ZN(new_n762));
  NOR2_X1   g0562(.A1(G13), .A2(G33), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n218), .B1(G20), .B2(new_n325), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n244), .A2(G45), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n707), .A2(new_n385), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(G45), .C2(new_n217), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n707), .A2(new_n588), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n772), .A2(G355), .B1(new_n599), .B2(new_n707), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n768), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n766), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n210), .A2(new_n323), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(G200), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n281), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G326), .ZN(new_n780));
  INV_X1    g0580(.A(G294), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n281), .A2(G179), .A3(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n210), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n210), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT95), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n786), .A2(new_n787), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n784), .A2(KEYINPUT96), .B1(new_n791), .B2(G303), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n776), .A2(G190), .A3(new_n299), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n785), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n794), .A2(G322), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n776), .A2(new_n795), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n588), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n777), .A2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n785), .A2(new_n281), .A3(G200), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n792), .B(new_n808), .C1(KEYINPUT96), .C2(new_n784), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n803), .A2(new_n220), .B1(new_n779), .B2(new_n202), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n783), .A2(new_n205), .B1(new_n806), .B2(new_n206), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n791), .A2(G87), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n796), .A2(new_n259), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT32), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n385), .B1(new_n793), .B2(new_n256), .ZN(new_n816));
  INV_X1    g0616(.A(new_n800), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(G77), .B2(new_n817), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n775), .B1(new_n809), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n760), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n774), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n765), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n702), .B2(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n762), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G396));
  AOI22_X1  g0626(.A1(new_n794), .A2(G143), .B1(new_n817), .B2(G159), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n827), .B1(new_n779), .B2(new_n828), .C1(new_n829), .C2(new_n803), .ZN(new_n830));
  XOR2_X1   g0630(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT98), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n830), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n791), .A2(G50), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n385), .B1(new_n796), .B2(new_n836), .C1(new_n783), .C2(new_n256), .ZN(new_n837));
  INV_X1    g0637(.A(new_n806), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n837), .B1(G68), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n790), .A2(new_n206), .ZN(new_n841));
  INV_X1    g0641(.A(new_n783), .ZN(new_n842));
  AOI22_X1  g0642(.A1(G97), .A2(new_n842), .B1(new_n778), .B2(G303), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n806), .A2(new_n483), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G283), .B2(new_n802), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n385), .B1(new_n797), .B2(G311), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n794), .A2(G294), .B1(new_n817), .B2(G116), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n843), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n840), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n775), .B1(new_n849), .B2(KEYINPUT99), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(KEYINPUT99), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n766), .A2(new_n763), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n821), .B1(new_n223), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n434), .A2(new_n436), .A3(new_n695), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n441), .A2(new_n442), .B1(new_n425), .B2(new_n695), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n437), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n851), .B(new_n853), .C1(new_n856), .C2(new_n764), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n663), .A2(new_n695), .A3(new_n856), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT100), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n663), .B2(new_n695), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n859), .B(new_n860), .Z(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n821), .B1(new_n862), .B2(new_n753), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n861), .A2(new_n752), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n857), .B1(new_n863), .B2(new_n864), .ZN(G384));
  INV_X1    g0665(.A(new_n679), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n667), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n854), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n858), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT101), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n383), .A2(new_n669), .A3(new_n376), .A4(new_n373), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n347), .A2(new_n695), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n872), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n380), .A2(new_n383), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n380), .A2(new_n870), .A3(new_n383), .A4(new_n874), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n869), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n318), .B1(new_n333), .B2(new_n327), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n333), .A2(new_n679), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n321), .A2(new_n328), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n321), .A2(new_n866), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .A4(new_n318), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n336), .A2(new_n882), .ZN(new_n889));
  AND3_X1   g0689(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n880), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n889), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n895), .A2(KEYINPUT102), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n867), .B1(new_n879), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n895), .A2(KEYINPUT104), .A3(new_n896), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n893), .A2(KEYINPUT104), .A3(new_n894), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n896), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n670), .A2(new_n348), .A3(new_n695), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT103), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT105), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT105), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n899), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n449), .A2(new_n722), .A3(new_n715), .A4(new_n721), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(new_n674), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n913), .B(new_n915), .Z(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n892), .A2(new_n897), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n741), .A2(new_n681), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT106), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT31), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n741), .A2(KEYINPUT106), .A3(new_n681), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT107), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n743), .B1(new_n627), .B2(new_n695), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(KEYINPUT107), .A3(new_n922), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n928), .A2(new_n856), .A3(new_n876), .A4(new_n877), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n917), .B1(new_n918), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT108), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND3_X1   g0732(.A1(new_n921), .A2(KEYINPUT107), .A3(new_n922), .ZN(new_n933));
  AOI21_X1  g0733(.A(KEYINPUT107), .B1(new_n921), .B2(new_n922), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n750), .A2(new_n742), .ZN(new_n935));
  NOR3_X1   g0735(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n876), .A2(new_n856), .A3(new_n877), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n898), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n939), .A2(KEYINPUT108), .A3(new_n917), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT40), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n932), .A2(new_n940), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n449), .A2(new_n928), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(G330), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n943), .A2(new_n944), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n916), .A2(new_n949), .B1(new_n209), .B2(new_n757), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n949), .B2(new_n916), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n563), .A2(KEYINPUT35), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n563), .A2(KEYINPUT35), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n218), .A2(new_n210), .A3(new_n599), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT36), .Z(new_n956));
  OR3_X1    g0756(.A1(new_n257), .A2(new_n217), .A3(new_n223), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n202), .A2(G68), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n209), .B(G13), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n951), .A2(new_n956), .A3(new_n959), .ZN(G367));
  INV_X1    g0760(.A(KEYINPUT42), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n634), .B1(new_n633), .B2(new_n695), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n646), .A2(new_n695), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n697), .A2(new_n961), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT109), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n698), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n681), .B1(new_n967), .B2(new_n579), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n697), .A2(new_n964), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(new_n969), .B2(KEYINPUT42), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n485), .A2(new_n695), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n655), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(new_n481), .A3(new_n648), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI22_X1  g0774(.A1(new_n966), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(KEYINPUT43), .B2(new_n974), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT43), .ZN(new_n977));
  INV_X1    g0777(.A(new_n974), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n966), .A2(new_n977), .A3(new_n978), .A4(new_n970), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n704), .A2(new_n964), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n983), .B2(new_n982), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n980), .A2(KEYINPUT110), .A3(new_n981), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n708), .B(KEYINPUT41), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n756), .B1(new_n697), .B2(KEYINPUT111), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n697), .A2(KEYINPUT111), .A3(new_n756), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n693), .A2(new_n696), .ZN(new_n992));
  NOR3_X1   g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n992), .ZN(new_n994));
  INV_X1    g0794(.A(new_n991), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(new_n995), .B2(new_n989), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(KEYINPUT112), .A3(new_n754), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n699), .A2(new_n964), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT45), .B1(new_n699), .B2(new_n964), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n697), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n533), .B2(new_n681), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n964), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT44), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n699), .A2(new_n1008), .A3(new_n964), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1003), .A2(new_n1010), .A3(new_n705), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT112), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n993), .A2(new_n996), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n754), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n1001), .A2(new_n1002), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n704), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n998), .A2(new_n1011), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n988), .B1(new_n1018), .B2(new_n754), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n986), .B(new_n987), .C1(new_n1019), .C2(new_n759), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n770), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n767), .B1(new_n213), .B2(new_n418), .C1(new_n1021), .C2(new_n239), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1022), .A2(new_n760), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n800), .A2(new_n202), .B1(new_n796), .B2(new_n828), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n588), .B(new_n1024), .C1(G150), .C2(new_n794), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n791), .A2(G58), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G143), .A2(new_n778), .B1(new_n802), .B2(G159), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n783), .A2(new_n220), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G77), .B2(new_n838), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G107), .A2(new_n842), .B1(new_n802), .B2(G294), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n793), .A2(new_n589), .B1(new_n800), .B2(new_n805), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n385), .B(new_n1032), .C1(G317), .C2(new_n797), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT46), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n790), .B2(new_n599), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n778), .A2(G311), .B1(new_n838), .B2(G97), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1033), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n790), .A2(new_n1034), .A3(new_n599), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1030), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT47), .Z(new_n1040));
  OAI221_X1 g0840(.A(new_n1023), .B1(new_n974), .B2(new_n823), .C1(new_n775), .C2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1020), .A2(new_n1041), .ZN(G387));
  INV_X1    g0842(.A(new_n998), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1015), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n708), .B1(new_n754), .B2(new_n997), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n693), .A2(new_n765), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n710), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n772), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(G107), .B2(new_n213), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n236), .A2(new_n468), .ZN(new_n1050));
  AOI211_X1 g0850(.A(G45), .B(new_n1047), .C1(G68), .C2(G77), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n309), .A2(new_n202), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT50), .Z(new_n1053));
  AOI21_X1  g0853(.A(new_n1021), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1049), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n760), .B1(new_n1055), .B2(new_n768), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n793), .A2(new_n202), .B1(new_n796), .B2(new_n829), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n588), .B(new_n1057), .C1(G68), .C2(new_n817), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n791), .A2(G77), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n842), .A2(new_n417), .B1(new_n838), .B2(G97), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(G159), .A2(new_n778), .B1(new_n802), .B2(new_n309), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(G317), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n793), .A2(new_n1063), .B1(new_n800), .B2(new_n589), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT113), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(KEYINPUT113), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G311), .A2(new_n802), .B1(new_n778), .B2(G322), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT48), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n790), .A2(new_n781), .B1(new_n805), .B2(new_n783), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1070), .A2(KEYINPUT49), .A3(new_n1072), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n588), .B1(new_n796), .B2(new_n780), .C1(new_n599), .C2(new_n806), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT114), .Z(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT49), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1062), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1056), .B1(new_n1078), .B2(new_n766), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n997), .A2(new_n759), .B1(new_n1046), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1045), .A2(new_n1080), .ZN(G393));
  INV_X1    g0881(.A(new_n1017), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1016), .A2(new_n704), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1082), .A2(new_n1083), .A3(new_n758), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1006), .A2(new_n765), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n767), .B1(new_n205), .B2(new_n213), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n770), .B2(new_n247), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n385), .B1(new_n797), .B2(G322), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n206), .B2(new_n806), .C1(new_n790), .C2(new_n805), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT115), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n779), .A2(new_n1063), .B1(new_n799), .B2(new_n793), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n802), .A2(G303), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n842), .A2(G116), .B1(new_n817), .B2(G294), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G150), .A2(new_n778), .B1(new_n794), .B2(G159), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n783), .A2(new_n223), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n844), .B(new_n1098), .C1(G50), .C2(new_n802), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n791), .A2(G68), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n797), .A2(G143), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n588), .B1(new_n817), .B2(new_n309), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1090), .A2(new_n1095), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n821), .B(new_n1087), .C1(new_n1104), .C2(new_n766), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1084), .B1(new_n1085), .B2(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1043), .A2(new_n1044), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n1018), .A3(new_n708), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(G390));
  NAND2_X1  g0909(.A1(new_n858), .A2(new_n868), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1110), .A2(new_n876), .A3(new_n877), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n903), .A2(new_n904), .B1(new_n1111), .B2(new_n906), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n900), .A2(new_n901), .A3(new_n906), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT116), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n876), .A2(new_n1114), .A3(new_n877), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n876), .B2(new_n877), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n855), .A2(new_n437), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n720), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n868), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1113), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n937), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n928), .A2(G330), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n753), .C1(new_n1123), .C2(KEYINPUT117), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1112), .A2(new_n1121), .A3(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n934), .A2(new_n935), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n947), .B1(new_n1126), .B2(new_n927), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n1127), .A2(new_n1122), .A3(KEYINPUT117), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n900), .A2(new_n901), .A3(new_n906), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1116), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n876), .A2(new_n1114), .A3(new_n877), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n854), .B1(new_n720), .B2(new_n1118), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1129), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n903), .A2(new_n904), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1111), .A2(new_n906), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1128), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1125), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n449), .A2(new_n1127), .ZN(new_n1140));
  AND3_X1   g0940(.A1(new_n914), .A2(new_n674), .A3(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n751), .A2(G330), .A3(new_n856), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(new_n878), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1143), .A2(KEYINPUT118), .B1(new_n1127), .B2(new_n1122), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT118), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1142), .A2(new_n1145), .A3(new_n878), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n869), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1133), .B1(new_n752), .B2(new_n937), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1127), .A2(new_n856), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n1132), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1141), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n709), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n793), .A2(new_n599), .B1(new_n800), .B2(new_n205), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n385), .B(new_n1154), .C1(G294), .C2(new_n797), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1098), .B1(G68), .B2(new_n838), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G107), .A2(new_n802), .B1(new_n778), .B2(G283), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1155), .A2(new_n813), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G159), .A2(new_n842), .B1(new_n802), .B2(G137), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n793), .A2(new_n836), .B1(new_n800), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n588), .B(new_n1161), .C1(G125), .C2(new_n797), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT53), .B1(new_n790), .B2(new_n829), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n778), .A2(G128), .B1(new_n838), .B2(G50), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1159), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n790), .A2(KEYINPUT53), .A3(new_n829), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1158), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n766), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n852), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n760), .C1(new_n309), .C2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1135), .B2(new_n763), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1139), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n759), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1153), .A2(new_n1173), .ZN(G378));
  OAI21_X1  g0974(.A(G330), .B1(new_n929), .B2(new_n941), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT119), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n405), .A2(new_n866), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n412), .A2(new_n416), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1178), .B1(new_n412), .B2(new_n416), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n412), .A2(new_n416), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1178), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1182), .B1(new_n1187), .B2(new_n1179), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1177), .B1(new_n1184), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1183), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1187), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1190), .A2(new_n1191), .A3(KEYINPUT119), .A4(KEYINPUT120), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT108), .B1(new_n939), .B2(new_n917), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n931), .B(KEYINPUT40), .C1(new_n938), .C2(new_n898), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1176), .B(new_n1193), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1175), .B1(new_n932), .B2(new_n940), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1190), .A2(KEYINPUT120), .A3(new_n1191), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1196), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n913), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n913), .B(new_n1196), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n759), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1189), .ZN(new_n1204));
  NOR3_X1   g1004(.A1(new_n1184), .A2(new_n1188), .A3(new_n1177), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n763), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n760), .B1(G50), .B2(new_n1169), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1208));
  INV_X1    g1008(.A(G41), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1208), .B1(new_n588), .B2(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n418), .A2(new_n800), .B1(new_n206), .B2(new_n793), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n588), .B(new_n1209), .C1(new_n796), .C2(new_n805), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1028), .B1(G58), .B2(new_n838), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G97), .A2(new_n802), .B1(new_n778), .B2(G116), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1059), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT58), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1210), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G128), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n793), .A2(new_n1219), .B1(new_n800), .B2(new_n828), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G132), .B2(new_n802), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G150), .A2(new_n842), .B1(new_n778), .B2(G125), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n790), .C2(new_n1160), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n838), .A2(G159), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1218), .B1(new_n1217), .B2(new_n1216), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1207), .B1(new_n1229), .B2(new_n766), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1206), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1203), .A2(KEYINPUT121), .A3(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT121), .B1(new_n1203), .B2(new_n1231), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1141), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1201), .A2(new_n1235), .A3(new_n1202), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT57), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1201), .A2(new_n1235), .A3(new_n1202), .A4(KEYINPUT57), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n708), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1234), .A2(new_n1240), .ZN(G375));
  AOI21_X1  g1041(.A(new_n821), .B1(new_n220), .B2(new_n852), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n794), .A2(G283), .B1(new_n797), .B2(G303), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1243), .B(new_n588), .C1(new_n206), .C2(new_n800), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n842), .A2(new_n417), .B1(new_n838), .B2(G77), .ZN(new_n1245));
  OAI221_X1 g1045(.A(new_n1245), .B1(new_n599), .B2(new_n803), .C1(new_n781), .C2(new_n779), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1244), .B(new_n1246), .C1(G97), .C2(new_n791), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n783), .A2(new_n202), .B1(new_n800), .B2(new_n829), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT123), .Z(new_n1249));
  NAND2_X1  g1049(.A1(new_n778), .A2(G132), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n828), .B2(new_n793), .C1(new_n803), .C2(new_n1160), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n385), .B1(new_n256), .B2(new_n806), .C1(new_n1251), .C2(KEYINPUT122), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1249), .B(new_n1252), .C1(KEYINPUT122), .C2(new_n1251), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n790), .A2(new_n259), .B1(new_n1219), .B2(new_n796), .ZN(new_n1254));
  XOR2_X1   g1054(.A(new_n1254), .B(KEYINPUT124), .Z(new_n1255));
  AOI21_X1  g1055(.A(new_n1247), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n1242), .B1(new_n775), .B2(new_n1256), .C1(new_n1117), .C2(new_n764), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n758), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1151), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1260), .A2(new_n988), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1141), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1259), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(G381));
  INV_X1    g1065(.A(G390), .ZN(new_n1266));
  INV_X1    g1066(.A(G384), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1045), .A2(new_n825), .A3(new_n1080), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1264), .A4(new_n1268), .ZN(new_n1269));
  OR4_X1    g1069(.A1(G387), .A2(new_n1269), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1070(.A(G378), .ZN(new_n1271));
  INV_X1    g1071(.A(G213), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(G343), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(G375), .C2(new_n1274), .ZN(G409));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1259), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1151), .A2(KEYINPUT60), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1278), .A2(new_n1263), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1258), .A2(KEYINPUT60), .A3(new_n1262), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n708), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1277), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1267), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1273), .A2(G2897), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1283), .B(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1240), .B(G378), .C1(new_n1233), .C2(new_n1232), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1203), .B(new_n1231), .C1(new_n1236), .C2(new_n988), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1271), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1273), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1276), .B1(new_n1285), .B2(new_n1289), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1273), .B(new_n1283), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(KEYINPUT63), .B2(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1291), .A2(KEYINPUT63), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n825), .B1(new_n1045), .B2(new_n1080), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1268), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G387), .A2(new_n1266), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G390), .A2(new_n1020), .A3(new_n1041), .ZN(new_n1298));
  AND4_X1   g1098(.A1(KEYINPUT125), .A2(new_n1296), .A3(new_n1297), .A4(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT125), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1297), .A2(new_n1300), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1301), .A2(new_n1296), .B1(new_n1298), .B2(new_n1297), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1292), .B(new_n1293), .C1(new_n1299), .C2(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1299), .ZN(new_n1304));
  OAI21_X1  g1104(.A(KEYINPUT62), .B1(new_n1291), .B2(KEYINPUT126), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1283), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1273), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT126), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1290), .B1(new_n1305), .B2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1304), .B1(new_n1313), .B2(KEYINPUT127), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT127), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n1315), .B(new_n1290), .C1(new_n1305), .C2(new_n1312), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1303), .B1(new_n1314), .B2(new_n1316), .ZN(G405));
  AOI21_X1  g1117(.A(G378), .B1(new_n1234), .B2(new_n1240), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1286), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(new_n1283), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(new_n1304), .B(new_n1321), .ZN(G402));
endmodule


