//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n207), .A2(KEYINPUT75), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(KEYINPUT75), .ZN(new_n209));
  INV_X1    g008(.A(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT76), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n217), .B1(new_n207), .B2(KEYINPUT2), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n207), .A2(new_n217), .A3(KEYINPUT2), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n215), .B1(KEYINPUT2), .B2(new_n207), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n212), .A2(new_n207), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n214), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n225));
  INV_X1    g024(.A(G113gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G120gat), .ZN(new_n227));
  INV_X1    g026(.A(G120gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G113gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231));
  INV_X1    g030(.A(G127gat), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n231), .A2(new_n232), .A3(G134gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n234), .A2(new_n225), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(new_n226), .B2(G120gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT70), .B1(new_n228), .B2(G113gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(new_n226), .A3(G120gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n228), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n238), .A2(new_n239), .A3(new_n241), .A4(new_n242), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n230), .A2(new_n235), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n236), .A2(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n234), .A2(new_n231), .ZN(new_n247));
  INV_X1    g046(.A(new_n233), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n230), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n251), .A3(new_n223), .ZN(new_n252));
  INV_X1    g051(.A(new_n220), .ZN(new_n253));
  NOR3_X1   g052(.A1(new_n253), .A2(new_n215), .A3(new_n218), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n254), .B2(new_n213), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n245), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT78), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n261));
  AOI211_X1 g060(.A(new_n261), .B(new_n258), .C1(new_n245), .C2(new_n256), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT5), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT4), .B1(new_n250), .B2(new_n255), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n224), .A2(new_n244), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n259), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n224), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n255), .A2(KEYINPUT3), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n270), .A3(new_n250), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n267), .A2(KEYINPUT77), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT77), .B1(new_n267), .B2(new_n271), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n263), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n245), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(new_n266), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n275), .B(new_n271), .C1(new_n276), .C2(KEYINPUT79), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n277), .A2(KEYINPUT5), .A3(new_n259), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n206), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n280));
  INV_X1    g079(.A(new_n260), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n257), .A2(KEYINPUT78), .A3(new_n259), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n271), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n267), .A2(KEYINPUT77), .A3(new_n271), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n283), .A2(new_n286), .A3(KEYINPUT5), .A4(new_n287), .ZN(new_n288));
  OR3_X1    g087(.A1(new_n277), .A2(KEYINPUT5), .A3(new_n259), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n205), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n279), .A2(new_n280), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT80), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n289), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT6), .B1(new_n293), .B2(new_n206), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n295), .A3(new_n290), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n205), .B1(new_n288), .B2(new_n289), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT65), .ZN(new_n301));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT26), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(new_n302), .B2(new_n303), .ZN(new_n306));
  OAI211_X1 g105(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n301), .A2(new_n304), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT27), .B(G183gat), .ZN(new_n310));
  INV_X1    g109(.A(G190gat), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n310), .A2(KEYINPUT28), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT28), .B1(new_n310), .B2(new_n311), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n308), .B(new_n309), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n302), .B(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n309), .ZN(new_n318));
  NAND4_X1  g117(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n316), .A2(new_n323), .A3(new_n301), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n318), .A2(new_n320), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n316), .A2(new_n326), .A3(new_n301), .A4(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n314), .A2(new_n325), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n244), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n316), .A2(new_n327), .A3(new_n301), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n331), .A2(new_n326), .B1(new_n324), .B2(KEYINPUT25), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n250), .A3(new_n314), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT64), .ZN(new_n337));
  NOR3_X1   g136(.A1(new_n335), .A2(KEYINPUT34), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT34), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n334), .B2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n330), .A2(new_n333), .A3(new_n337), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT32), .ZN(new_n346));
  XOR2_X1   g145(.A(G71gat), .B(G99gat), .Z(new_n347));
  XNOR2_X1  g146(.A(G15gat), .B(G43gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT33), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT71), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(KEYINPUT71), .A3(new_n351), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n350), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n346), .B1(KEYINPUT33), .B2(new_n349), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n343), .B(new_n344), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G22gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G228gat), .ZN(new_n362));
  INV_X1    g161(.A(G233gat), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G211gat), .B(G218gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(G211gat), .A2(G218gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(G197gat), .A2(G204gat), .ZN(new_n369));
  AND2_X1   g168(.A1(G197gat), .A2(G204gat), .ZN(new_n370));
  OAI22_X1  g169(.A1(new_n368), .A2(KEYINPUT22), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n367), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT3), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n364), .B1(new_n374), .B2(new_n224), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT82), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n372), .B1(new_n269), .B2(new_n373), .ZN(new_n377));
  OR3_X1    g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n364), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n371), .A2(KEYINPUT81), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n382), .A2(new_n383), .A3(new_n365), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n371), .A2(KEYINPUT81), .A3(new_n365), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n373), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n224), .B1(new_n386), .B2(new_n268), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n381), .B1(new_n387), .B2(new_n377), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT31), .B(G50gat), .Z(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n380), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n380), .B2(new_n388), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n361), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n380), .A2(new_n388), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n389), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n388), .A3(new_n390), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n360), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n354), .A2(new_n355), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n398), .A2(new_n346), .A3(new_n349), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n344), .B1(new_n338), .B2(new_n341), .ZN(new_n400));
  INV_X1    g199(.A(new_n357), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AND4_X1   g201(.A1(new_n358), .A2(new_n393), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n372), .ZN(new_n404));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n329), .A2(new_n406), .ZN(new_n407));
  AOI22_X1  g206(.A1(new_n332), .A2(new_n314), .B1(new_n373), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n329), .B1(KEYINPUT29), .B2(new_n406), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n332), .A2(new_n405), .A3(new_n314), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n372), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT74), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT74), .B(new_n404), .C1(new_n407), .C2(new_n408), .ZN(new_n415));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(new_n415), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT30), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n414), .B2(new_n415), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n299), .A2(new_n403), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT35), .ZN(new_n425));
  AOI211_X1 g224(.A(new_n280), .B(new_n205), .C1(new_n288), .C2(new_n289), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n294), .B2(new_n290), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n393), .A2(new_n397), .ZN(new_n428));
  NOR3_X1   g227(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT35), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n421), .B(new_n422), .Z(new_n430));
  NAND3_X1  g229(.A1(new_n399), .A2(new_n343), .A3(new_n401), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n342), .B(new_n339), .C1(new_n356), .C2(new_n357), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n358), .A2(new_n402), .A3(KEYINPUT36), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT36), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n431), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT40), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n277), .A2(new_n259), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n205), .B1(new_n442), .B2(KEYINPUT39), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT39), .B1(new_n257), .B2(new_n259), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n277), .B2(new_n259), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n443), .A2(new_n441), .A3(new_n445), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n447), .A2(new_n448), .A3(new_n297), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n428), .B1(new_n430), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT83), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n412), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n409), .A2(new_n412), .A3(new_n451), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT38), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n419), .A2(KEYINPUT37), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n420), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n422), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n414), .A2(new_n415), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT37), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT38), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n460), .A2(KEYINPUT37), .B1(new_n420), .B2(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT38), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT84), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n427), .A2(new_n459), .A3(new_n464), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n440), .B1(new_n450), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n299), .A2(new_n423), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n428), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n436), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G22gat), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n474), .A2(G1gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT16), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n474), .B1(new_n476), .B2(G1gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(KEYINPUT87), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G8gat), .ZN(new_n479));
  INV_X1    g278(.A(G8gat), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n475), .A2(KEYINPUT87), .A3(new_n480), .A4(new_n477), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G36gat), .ZN(new_n483));
  AND2_X1   g282(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n484));
  NOR2_X1   g283(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G29gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n487), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g288(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(KEYINPUT15), .ZN(new_n491));
  XNOR2_X1  g290(.A(G43gat), .B(G50gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n491), .A2(new_n492), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(KEYINPUT17), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n482), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n479), .A2(KEYINPUT88), .A3(new_n481), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT88), .B1(new_n479), .B2(new_n481), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n495), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n499), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT90), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT18), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT86), .ZN(new_n511));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(G169gat), .B(G197gat), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT12), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(new_n500), .ZN(new_n518));
  INV_X1    g317(.A(new_n503), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n501), .A2(new_n502), .A3(new_n495), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n499), .A2(KEYINPUT18), .A3(new_n500), .A4(new_n503), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n504), .A2(new_n506), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n521), .A3(new_n522), .ZN(new_n525));
  INV_X1    g324(.A(new_n516), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n509), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n473), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G134gat), .B(G162gat), .Z(new_n530));
  AND2_X1   g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(KEYINPUT41), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n530), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT96), .ZN(new_n534));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT93), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(G99gat), .A2(G106gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(G85gat), .ZN(new_n548));
  INV_X1    g347(.A(G92gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(KEYINPUT8), .A2(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n545), .B1(new_n544), .B2(new_n546), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n543), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n537), .A2(KEYINPUT93), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n535), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n553), .B1(new_n560), .B2(new_n551), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n496), .B2(new_n498), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT95), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n495), .A2(new_n562), .B1(KEYINPUT41), .B2(new_n531), .ZN(new_n566));
  XOR2_X1   g365(.A(G190gat), .B(G218gat), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n565), .B2(new_n566), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n534), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n566), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n567), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n533), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n581), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(KEYINPUT9), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n582), .B(KEYINPUT91), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(G57gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(G64gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(G57gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n588), .A2(new_n590), .B1(new_n591), .B2(new_n581), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT91), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n580), .A2(new_n593), .A3(new_n581), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT91), .B1(new_n583), .B2(new_n579), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n586), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G127gat), .B(G155gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI211_X1 g404(.A(new_n502), .B(new_n501), .C1(KEYINPUT21), .C2(new_n597), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n554), .B1(new_n543), .B2(new_n552), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n560), .A2(new_n553), .A3(new_n551), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n597), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n586), .A2(new_n596), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(new_n555), .A3(new_n561), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G230gat), .A2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT98), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n614), .A2(new_n626), .A3(new_n616), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n562), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n619), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(KEYINPUT97), .A3(new_n628), .ZN(new_n632));
  AOI211_X1 g431(.A(new_n621), .B(new_n625), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n625), .B1(new_n621), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n578), .A2(new_n611), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT99), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n611), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n571), .A2(new_n577), .ZN(new_n642));
  INV_X1    g441(.A(new_n637), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT99), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n529), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n299), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g449(.A(KEYINPUT16), .B(G8gat), .Z(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n430), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  OAI21_X1  g452(.A(G8gat), .B1(new_n653), .B2(new_n423), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n652), .ZN(new_n655));
  MUX2_X1   g454(.A(new_n652), .B(new_n655), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g455(.A1(new_n437), .A2(new_n439), .ZN(new_n657));
  OAI21_X1  g456(.A(G15gat), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n433), .A2(G15gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n658), .B1(new_n653), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n647), .A2(new_n428), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n425), .A2(new_n435), .B1(new_n469), .B2(new_n471), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n664), .B1(new_n665), .B2(new_n642), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n464), .A2(new_n467), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n291), .A2(new_n459), .A3(new_n298), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n393), .A2(new_n397), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n448), .A2(new_n297), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n446), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n672), .B2(new_n423), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n657), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n670), .B1(new_n299), .B2(new_n423), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n424), .A2(KEYINPUT35), .B1(new_n429), .B2(new_n434), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT44), .B(new_n578), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n666), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n528), .A2(KEYINPUT100), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n527), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n611), .A2(new_n643), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n487), .B1(new_n686), .B2(new_n648), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n684), .A2(new_n642), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n473), .A2(new_n528), .A3(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(G29gat), .A3(new_n299), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n687), .A2(new_n691), .ZN(G1328gat));
  NAND3_X1  g491(.A1(new_n679), .A2(new_n430), .A3(new_n685), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n483), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n694), .B2(new_n693), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n689), .A2(G36gat), .A3(new_n423), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(G1329gat));
  NAND4_X1  g498(.A1(new_n666), .A2(new_n440), .A3(new_n678), .A4(new_n685), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G43gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n433), .A2(G43gat), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n473), .A2(new_n528), .A3(new_n688), .A4(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n701), .A2(KEYINPUT47), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n703), .B(KEYINPUT103), .Z(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n706), .B2(new_n701), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT104), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  AOI211_X1 g508(.A(new_n709), .B(new_n705), .C1(new_n706), .C2(new_n701), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n704), .B1(new_n708), .B2(new_n710), .ZN(G1330gat));
  NAND3_X1  g510(.A1(new_n679), .A2(new_n428), .A3(new_n685), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n689), .A2(G50gat), .A3(new_n670), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT48), .B1(new_n714), .B2(KEYINPUT105), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1331gat));
  INV_X1    g516(.A(new_n683), .ZN(new_n718));
  NOR4_X1   g517(.A1(new_n718), .A2(new_n611), .A3(new_n578), .A4(new_n643), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n473), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n720), .A2(new_n299), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(new_n587), .ZN(G1332gat));
  XOR2_X1   g521(.A(new_n720), .B(KEYINPUT106), .Z(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n423), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n720), .B2(new_n433), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n440), .A2(G71gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n723), .A2(new_n428), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT107), .B(G78gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n718), .A2(new_n641), .A3(new_n643), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n679), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n299), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n718), .A2(new_n641), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n578), .B(new_n741), .C1(new_n676), .C2(new_n677), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT51), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n473), .A2(KEYINPUT51), .A3(new_n578), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n299), .A2(G85gat), .A3(new_n643), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT108), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n740), .A2(new_n749), .ZN(G1336gat));
  NAND4_X1  g549(.A1(new_n666), .A2(new_n430), .A3(new_n678), .A4(new_n738), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n423), .A2(new_n643), .A3(G92gat), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n754), .B1(new_n744), .B2(new_n745), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(KEYINPUT109), .B2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n755), .A2(KEYINPUT109), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT52), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(KEYINPUT110), .B(KEYINPUT52), .C1(new_n756), .C2(new_n757), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(new_n755), .B2(KEYINPUT111), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n762), .B(new_n752), .C1(KEYINPUT111), .C2(new_n755), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n739), .B2(new_n657), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n433), .A2(G99gat), .A3(new_n643), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n746), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1338gat));
  NOR3_X1   g567(.A1(new_n670), .A2(G106gat), .A3(new_n643), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT112), .Z(new_n770));
  NAND2_X1  g569(.A1(new_n746), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n666), .A2(new_n428), .A3(new_n678), .A4(new_n738), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774));
  AND3_X1   g573(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n774), .B1(new_n771), .B2(new_n773), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT113), .B1(new_n772), .B2(G106gat), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n771), .A2(new_n773), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT114), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n777), .B1(new_n773), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n779), .A2(new_n785), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n509), .A2(new_n523), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n519), .A2(new_n520), .A3(new_n518), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n500), .B1(new_n499), .B2(new_n503), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n515), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n571), .A2(new_n577), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n624), .B1(new_n635), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n627), .A2(KEYINPUT97), .A3(new_n628), .ZN(new_n794));
  AOI21_X1  g593(.A(KEYINPUT97), .B1(new_n627), .B2(new_n628), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n619), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n627), .A2(new_n619), .A3(new_n628), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT54), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n633), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n619), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n629), .A2(new_n792), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n625), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n631), .A2(new_n632), .ZN(new_n805));
  INV_X1    g604(.A(new_n798), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT115), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n798), .B1(new_n631), .B2(new_n632), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  NOR4_X1   g609(.A1(new_n809), .A2(new_n804), .A3(new_n810), .A4(new_n800), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n801), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n791), .A2(KEYINPUT116), .A3(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT116), .B1(new_n791), .B2(new_n812), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n812), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n680), .A2(new_n682), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n787), .A2(new_n790), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(new_n643), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n578), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n611), .B1(new_n815), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n638), .A2(new_n683), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n428), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n648), .A3(new_n434), .ZN(new_n825));
  OAI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n527), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n823), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n648), .A2(new_n403), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n827), .A2(new_n423), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n226), .A3(new_n718), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g630(.A(new_n831), .B(KEYINPUT117), .Z(G1340gat));
  OAI21_X1  g631(.A(G120gat), .B1(new_n825), .B2(new_n643), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n637), .A2(new_n228), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT118), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n825), .B2(new_n611), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n232), .A3(new_n641), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g639(.A(new_n840), .B(KEYINPUT119), .Z(G1342gat));
  INV_X1    g640(.A(G134gat), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n642), .A2(new_n430), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n842), .A3(new_n828), .A4(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT56), .Z(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n825), .B2(new_n642), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  NOR3_X1   g646(.A1(new_n440), .A2(new_n299), .A3(new_n430), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n670), .B1(new_n822), .B2(new_n823), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(KEYINPUT57), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n527), .B1(new_n812), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n801), .B(KEYINPUT120), .C1(new_n808), .C2(new_n811), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n819), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n578), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n611), .B1(new_n856), .B2(new_n815), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n851), .B(new_n670), .C1(new_n857), .C2(new_n823), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n848), .B1(new_n850), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G141gat), .B1(new_n859), .B2(new_n527), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n849), .A2(new_n648), .A3(new_n657), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n430), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n527), .A2(G141gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n718), .B(new_n848), .C1(new_n850), .C2(new_n858), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n867), .A2(G141gat), .B1(new_n862), .B2(new_n863), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(G1344gat));
  OAI21_X1  g669(.A(G148gat), .B1(new_n859), .B2(new_n643), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(G148gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n862), .A2(new_n874), .A3(new_n637), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n848), .A2(new_n637), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n640), .A2(new_n645), .A3(new_n527), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n791), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n816), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n855), .B2(new_n578), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n641), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI211_X1 g682(.A(KEYINPUT122), .B(new_n880), .C1(new_n855), .C2(new_n578), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n851), .B1(new_n885), .B2(new_n670), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n670), .A2(new_n851), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n827), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n876), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n873), .B(new_n875), .C1(new_n889), .C2(new_n890), .ZN(G1345gat));
  OAI21_X1  g690(.A(G155gat), .B1(new_n859), .B2(new_n611), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n862), .A2(new_n210), .A3(new_n641), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n859), .B2(new_n642), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n843), .A2(new_n211), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n861), .B2(new_n896), .ZN(G1347gat));
  INV_X1    g696(.A(new_n433), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n648), .A2(new_n423), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n824), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n527), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n648), .B1(new_n822), .B2(new_n823), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n403), .A2(new_n430), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT123), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n905), .A2(G169gat), .A3(new_n683), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n906), .A2(new_n907), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  OAI21_X1  g709(.A(G176gat), .B1(new_n900), .B2(new_n643), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n643), .A2(G176gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n911), .B1(new_n905), .B2(new_n912), .ZN(G1349gat));
  INV_X1    g712(.A(new_n905), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n310), .A3(new_n641), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n900), .B2(new_n611), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n918));
  XOR2_X1   g717(.A(new_n917), .B(new_n918), .Z(G1350gat));
  NAND3_X1  g718(.A1(new_n914), .A2(new_n311), .A3(new_n578), .ZN(new_n920));
  OAI21_X1  g719(.A(G190gat), .B1(new_n900), .B2(new_n642), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(KEYINPUT61), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(KEYINPUT61), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(G1351gat));
  NOR3_X1   g723(.A1(new_n440), .A2(new_n423), .A3(new_n670), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n902), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(G197gat), .B1(new_n927), .B2(new_n718), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n899), .A2(new_n657), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n929), .B1(new_n886), .B2(new_n888), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n528), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  AOI21_X1  g732(.A(G204gat), .B1(new_n933), .B2(KEYINPUT62), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n927), .A2(new_n637), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n933), .A2(KEYINPUT62), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n930), .A2(new_n637), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G204gat), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1353gat));
  OR3_X1    g739(.A1(new_n926), .A2(G211gat), .A3(new_n611), .ZN(new_n941));
  INV_X1    g740(.A(new_n929), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n881), .A2(new_n882), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n611), .A3(new_n884), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n877), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT57), .B1(new_n945), .B2(new_n428), .ZN(new_n946));
  INV_X1    g745(.A(new_n888), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n641), .B(new_n942), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n941), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952));
  INV_X1    g751(.A(G218gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n953), .B1(new_n930), .B2(new_n578), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n926), .A2(G218gat), .A3(new_n642), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n578), .B(new_n942), .C1(new_n946), .C2(new_n947), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G218gat), .ZN(new_n958));
  INV_X1    g757(.A(new_n955), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n958), .A2(KEYINPUT127), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n956), .A2(new_n960), .ZN(G1355gat));
endmodule


