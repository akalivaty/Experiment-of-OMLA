//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1201, new_n1202, new_n1203;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(new_n469), .B1(G113), .B2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(KEYINPUT66), .A3(G125), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n472), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n467), .A2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n462), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n481));
  OAI22_X1  g056(.A1(new_n478), .A2(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(G136), .B2(new_n473), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT67), .ZN(G162));
  NAND3_X1  g059(.A1(new_n467), .A2(G126), .A3(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n467), .A2(new_n462), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n473), .A2(new_n492), .A3(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT68), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n495), .A3(G543), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OR3_X1    g078(.A1(new_n502), .A2(KEYINPUT69), .A3(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT69), .B1(new_n502), .B2(new_n503), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  INV_X1    g081(.A(new_n496), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n499), .B1(new_n495), .B2(G543), .ZN(new_n508));
  NOR3_X1   g083(.A1(new_n497), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  OR2_X1    g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n497), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(G88), .B1(G50), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n504), .A2(new_n505), .A3(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  XNOR2_X1  g092(.A(KEYINPUT70), .B(KEYINPUT7), .ZN(new_n518));
  AND3_X1   g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n501), .A2(G89), .A3(new_n506), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n514), .A2(G51), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n526));
  AND2_X1   g101(.A1(G77), .A2(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n501), .B2(G64), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n526), .B1(new_n528), .B2(new_n503), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n514), .A2(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n510), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  AOI211_X1 g109(.A(new_n534), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n535));
  OAI211_X1 g110(.A(KEYINPUT71), .B(G651), .C1(new_n535), .C2(new_n527), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n529), .A2(new_n533), .A3(new_n536), .ZN(G171));
  XOR2_X1   g112(.A(KEYINPUT73), .B(G43), .Z(new_n538));
  AOI22_X1  g113(.A1(new_n511), .A2(G81), .B1(new_n514), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n501), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n540), .A2(KEYINPUT72), .ZN(new_n541));
  OAI21_X1  g116(.A(G651), .B1(new_n540), .B2(KEYINPUT72), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  INV_X1    g124(.A(new_n513), .ZN(new_n550));
  NOR2_X1   g125(.A1(KEYINPUT6), .A2(G651), .ZN(new_n551));
  OAI211_X1 g126(.A(G53), .B(G543), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n554), .A2(KEYINPUT74), .ZN(new_n555));
  NOR3_X1   g130(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n498), .A2(new_n500), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n557), .A2(G65), .A3(new_n507), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n556), .B1(new_n560), .B2(G651), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n510), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n501), .A2(KEYINPUT76), .A3(new_n506), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(G91), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n554), .B1(new_n552), .B2(KEYINPUT74), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n552), .A2(new_n553), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n561), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G299));
  OAI21_X1  g145(.A(G651), .B1(new_n535), .B2(new_n527), .ZN(new_n571));
  AOI21_X1  g146(.A(new_n532), .B1(new_n571), .B2(new_n526), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(new_n536), .ZN(G301));
  OR2_X1    g148(.A1(new_n501), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G49), .B2(new_n514), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n563), .A2(G87), .A3(new_n564), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n563), .A2(G86), .A3(new_n564), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n563), .A2(KEYINPUT79), .A3(G86), .A4(new_n564), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  OAI211_X1 g159(.A(G61), .B(new_n507), .C1(new_n508), .C2(new_n509), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n584), .B1(new_n587), .B2(G651), .ZN(new_n588));
  AOI211_X1 g163(.A(KEYINPUT77), .B(new_n503), .C1(new_n585), .C2(new_n586), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n583), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n586), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n501), .B2(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT77), .B1(new_n592), .B2(new_n503), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI211_X1 g169(.A(new_n594), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n595));
  OAI211_X1 g170(.A(new_n584), .B(G651), .C1(new_n595), .C2(new_n591), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n596), .A3(KEYINPUT78), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n514), .A2(G48), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n582), .A2(new_n590), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(KEYINPUT80), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n596), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n583), .A2(new_n602), .B1(new_n580), .B2(new_n581), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n597), .A2(new_n598), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n600), .A2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n503), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n514), .A2(G47), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n510), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n563), .A2(G92), .A3(new_n564), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g192(.A1(new_n563), .A2(KEYINPUT10), .A3(G92), .A4(new_n564), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n501), .A2(G66), .ZN(new_n620));
  INV_X1    g195(.A(G79), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n497), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n622), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n614), .B1(new_n625), .B2(G868), .ZN(G284));
  OAI21_X1  g201(.A(new_n614), .B1(new_n625), .B2(G868), .ZN(G321));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n569), .B2(G868), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(new_n569), .B2(G868), .ZN(G280));
  XNOR2_X1  g205(.A(KEYINPUT81), .B(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n625), .B1(G860), .B2(new_n631), .ZN(G148));
  OAI21_X1  g207(.A(KEYINPUT82), .B1(new_n544), .B2(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n631), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  MUX2_X1   g210(.A(KEYINPUT82), .B(new_n633), .S(new_n635), .Z(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n467), .A2(new_n474), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT83), .B(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n473), .A2(G135), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n646), .C1(new_n647), .C2(new_n478), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n643), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT15), .B(G2435), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2438), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2430), .Z(new_n654));
  AOI21_X1  g229(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n653), .B2(new_n654), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2451), .B(G2454), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n656), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n663), .A2(G14), .A3(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n668), .B(KEYINPUT17), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n670), .C1(new_n667), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n667), .A3(new_n669), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n683), .A2(new_n684), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n682), .A2(new_n687), .A3(new_n685), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n690));
  AOI211_X1 g265(.A(new_n686), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n689), .B2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(G1981), .B(G1986), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(G229));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT32), .B(G1981), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NOR2_X1   g279(.A1(G16), .A2(G22), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G166), .B2(G16), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1971), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT33), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(KEYINPUT33), .ZN(new_n714));
  OR3_X1    g289(.A1(new_n713), .A2(G1976), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(G1976), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n707), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n703), .A2(new_n704), .A3(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT34), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n708), .A2(G24), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT88), .Z(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n612), .B2(new_n708), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT89), .B(G1986), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(KEYINPUT90), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT87), .B(G29), .Z(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G25), .ZN(new_n730));
  INV_X1    g305(.A(new_n478), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G119), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n473), .A2(G131), .ZN(new_n733));
  OR2_X1    g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(new_n729), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(KEYINPUT36), .ZN(new_n743));
  AND3_X1   g318(.A1(new_n726), .A2(new_n727), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n719), .A2(new_n720), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n742), .A2(KEYINPUT36), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT26), .Z(new_n750));
  INV_X1    g325(.A(G129), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n478), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n474), .A2(G105), .ZN(new_n753));
  INV_X1    g328(.A(G141), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n489), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G29), .B2(G32), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT27), .B(G1996), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT96), .ZN(new_n762));
  INV_X1    g337(.A(G33), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G29), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT25), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n467), .A2(G127), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n462), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n770));
  AOI211_X1 g345(.A(new_n766), .B(new_n770), .C1(G139), .C2(new_n473), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n764), .B1(new_n773), .B2(G29), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(new_n442), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(new_n442), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(G34), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n777), .A2(G34), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n729), .ZN(new_n780));
  AOI22_X1  g355(.A1(G160), .A2(G29), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G2084), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n762), .A2(new_n775), .A3(new_n776), .A4(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT97), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(KEYINPUT97), .ZN(new_n785));
  NOR2_X1   g360(.A1(G171), .A2(new_n708), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G5), .B2(new_n708), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT100), .Z(new_n790));
  NAND3_X1  g365(.A1(new_n784), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n708), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n544), .B2(new_n708), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1341), .Z(new_n794));
  NAND2_X1  g369(.A1(new_n708), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n624), .A2(G16), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n708), .A2(G4), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G1348), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n794), .B(new_n798), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n729), .A2(G35), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G162), .B2(new_n729), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT29), .Z(new_n806));
  INV_X1    g381(.A(G2090), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n787), .A2(new_n788), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n759), .A2(new_n760), .B1(G2084), .B2(new_n781), .ZN(new_n812));
  NOR2_X1   g387(.A1(G168), .A2(new_n708), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n708), .B2(G21), .ZN(new_n814));
  INV_X1    g389(.A(G1966), .ZN(new_n815));
  NOR2_X1   g390(.A1(G164), .A2(new_n728), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G27), .B2(new_n728), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n814), .A2(new_n815), .B1(new_n443), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n443), .B2(new_n817), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n728), .A2(G26), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT28), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n731), .A2(G128), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT92), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n825));
  INV_X1    g400(.A(G116), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G2105), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(G140), .B2(new_n473), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n821), .B1(new_n829), .B2(G29), .ZN(new_n830));
  INV_X1    g405(.A(G2067), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT31), .B(G11), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT98), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT99), .B(G28), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n835), .A2(KEYINPUT30), .ZN(new_n836));
  AOI21_X1  g411(.A(G29), .B1(new_n835), .B2(KEYINPUT30), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI221_X1 g413(.A(new_n838), .B1(new_n648), .B2(new_n728), .C1(new_n814), .C2(new_n815), .ZN(new_n839));
  NOR4_X1   g414(.A1(new_n812), .A2(new_n819), .A3(new_n832), .A4(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n801), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(G1348), .B2(new_n841), .ZN(new_n842));
  NOR4_X1   g417(.A1(new_n791), .A2(new_n803), .A3(new_n811), .A4(new_n842), .ZN(new_n843));
  AND3_X1   g418(.A1(new_n747), .A2(new_n748), .A3(new_n843), .ZN(G311));
  NAND3_X1  g419(.A1(new_n747), .A2(new_n748), .A3(new_n843), .ZN(G150));
  AND3_X1   g420(.A1(new_n557), .A2(G67), .A3(new_n507), .ZN(new_n846));
  AND2_X1   g421(.A1(G80), .A2(G543), .ZN(new_n847));
  OAI211_X1 g422(.A(KEYINPUT101), .B(G651), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n847), .B1(new_n501), .B2(G67), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n850), .B2(new_n503), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n501), .A2(G93), .A3(new_n506), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n514), .A2(G55), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n848), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT102), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n848), .A2(new_n851), .A3(new_n854), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  NAND2_X1  g436(.A1(new_n625), .A2(G559), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT38), .Z(new_n863));
  NAND3_X1  g438(.A1(new_n856), .A2(new_n543), .A3(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n544), .A2(new_n855), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n863), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n861), .B1(new_n869), .B2(new_n871), .ZN(G145));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n473), .A2(G142), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n462), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  INV_X1    g451(.A(G130), .ZN(new_n877));
  OAI221_X1 g452(.A(new_n874), .B1(new_n875), .B2(new_n876), .C1(new_n877), .C2(new_n478), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n639), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n829), .B(G164), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n737), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n491), .A2(new_n493), .ZN(new_n882));
  INV_X1    g457(.A(new_n488), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n829), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n736), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n879), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n881), .A2(new_n886), .A3(new_n879), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n773), .A2(new_n757), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n756), .B2(new_n773), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n889), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n894), .B2(new_n887), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G160), .B(new_n648), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(G162), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n873), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT103), .A4(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n896), .B2(new_n899), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n599), .A2(KEYINPUT80), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n603), .A2(new_n604), .A3(new_n601), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n909), .A2(new_n910), .A3(G303), .ZN(new_n911));
  AOI21_X1  g486(.A(G303), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  XNOR2_X1  g487(.A(G290), .B(G288), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NOR3_X1   g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(G166), .B1(new_n600), .B2(new_n605), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n909), .A2(new_n910), .A3(G303), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n908), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n914), .B1(new_n911), .B2(new_n912), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n913), .A3(new_n917), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT104), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n907), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT42), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n866), .B(new_n634), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n569), .A2(new_n619), .A3(new_n623), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n566), .A2(new_n567), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n503), .B1(new_n558), .B2(new_n559), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n928), .A2(new_n929), .A3(new_n556), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n619), .A2(new_n623), .B1(new_n565), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n927), .B2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n624), .A2(G299), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n569), .A2(new_n619), .A3(new_n623), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n933), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n925), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n940), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n923), .B2(new_n924), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(G868), .ZN(new_n945));
  INV_X1    g520(.A(new_n859), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(G868), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n906), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  AOI211_X1 g524(.A(KEYINPUT105), .B(new_n947), .C1(new_n944), .C2(G868), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(G295));
  NAND2_X1  g526(.A1(new_n945), .A2(new_n948), .ZN(G331));
  INV_X1    g527(.A(G37), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n920), .A2(KEYINPUT104), .A3(new_n921), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT104), .B1(new_n920), .B2(new_n921), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G286), .B1(new_n572), .B2(new_n536), .ZN(new_n957));
  AND4_X1   g532(.A1(G286), .A2(new_n529), .A3(new_n533), .A4(new_n536), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n959), .A2(new_n864), .A3(new_n865), .ZN(new_n960));
  INV_X1    g535(.A(new_n957), .ZN(new_n961));
  INV_X1    g536(.A(new_n958), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n864), .A2(new_n865), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n935), .B(new_n938), .C1(new_n960), .C2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n935), .A2(new_n938), .ZN(new_n967));
  INV_X1    g542(.A(new_n959), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n866), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n959), .A2(new_n864), .A3(new_n865), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(new_n971), .A3(KEYINPUT106), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n960), .A2(new_n963), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n932), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n966), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n953), .B1(new_n956), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n964), .A2(KEYINPUT107), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n967), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n979), .A3(new_n974), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(new_n919), .A3(new_n922), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT108), .B1(new_n976), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n919), .A2(new_n922), .ZN(new_n985));
  INV_X1    g560(.A(new_n975), .ZN(new_n986));
  AOI21_X1  g561(.A(G37), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n982), .A4(new_n981), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n969), .A2(new_n932), .A3(new_n970), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n973), .A2(new_n939), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(KEYINPUT106), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(new_n966), .C1(new_n954), .C2(new_n955), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n975), .A2(new_n919), .A3(new_n922), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n953), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT43), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n984), .A2(new_n989), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n982), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n987), .A2(KEYINPUT43), .A3(new_n981), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  MUX2_X1   g575(.A(new_n997), .B(new_n1000), .S(KEYINPUT44), .Z(G397));
  AOI21_X1  g576(.A(G1384), .B1(new_n882), .B2(new_n883), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n472), .A2(new_n1006), .A3(new_n476), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n829), .B(new_n831), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n756), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT125), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1008), .A2(G1996), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT46), .Z(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1015));
  XNOR2_X1  g590(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(G1996), .B1(new_n752), .B2(new_n755), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1009), .A2(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1012), .A2(KEYINPUT112), .A3(new_n757), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT112), .B1(new_n1012), .B2(new_n757), .ZN(new_n1020));
  OAI22_X1  g595(.A1(new_n1018), .A2(new_n1008), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT113), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1008), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n737), .A2(new_n739), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n736), .A2(new_n740), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1022), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(G290), .A2(G1986), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(new_n1008), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT48), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1016), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n824), .A2(new_n831), .A3(new_n828), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1008), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n569), .B(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(G1384), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n884), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1007), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1956), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1047), .A2(new_n1007), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT114), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1050), .B(new_n1003), .C1(G164), .C2(G1384), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT56), .B(G2072), .ZN(new_n1052));
  XOR2_X1   g627(.A(new_n1052), .B(KEYINPUT119), .Z(new_n1053));
  NAND4_X1  g628(.A1(new_n1048), .A2(new_n1049), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1039), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n470), .A2(new_n471), .ZN(new_n1056));
  OAI211_X1 g631(.A(G40), .B(new_n475), .C1(new_n1056), .C2(new_n462), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1002), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n831), .A2(new_n1059), .B1(new_n1044), .B2(new_n802), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(new_n624), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1049), .A2(new_n1051), .A3(new_n1007), .A4(new_n1047), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1053), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1046), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1038), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT58), .B(G1341), .Z(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1063), .B2(G1996), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT120), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1070), .C1(new_n1063), .C2(G1996), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1068), .B1(new_n1075), .B2(new_n544), .ZN(new_n1076));
  AOI211_X1 g651(.A(KEYINPUT59), .B(new_n543), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1055), .A2(new_n1066), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT61), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1060), .A2(new_n624), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT60), .B1(new_n1082), .B2(new_n1061), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1055), .A2(new_n1066), .A3(KEYINPUT61), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1060), .A2(new_n1085), .A3(new_n625), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1081), .A2(new_n1083), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1067), .B1(new_n1078), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1063), .B2(G2078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT45), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(G164), .B2(G1384), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1091), .A2(new_n1007), .A3(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1089), .A2(G2078), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1094), .A2(new_n1095), .B1(new_n1044), .B2(new_n788), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1090), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n1097), .B2(G171), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1044), .A2(new_n788), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(G40), .B(new_n1095), .C1(new_n475), .C2(KEYINPUT123), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n1102), .B(new_n472), .C1(KEYINPUT123), .C2(new_n475), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1047), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1101), .B(new_n1090), .C1(new_n1005), .C2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1105), .B2(G171), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1097), .A2(G171), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT121), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1097), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1109), .B(new_n1110), .C1(new_n1105), .C2(G171), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1106), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT116), .B1(new_n1094), .B2(G1966), .ZN(new_n1114));
  INV_X1    g689(.A(G2084), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1007), .A2(new_n1042), .A3(new_n1115), .A4(new_n1043), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1091), .A2(new_n1007), .A3(new_n1093), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1117), .A2(new_n1118), .A3(new_n815), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1114), .A2(G168), .A3(new_n1116), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1120), .A2(new_n1121), .A3(G8), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1119), .A2(new_n1116), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1118), .B1(new_n1117), .B2(new_n815), .ZN(new_n1124));
  OAI21_X1  g699(.A(G286), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(new_n1120), .A3(G8), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1122), .B1(KEYINPUT51), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G8), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1059), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(G1976), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(G288), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n710), .B2(G1976), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(KEYINPUT52), .B2(new_n1131), .ZN(new_n1135));
  INV_X1    g710(.A(G86), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n598), .B1(new_n510), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(G1981), .B1(new_n602), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n599), .B2(G1981), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT49), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1139), .A2(new_n1142), .A3(new_n1140), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1141), .B(new_n1129), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G1971), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1007), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1063), .A2(new_n1146), .B1(new_n1147), .B2(new_n807), .ZN(new_n1148));
  AND3_X1   g723(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1148), .A2(new_n1151), .A3(new_n1128), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1151), .B1(new_n1148), .B2(new_n1128), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1135), .A2(new_n1145), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1127), .A2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1088), .A2(new_n1113), .A3(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1135), .A2(new_n1145), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1148), .A2(new_n1128), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1151), .A2(KEYINPUT117), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1159), .B(new_n1160), .Z(new_n1161));
  NOR2_X1   g736(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1162), .A2(new_n1128), .A3(G286), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1158), .A2(new_n1161), .A3(KEYINPUT63), .A4(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1163), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1155), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1164), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1145), .A2(new_n1130), .A3(new_n710), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(G1981), .B2(new_n599), .ZN(new_n1170));
  AOI22_X1  g745(.A1(new_n1170), .A2(new_n1129), .B1(new_n1158), .B2(new_n1152), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1128), .B1(new_n1162), .B2(G168), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1121), .B1(new_n1172), .B2(new_n1125), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT62), .B1(new_n1173), .B2(new_n1122), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1155), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1122), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1126), .A2(KEYINPUT51), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1157), .A2(new_n1168), .A3(new_n1171), .A4(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT110), .ZN(new_n1184));
  NAND2_X1  g759(.A1(G290), .A2(G1986), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1029), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1186), .B(new_n1023), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT111), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1027), .A2(new_n1188), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1182), .A2(new_n1183), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1183), .B1(new_n1182), .B2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1036), .B1(new_n1190), .B2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1194));
  NOR3_X1   g768(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1195));
  OAI21_X1  g769(.A(new_n1195), .B1(new_n698), .B2(new_n699), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n902), .B2(new_n903), .ZN(new_n1197));
  AND3_X1   g771(.A1(new_n997), .A2(new_n1194), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1194), .B1(new_n997), .B2(new_n1197), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n1199), .ZN(G308));
  NAND2_X1  g774(.A1(new_n997), .A2(new_n1197), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1201), .A2(KEYINPUT127), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n997), .A2(new_n1197), .A3(new_n1194), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1202), .A2(new_n1203), .ZN(G225));
endmodule


