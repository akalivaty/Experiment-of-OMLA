//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939;
  XOR2_X1   g000(.A(KEYINPUT95), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT94), .B(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT15), .ZN(new_n205));
  NOR2_X1   g004(.A1(G29gat), .A2(G36gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT14), .ZN(new_n207));
  OR3_X1    g006(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n204), .B2(new_n207), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(new_n211), .A3(new_n209), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT17), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n215), .ZN(new_n218));
  XOR2_X1   g017(.A(new_n218), .B(G8gat), .Z(new_n219));
  XOR2_X1   g018(.A(KEYINPUT96), .B(KEYINPUT17), .Z(new_n220));
  OAI211_X1 g019(.A(new_n214), .B(new_n219), .C1(new_n213), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n213), .A2(new_n219), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT18), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n221), .A2(KEYINPUT18), .A3(new_n222), .A4(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n213), .A2(new_n219), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n222), .B(KEYINPUT13), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G169gat), .B(G197gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT93), .ZN(new_n234));
  INV_X1    g033(.A(G113gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT92), .B(KEYINPUT11), .Z(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G141gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n236), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(KEYINPUT12), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n231), .A4(new_n240), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT97), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(KEYINPUT97), .A3(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT27), .B(G183gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT27), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(G183gat), .ZN(new_n254));
  INV_X1    g053(.A(G183gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT27), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT69), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G190gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT28), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OR2_X1    g061(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n263));
  NAND2_X1  g062(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(G183gat), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g067(.A(new_n265), .B(new_n259), .C1(new_n268), .C2(new_n253), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n262), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(KEYINPUT26), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT26), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n277), .A2(new_n283), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n276), .A2(KEYINPUT65), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT65), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n278), .B2(KEYINPUT23), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n275), .B1(KEYINPUT23), .B2(new_n278), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT24), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n294), .A2(new_n296), .B1(new_n255), .B2(new_n259), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n285), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n280), .A2(new_n282), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT23), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT25), .B1(new_n273), .B2(new_n274), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n301), .B1(new_n287), .B2(new_n289), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n266), .A2(new_n259), .A3(new_n267), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n294), .A2(new_n296), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n272), .A2(new_n284), .B1(new_n298), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G134gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G127gat), .ZN(new_n309));
  INV_X1    g108(.A(G127gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G134gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT70), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(KEYINPUT70), .B2(new_n311), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n235), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(G113gat), .A2(G120gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT1), .B1(new_n317), .B2(KEYINPUT71), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n313), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT73), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT73), .B1(new_n309), .B2(new_n311), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT72), .ZN(new_n326));
  AND2_X1   g125(.A1(G113gat), .A2(G120gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(G113gat), .A2(G120gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n315), .A2(KEYINPUT72), .A3(new_n316), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n325), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT73), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n310), .A2(G134gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n308), .A2(G127gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT73), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT1), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(new_n330), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT74), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n321), .B1(new_n333), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n307), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n307), .A2(new_n342), .ZN(new_n345));
  INV_X1    g144(.A(G227gat), .ZN(new_n346));
  INV_X1    g145(.A(G233gat), .ZN(new_n347));
  OAI22_X1  g146(.A1(new_n344), .A2(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT34), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT34), .ZN(new_n350));
  OAI221_X1 g149(.A(new_n350), .B1(new_n346), .B2(new_n347), .C1(new_n344), .C2(new_n345), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(G15gat), .B(G43gat), .Z(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT67), .B(G183gat), .Z(new_n358));
  AOI21_X1  g157(.A(G190gat), .B1(new_n358), .B2(KEYINPUT27), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT28), .B1(new_n359), .B2(new_n265), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n260), .B1(new_n252), .B2(new_n257), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n284), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n298), .A2(new_n306), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n332), .B1(new_n325), .B2(new_n331), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n339), .A2(KEYINPUT74), .A3(new_n340), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n320), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n368), .A2(new_n343), .A3(G227gat), .A4(G233gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT75), .B(KEYINPUT33), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n357), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n369), .B(KEYINPUT32), .C1(new_n370), .C2(new_n357), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n352), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n352), .B1(new_n373), .B2(new_n374), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT36), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT36), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n373), .A2(new_n374), .ZN(new_n380));
  INV_X1    g179(.A(new_n352), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n352), .A2(new_n373), .A3(KEYINPUT78), .A4(new_n374), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G141gat), .B(G148gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT2), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(G155gat), .B2(G162gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G155gat), .B(G162gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n394), .B(new_n389), .C1(new_n390), .C2(new_n392), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(KEYINPUT3), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n396), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n388), .B1(new_n342), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n365), .A2(new_n366), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n397), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n402), .A2(new_n403), .A3(new_n321), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n367), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n401), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n404), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n342), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n367), .A2(new_n404), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT84), .A3(new_n412), .ZN(new_n413));
  OR3_X1    g212(.A1(new_n367), .A2(KEYINPUT84), .A3(new_n404), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n388), .A3(new_n414), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n401), .B(KEYINPUT83), .C1(new_n405), .C2(new_n406), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n409), .A2(KEYINPUT5), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n412), .A2(KEYINPUT4), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT85), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n367), .A2(new_n402), .A3(new_n404), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n367), .A2(KEYINPUT85), .A3(new_n402), .A4(new_n404), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n342), .A2(new_n400), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n388), .A2(KEYINPUT5), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G1gat), .B(G29gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT0), .ZN(new_n429));
  XNOR2_X1  g228(.A(G57gat), .B(G85gat), .ZN(new_n430));
  XOR2_X1   g229(.A(new_n429), .B(new_n430), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n431), .A3(new_n426), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT86), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n431), .B1(new_n417), .B2(new_n426), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT86), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT6), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n436), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G8gat), .B(G36gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(G64gat), .B(G92gat), .ZN(new_n444));
  XOR2_X1   g243(.A(new_n443), .B(new_n444), .Z(new_n445));
  XNOR2_X1  g244(.A(G211gat), .B(G218gat), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G197gat), .B(G204gat), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT22), .ZN(new_n450));
  INV_X1    g249(.A(G211gat), .ZN(new_n451));
  INV_X1    g250(.A(G218gat), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n446), .B(KEYINPUT79), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n456), .A2(new_n458), .A3(KEYINPUT80), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n464), .B(KEYINPUT81), .Z(new_n465));
  NAND2_X1  g264(.A1(new_n277), .A2(new_n283), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n293), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n271), .B2(new_n262), .ZN(new_n468));
  INV_X1    g267(.A(new_n297), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n290), .A3(new_n291), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n299), .A2(KEYINPUT23), .B1(new_n304), .B2(new_n303), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n470), .A2(new_n285), .B1(new_n471), .B2(new_n302), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n465), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT29), .B1(new_n362), .B2(new_n363), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n463), .B(new_n473), .C1(new_n474), .C2(new_n465), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n465), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n307), .B2(KEYINPUT29), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n463), .B1(new_n478), .B2(new_n473), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n445), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n461), .A2(new_n462), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n474), .A2(new_n465), .ZN(new_n482));
  INV_X1    g281(.A(new_n473), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n445), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n475), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n486), .A3(KEYINPUT30), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n488), .B(new_n445), .C1(new_n476), .C2(new_n479), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n442), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n399), .A2(KEYINPUT29), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n481), .A2(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n459), .A2(KEYINPUT29), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT3), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n404), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G78gat), .B(G106gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n493), .B2(new_n496), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G228gat), .A2(G233gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(G22gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G50gat), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n504), .B(new_n505), .Z(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n500), .A2(new_n501), .A3(new_n506), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n386), .B1(new_n491), .B2(new_n510), .ZN(new_n511));
  AND4_X1   g310(.A1(new_n440), .A2(new_n427), .A3(KEYINPUT6), .A4(new_n432), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n440), .B1(new_n439), .B2(KEYINPUT6), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT37), .B1(new_n476), .B2(new_n479), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n484), .A2(new_n516), .A3(new_n475), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n445), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT38), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n480), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n517), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(new_n519), .A3(new_n485), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n518), .A2(KEYINPUT89), .A3(new_n519), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n427), .A2(KEYINPUT88), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT88), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n417), .A2(new_n528), .A3(new_n426), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n432), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n435), .A2(new_n434), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n526), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n510), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n387), .B1(new_n421), .B2(new_n424), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n431), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n388), .B1(new_n413), .B2(new_n414), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT87), .B1(new_n541), .B2(KEYINPUT40), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n490), .B1(new_n541), .B2(KEYINPUT40), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT40), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n544), .B(new_n545), .C1(new_n538), .C2(new_n540), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n542), .A2(new_n543), .A3(new_n530), .A4(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n533), .A2(new_n534), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n511), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n510), .B1(new_n384), .B2(new_n383), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n442), .A2(new_n490), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT35), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n514), .A2(new_n532), .ZN(new_n553));
  INV_X1    g352(.A(new_n490), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n376), .B2(new_n377), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n380), .A2(new_n381), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT90), .A3(new_n375), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n553), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n552), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n549), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT91), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n562), .A3(KEYINPUT91), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n249), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT101), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(KEYINPUT102), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT7), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G99gat), .B(G106gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  OAI211_X1 g378(.A(new_n214), .B(new_n579), .C1(new_n213), .C2(new_n220), .ZN(new_n580));
  INV_X1    g379(.A(new_n213), .ZN(new_n581));
  INV_X1    g380(.A(new_n579), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n581), .A2(new_n582), .B1(KEYINPUT41), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n570), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n569), .A2(KEYINPUT102), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT103), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n585), .A2(new_n589), .ZN(new_n595));
  OR3_X1    g394(.A1(new_n591), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G57gat), .B(G64gat), .Z(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G71gat), .B(G78gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n597), .A2(new_n601), .B1(new_n602), .B2(KEYINPUT98), .ZN(new_n603));
  INV_X1    g402(.A(new_n602), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT98), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n604), .A2(new_n597), .A3(new_n605), .A4(new_n601), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n310), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n609), .B(KEYINPUT100), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT21), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n219), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n616), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT99), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G155gat), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n617), .A2(new_n618), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n623), .B1(new_n617), .B2(new_n618), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G230gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n347), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n609), .B1(KEYINPUT104), .B2(new_n578), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n582), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT10), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n614), .A2(new_n631), .A3(new_n579), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n628), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n629), .B(new_n579), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n635), .B1(new_n628), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n638), .B(new_n639), .Z(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n637), .B(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n594), .B1(new_n591), .B2(new_n595), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n596), .A2(new_n626), .A3(new_n642), .A4(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n567), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n442), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n647), .B(G1gat), .Z(G1324gat));
  OAI21_X1  g447(.A(G8gat), .B1(new_n646), .B2(new_n490), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT106), .Z(new_n650));
  NOR2_X1   g449(.A1(new_n646), .A2(new_n490), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT42), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT16), .B(G8gat), .Z(new_n653));
  AND4_X1   g452(.A1(KEYINPUT105), .A2(new_n651), .A3(new_n652), .A4(new_n653), .ZN(new_n654));
  OR3_X1    g453(.A1(new_n646), .A2(KEYINPUT105), .A3(new_n490), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n655), .A2(new_n652), .B1(new_n651), .B2(new_n653), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n654), .B2(new_n656), .ZN(G1325gat));
  INV_X1    g456(.A(new_n386), .ZN(new_n658));
  OAI21_X1  g457(.A(G15gat), .B1(new_n646), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n556), .A2(new_n558), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(G15gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n659), .B1(new_n646), .B2(new_n662), .ZN(G1326gat));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n534), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT43), .B(G22gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1327gat));
  INV_X1    g465(.A(KEYINPUT45), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n637), .B(new_n640), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n626), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n596), .A2(new_n643), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n567), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n442), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n203), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n667), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n674), .A2(new_n667), .A3(new_n676), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n565), .A2(new_n566), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n671), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n563), .A2(KEYINPUT107), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n549), .B2(new_n562), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n671), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n682), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n244), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(new_n442), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n677), .B(new_n678), .C1(new_n693), .C2(new_n203), .ZN(G1328gat));
  AND4_X1   g493(.A1(new_n554), .A2(new_n567), .A3(new_n202), .A4(new_n673), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT46), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n692), .A2(new_n490), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n202), .ZN(G1329gat));
  NAND2_X1  g497(.A1(new_n386), .A2(G43gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n674), .A2(new_n661), .ZN(new_n700));
  OAI22_X1  g499(.A1(new_n692), .A2(new_n699), .B1(G43gat), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  INV_X1    g502(.A(new_n691), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n534), .B(new_n704), .C1(new_n681), .C2(new_n688), .ZN(new_n705));
  INV_X1    g504(.A(G50gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n567), .A2(new_n706), .A3(new_n510), .A4(new_n673), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n705), .B2(new_n706), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT48), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  OAI221_X1 g510(.A(new_n708), .B1(new_n703), .B2(KEYINPUT48), .C1(new_n705), .C2(new_n706), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(G1331gat));
  NOR2_X1   g512(.A1(new_n682), .A2(new_n684), .ZN(new_n714));
  INV_X1    g513(.A(new_n626), .ZN(new_n715));
  NOR4_X1   g514(.A1(new_n671), .A2(new_n715), .A3(new_n244), .A4(new_n642), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n675), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  OAI22_X1  g519(.A1(new_n717), .A2(new_n490), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n554), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT109), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n717), .B2(new_n658), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n660), .A2(new_n599), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n717), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g528(.A1(new_n717), .A2(new_n534), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT110), .B(G78gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1335gat));
  NAND2_X1  g531(.A1(new_n690), .A2(new_n715), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n642), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n689), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735), .B2(new_n442), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n733), .A2(new_n672), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n563), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT51), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT51), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n563), .A2(new_n740), .A3(new_n737), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n742), .A2(new_n574), .A3(new_n675), .A4(new_n668), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(G1336gat));
  NOR2_X1   g543(.A1(new_n490), .A2(G92gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n668), .A3(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n689), .A2(new_n554), .A3(new_n734), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n752), .A2(G92gat), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n740), .A2(KEYINPUT111), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n738), .B(new_n754), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n755), .A2(new_n668), .A3(new_n745), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n756), .B1(new_n752), .B2(G92gat), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n751), .A2(new_n753), .B1(new_n757), .B2(new_n749), .ZN(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n735), .B2(new_n658), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n661), .A2(G99gat), .A3(new_n642), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT113), .Z(new_n761));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(G1338gat));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n534), .A2(G106gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n739), .A2(new_n668), .A3(new_n741), .A4(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n767), .B2(new_n766), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n685), .B1(new_n679), .B2(new_n671), .ZN(new_n770));
  OAI211_X1 g569(.A(new_n510), .B(new_n734), .C1(new_n770), .C2(new_n687), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G106gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n771), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT114), .B1(new_n771), .B2(G106gat), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n642), .A2(G106gat), .A3(new_n534), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n755), .A2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n755), .A2(KEYINPUT115), .A3(new_n776), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n774), .A2(new_n775), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n773), .B1(new_n782), .B2(new_n764), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n637), .A2(new_n640), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n640), .B1(new_n635), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n636), .A2(KEYINPUT10), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n788), .A2(new_n633), .B1(new_n627), .B2(new_n347), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n632), .A2(new_n628), .A3(new_n634), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(KEYINPUT54), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n785), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT55), .B1(new_n787), .B2(new_n791), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n784), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n794), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n796), .A2(KEYINPUT118), .A3(new_n785), .A4(new_n792), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n797), .A3(new_n244), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n222), .B1(new_n221), .B2(new_n223), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n229), .A2(new_n230), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n239), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n243), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n668), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n671), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  AND4_X1   g603(.A1(new_n671), .A2(new_n795), .A3(new_n802), .A4(new_n797), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n715), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n645), .B2(new_n690), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n644), .A2(new_n808), .A3(new_n244), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n442), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n811), .A2(new_n534), .A3(new_n559), .ZN(new_n812));
  OAI21_X1  g611(.A(G113gat), .B1(new_n812), .B2(new_n249), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT119), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n811), .A2(new_n550), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n554), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n235), .A3(new_n244), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(G1340gat));
  NOR3_X1   g617(.A1(new_n812), .A2(new_n314), .A3(new_n642), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(new_n668), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n314), .ZN(G1341gat));
  NAND3_X1  g620(.A1(new_n816), .A2(new_n310), .A3(new_n626), .ZN(new_n822));
  OAI21_X1  g621(.A(G127gat), .B1(new_n812), .B2(new_n715), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1342gat));
  NAND2_X1  g623(.A1(new_n671), .A2(new_n490), .ZN(new_n825));
  OR3_X1    g624(.A1(new_n815), .A2(G134gat), .A3(new_n825), .ZN(new_n826));
  OR2_X1    g625(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n827));
  OAI21_X1  g626(.A(G134gat), .B1(new_n812), .B2(new_n672), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(KEYINPUT56), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G1343gat));
  OR2_X1    g629(.A1(new_n811), .A2(KEYINPUT121), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n811), .A2(KEYINPUT121), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n831), .A2(new_n510), .A3(new_n658), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n554), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n249), .A2(G141gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n386), .A2(new_n442), .A3(new_n554), .ZN(new_n838));
  XOR2_X1   g637(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n806), .A2(new_n810), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n510), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n793), .A2(new_n794), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n242), .A2(KEYINPUT97), .A3(new_n243), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT97), .B1(new_n242), .B2(new_n243), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n671), .B1(new_n847), .B2(new_n803), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n715), .B1(new_n848), .B2(new_n805), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n843), .B(new_n534), .C1(new_n849), .C2(new_n810), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n838), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n249), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n837), .A3(new_n852), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n851), .A2(new_n690), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n834), .A2(new_n835), .B1(new_n854), .B2(G141gat), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n837), .ZN(G1344gat));
  XNOR2_X1  g655(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n645), .A2(KEYINPUT123), .A3(new_n246), .A4(new_n247), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n248), .B2(new_n644), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n803), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n248), .B2(new_n844), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n671), .A2(new_n802), .ZN(new_n864));
  INV_X1    g663(.A(new_n844), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n863), .A2(new_n671), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n861), .B1(new_n866), .B2(new_n715), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n843), .B1(new_n867), .B2(new_n534), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n841), .A2(new_n510), .A3(new_n840), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n870), .A2(new_n668), .A3(new_n838), .ZN(new_n871));
  INV_X1    g670(.A(G148gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n857), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(KEYINPUT59), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n851), .B2(new_n642), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n834), .A2(new_n872), .A3(new_n668), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1345gat));
  INV_X1    g677(.A(G155gat), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n834), .A2(new_n879), .A3(new_n626), .ZN(new_n880));
  OAI21_X1  g679(.A(G155gat), .B1(new_n851), .B2(new_n715), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n851), .B2(new_n672), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n825), .A2(G162gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n833), .B2(new_n884), .ZN(G1347gat));
  AOI211_X1 g684(.A(new_n675), .B(new_n490), .C1(new_n806), .C2(new_n810), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(new_n550), .ZN(new_n887));
  AOI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n244), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n534), .A3(new_n660), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(new_n273), .A3(new_n249), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n888), .A2(new_n890), .ZN(G1348gat));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n274), .A3(new_n668), .ZN(new_n892));
  OAI21_X1  g691(.A(G176gat), .B1(new_n889), .B2(new_n642), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT124), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n887), .A2(new_n258), .A3(new_n626), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n268), .B1(new_n889), .B2(new_n715), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n896), .A2(new_n897), .B1(KEYINPUT125), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(KEYINPUT125), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n899), .B(new_n900), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n889), .B2(new_n672), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT61), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n259), .A3(new_n671), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(G1351gat));
  NOR3_X1   g704(.A1(new_n675), .A2(new_n386), .A3(new_n490), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n864), .A2(new_n865), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n715), .B1(new_n848), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n860), .A3(new_n858), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n510), .ZN(new_n910));
  AOI211_X1 g709(.A(new_n534), .B(new_n839), .C1(new_n806), .C2(new_n810), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n248), .B(new_n906), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n870), .A2(new_n914), .A3(new_n248), .A4(new_n906), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n913), .A2(new_n915), .A3(G197gat), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n886), .A2(new_n510), .A3(new_n658), .ZN(new_n917));
  INV_X1    g716(.A(G197gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n244), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n916), .A2(KEYINPUT127), .A3(new_n919), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1352gat));
  INV_X1    g723(.A(G204gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n925), .A3(new_n668), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n870), .A2(new_n906), .ZN(new_n928));
  OAI21_X1  g727(.A(G204gat), .B1(new_n928), .B2(new_n642), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(KEYINPUT62), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(G1353gat));
  NAND3_X1  g730(.A1(new_n917), .A2(new_n451), .A3(new_n626), .ZN(new_n932));
  OAI21_X1  g731(.A(G211gat), .B1(new_n928), .B2(new_n715), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(G1354gat));
  OAI21_X1  g736(.A(G218gat), .B1(new_n928), .B2(new_n672), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n452), .A3(new_n671), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1355gat));
endmodule


