//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n549, new_n550, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT66), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2105), .ZN(new_n457));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(G125), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n457), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n457), .C1(new_n458), .C2(new_n459), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n462), .A2(new_n467), .ZN(G160));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n457), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G136), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n457), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  OR2_X1    g051(.A1(G100), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G112), .C2(new_n457), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n472), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  OAI211_X1 g055(.A(G126), .B(G2105), .C1(new_n458), .C2(new_n459), .ZN(new_n481));
  INV_X1    g056(.A(G114), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n458), .B2(new_n459), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n469), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n485), .B1(new_n489), .B2(new_n491), .ZN(G164));
  INV_X1    g067(.A(G651), .ZN(new_n493));
  AND2_X1   g068(.A1(KEYINPUT5), .A2(G543), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT5), .A2(G543), .ZN(new_n495));
  OAI21_X1  g070(.A(G62), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n496), .A2(KEYINPUT69), .B1(G75), .B2(G543), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G62), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n493), .B1(new_n497), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT68), .A3(G50), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(G50), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n498), .A2(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(new_n514), .B1(G88), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n504), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(G89), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n495), .A2(new_n494), .B1(new_n510), .B2(new_n511), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT70), .B(G51), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n508), .A2(new_n527), .B1(new_n500), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  AOI22_X1  g106(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n493), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n506), .A2(new_n507), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n522), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n533), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n493), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n535), .A2(new_n542), .B1(new_n522), .B2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(KEYINPUT9), .B1(new_n535), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n508), .A2(new_n552), .A3(new_n555), .A4(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n494), .A2(new_n495), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(new_n515), .B2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n557), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G74), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n498), .A2(new_n565), .A3(new_n499), .ZN(new_n566));
  AOI22_X1  g141(.A1(G49), .A2(new_n508), .B1(new_n566), .B2(G651), .ZN(new_n567));
  INV_X1    g142(.A(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT74), .B1(new_n522), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n500), .A2(new_n534), .A3(new_n570), .A4(G87), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(G288));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  OAI211_X1 g148(.A(G48), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n522), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(G61), .B1(new_n494), .B2(new_n495), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n493), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n573), .B1(new_n576), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n498), .B2(new_n499), .ZN(new_n582));
  INV_X1    g157(.A(new_n578), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n500), .A2(new_n534), .A3(G86), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n584), .A2(KEYINPUT75), .A3(new_n585), .A4(new_n574), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(new_n493), .ZN(new_n590));
  INV_X1    g165(.A(G47), .ZN(new_n591));
  INV_X1    g166(.A(G85), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n535), .A2(new_n591), .B1(new_n522), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n515), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n559), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n508), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n596), .B1(new_n605), .B2(G868), .ZN(G321));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NAND2_X1  g183(.A1(G299), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G168), .B2(new_n608), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n605), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n605), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI22_X1  g190(.A1(new_n615), .A2(KEYINPUT77), .B1(G868), .B2(new_n545), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(KEYINPUT77), .B2(new_n615), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n469), .A2(new_n464), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT80), .B(G2100), .Z(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n475), .A2(G123), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT81), .ZN(new_n627));
  INV_X1    g202(.A(G2096), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n471), .B2(G135), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n627), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n623), .A2(new_n624), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n627), .A2(new_n632), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G2096), .ZN(new_n636));
  NAND4_X1  g211(.A1(new_n625), .A2(new_n633), .A3(new_n634), .A4(new_n636), .ZN(G156));
  INV_X1    g212(.A(G14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n644), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n638), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n649), .A2(new_n650), .ZN(new_n655));
  AOI21_X1  g230(.A(KEYINPUT82), .B1(new_n655), .B2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n657));
  AOI211_X1 g232(.A(new_n657), .B(new_n653), .C1(new_n649), .C2(new_n650), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n657), .B1(new_n651), .B2(new_n653), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n655), .A2(KEYINPUT82), .A3(new_n652), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n664), .A2(KEYINPUT83), .A3(new_n654), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n661), .A2(new_n665), .ZN(G401));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT84), .ZN(new_n668));
  NOR2_X1   g243(.A1(G2072), .A2(G2078), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n442), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2084), .B(G2090), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n668), .A2(new_n670), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n670), .B(KEYINPUT17), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n671), .C1(new_n668), .C2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n671), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n668), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n628), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT85), .B(G2100), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(G2096), .ZN(new_n683));
  INV_X1    g258(.A(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT88), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1956), .B(G2474), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT86), .ZN(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(new_n691), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n693), .A2(new_n694), .ZN(new_n697));
  MUX2_X1   g272(.A(new_n691), .B(new_n696), .S(new_n697), .Z(new_n698));
  NOR2_X1   g273(.A1(new_n695), .A2(new_n691), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n702), .B1(new_n698), .B2(new_n701), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n689), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(new_n689), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n707), .A2(new_n708), .A3(new_n703), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n706), .A2(new_n709), .A3(new_n711), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(G229));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n580), .B2(new_n586), .ZN(new_n717));
  NOR2_X1   g292(.A1(G6), .A2(G16), .ZN(new_n718));
  OR3_X1    g293(.A1(new_n717), .A2(KEYINPUT91), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(KEYINPUT91), .B1(new_n717), .B2(new_n718), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT32), .B(G1981), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(new_n722), .A3(new_n720), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n716), .A2(G22), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G166), .B2(new_n716), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G1971), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT33), .B(G1976), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT93), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G288), .A2(G16), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT92), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n716), .A2(G23), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n734), .B1(new_n733), .B2(new_n735), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n732), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(new_n738), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n740), .A2(new_n731), .A3(new_n736), .ZN(new_n741));
  INV_X1    g316(.A(G1971), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n742), .B(new_n727), .C1(G166), .C2(new_n716), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n729), .A2(new_n739), .A3(new_n741), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n726), .A2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT34), .ZN(new_n746));
  OAI21_X1  g321(.A(KEYINPUT94), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT89), .B(G29), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n749), .A2(G25), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n471), .A2(G131), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n475), .A2(G119), .ZN(new_n752));
  OR2_X1    g327(.A1(G95), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G107), .C2(new_n457), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n750), .B1(new_n756), .B2(new_n749), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT35), .B(G1991), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n716), .A2(G24), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n594), .B2(new_n716), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT90), .B(G1986), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n759), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n745), .B2(new_n746), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n766), .B(KEYINPUT34), .C1(new_n726), .C2(new_n744), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n747), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(KEYINPUT36), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT36), .ZN(new_n770));
  NAND4_X1  g345(.A1(new_n747), .A2(new_n765), .A3(new_n770), .A4(new_n767), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G160), .A2(G29), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT24), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n774), .A2(G34), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n774), .A2(G34), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n748), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT98), .Z(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n716), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n716), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n779), .A2(new_n780), .B1(new_n782), .B2(G1966), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G1966), .B2(new_n782), .ZN(new_n784));
  INV_X1    g359(.A(G29), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G32), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n475), .A2(G129), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n464), .A2(G105), .ZN(new_n791));
  INV_X1    g366(.A(G141), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n470), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n790), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT99), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n786), .B1(new_n796), .B2(new_n785), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT100), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT27), .B(G1996), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n784), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  NOR2_X1   g376(.A1(G16), .A2(G19), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n545), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1341), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n785), .A2(G33), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT25), .ZN(new_n807));
  NAND2_X1  g382(.A1(G103), .A2(G2104), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G2105), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n457), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n471), .A2(G139), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n469), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(new_n457), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n806), .B1(new_n814), .B2(new_n785), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT97), .B(G2072), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n716), .A2(G4), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n605), .B2(new_n716), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n817), .B1(new_n819), .B2(G1348), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(G1348), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n475), .A2(G128), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n457), .A2(G116), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n824));
  INV_X1    g399(.A(G140), .ZN(new_n825));
  OAI221_X1 g400(.A(new_n822), .B1(new_n823), .B2(new_n824), .C1(new_n825), .C2(new_n470), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G29), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n748), .A2(G26), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G2067), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n821), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n805), .A2(new_n820), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT31), .B(G11), .Z(new_n836));
  INV_X1    g411(.A(G28), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT30), .ZN(new_n838));
  AOI21_X1  g413(.A(G29), .B1(new_n837), .B2(KEYINPUT30), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n836), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(G171), .A2(new_n716), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G5), .B2(new_n716), .ZN(new_n842));
  INV_X1    g417(.A(G1961), .ZN(new_n843));
  OAI221_X1 g418(.A(new_n840), .B1(new_n635), .B2(new_n748), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n748), .A2(G35), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G162), .B2(new_n748), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT29), .B(G2090), .Z(new_n847));
  XOR2_X1   g422(.A(new_n846), .B(new_n847), .Z(new_n848));
  AND2_X1   g423(.A1(new_n842), .A2(new_n843), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n749), .A2(G27), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(G164), .B2(new_n749), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(G2078), .ZN(new_n852));
  NOR4_X1   g427(.A1(new_n844), .A2(new_n848), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n716), .A2(G20), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT101), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT23), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G299), .B2(G16), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT102), .B(G1956), .Z(new_n858));
  XOR2_X1   g433(.A(new_n857), .B(new_n858), .Z(new_n859));
  OR2_X1    g434(.A1(new_n779), .A2(new_n780), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n835), .A2(new_n853), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n801), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n772), .A2(KEYINPUT103), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT103), .B1(new_n772), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(G311));
  NAND2_X1  g440(.A1(new_n772), .A2(new_n862), .ZN(G150));
  NAND2_X1  g441(.A1(new_n605), .A2(G559), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT38), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n515), .A2(G93), .B1(new_n508), .B2(G55), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT104), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(new_n493), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n545), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(new_n545), .A3(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n868), .B(new_n877), .Z(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n879), .A2(new_n880), .A3(G860), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n873), .A2(G860), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT37), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n881), .A2(new_n883), .ZN(G145));
  XNOR2_X1  g459(.A(new_n479), .B(G160), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n635), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n475), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n457), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(G142), .ZN(new_n891));
  OAI221_X1 g466(.A(new_n888), .B1(new_n889), .B2(new_n890), .C1(new_n891), .C2(new_n470), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT107), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n755), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n826), .B(G164), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n621), .B(KEYINPUT106), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n893), .B(new_n756), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n489), .A2(new_n491), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n481), .A2(new_n484), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n826), .B(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(new_n896), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n899), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n794), .A2(KEYINPUT105), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n907));
  INV_X1    g482(.A(new_n794), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n814), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n906), .A2(new_n909), .B1(new_n795), .B2(new_n814), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n898), .A2(new_n905), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n898), .B2(new_n905), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n887), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n898), .A2(new_n905), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n898), .A2(new_n905), .A3(new_n911), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n886), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(G37), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n921), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT40), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT40), .B1(new_n922), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(G395));
  XOR2_X1   g501(.A(G303), .B(G288), .Z(new_n927));
  NAND2_X1  g502(.A1(G305), .A2(G290), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n587), .A2(new_n594), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G303), .B(G288), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n928), .A3(new_n929), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(KEYINPUT109), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT110), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n877), .B(new_n614), .Z(new_n937));
  XNOR2_X1  g512(.A(new_n604), .B(G299), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n877), .B(new_n614), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n938), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n946), .A3(new_n943), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n936), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n936), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n873), .A2(new_n608), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(G295));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n951), .ZN(G331));
  NAND2_X1  g528(.A1(G286), .A2(G301), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n525), .A2(G171), .A3(new_n526), .A4(new_n529), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n938), .B1(new_n877), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n875), .A2(new_n876), .A3(new_n954), .A4(new_n955), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n877), .A2(new_n956), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OR2_X1    g536(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n934), .B(new_n959), .C1(new_n964), .C2(new_n940), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n965), .A2(new_n919), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n959), .B1(new_n964), .B2(new_n940), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n931), .A2(new_n933), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT112), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT43), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n938), .B(new_n961), .C1(new_n962), .C2(new_n963), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n940), .B1(new_n960), .B2(new_n958), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  AND4_X1   g549(.A1(KEYINPUT43), .A2(new_n974), .A3(new_n919), .A4(new_n965), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT44), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT43), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n966), .B2(new_n970), .ZN(new_n979));
  AND4_X1   g554(.A1(new_n978), .A2(new_n974), .A3(new_n919), .A4(new_n965), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n976), .A2(new_n981), .ZN(G397));
  INV_X1    g557(.A(G1384), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n902), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n462), .A2(new_n467), .A3(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n984), .A2(new_n985), .A3(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT46), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT126), .Z(new_n992));
  XNOR2_X1  g567(.A(new_n826), .B(G2067), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n908), .B(new_n993), .C1(KEYINPUT46), .C2(new_n990), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT47), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n795), .A2(G1996), .A3(new_n988), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT113), .Z(new_n998));
  AND2_X1   g573(.A1(new_n989), .A2(new_n993), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n988), .A2(new_n990), .A3(new_n794), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT114), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n756), .A2(new_n758), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n756), .A2(new_n758), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n989), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n988), .A2(G1986), .A3(G290), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1009));
  XNOR2_X1  g584(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n996), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n826), .A2(G2067), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT125), .ZN(new_n1014));
  OR2_X1    g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n988), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n594), .B(G1986), .Z(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n989), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1002), .A2(new_n1019), .A3(new_n1006), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n985), .B1(G164), .B2(G1384), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n902), .A2(KEYINPUT45), .A3(new_n983), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n987), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G1966), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n1026));
  AOI21_X1  g601(.A(G1384), .B1(new_n900), .B2(new_n901), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1026), .A2(new_n1029), .A3(new_n780), .A4(new_n987), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(G168), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(G168), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT51), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1031), .A2(new_n1035), .A3(G8), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT62), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT62), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1034), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(G1981), .B1(new_n576), .B2(new_n579), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n584), .A2(new_n1042), .A3(new_n585), .A4(new_n574), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT117), .B(KEYINPUT49), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT118), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1027), .B2(new_n987), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1051), .A3(new_n1046), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1041), .A2(new_n1043), .A3(KEYINPUT49), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1048), .A2(new_n1050), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G288), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(KEYINPUT116), .A3(new_n1057), .ZN(new_n1061));
  OR2_X1    g636(.A1(G288), .A2(new_n1055), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1050), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1054), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n509), .A2(new_n514), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n515), .A2(G88), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(G8), .B1(new_n1069), .B2(new_n503), .ZN(new_n1070));
  NAND2_X1  g645(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1071), .ZN(new_n1074));
  OAI221_X1 g649(.A(G8), .B1(new_n1073), .B2(new_n1074), .C1(new_n1069), .C2(new_n503), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n987), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1078));
  NOR3_X1   g653(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2090), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1080), .A2(new_n1081), .B1(new_n1023), .B2(new_n742), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1077), .B1(new_n1082), .B2(new_n1049), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n987), .B1(new_n1027), .B2(KEYINPUT45), .ZN(new_n1084));
  NOR3_X1   g659(.A1(G164), .A2(new_n985), .A3(G1384), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n742), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1026), .A2(new_n1029), .A3(new_n1081), .A4(new_n987), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(G8), .A3(new_n1076), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1066), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G2078), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1021), .A2(new_n1022), .A3(new_n1091), .A4(new_n987), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n843), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT53), .B1(new_n1092), .B2(new_n1096), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1094), .B(new_n1095), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1090), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1038), .A2(new_n1040), .A3(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1043), .B(KEYINPUT120), .ZN(new_n1103));
  NOR2_X1   g678(.A1(G288), .A2(G1976), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1054), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(new_n1050), .B(KEYINPUT119), .Z(new_n1106));
  NAND3_X1  g681(.A1(new_n1054), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1089), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1049), .B(G286), .C1(new_n1025), .C2(new_n1030), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1066), .A2(new_n1083), .A3(new_n1089), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT63), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI221_X4 g687(.A(new_n1049), .B1(new_n1072), .B2(new_n1075), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(new_n1107), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1114), .A2(KEYINPUT63), .A3(new_n1083), .A4(new_n1109), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1108), .B1(new_n1112), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1102), .A2(new_n1116), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1066), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1095), .B1(new_n1093), .B2(new_n1092), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1094), .ZN(new_n1120));
  OAI21_X1  g695(.A(G171), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1094), .A2(G301), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1121), .B(KEYINPUT54), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1037), .A2(new_n1118), .A3(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1123), .A2(new_n1119), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT54), .B1(new_n1100), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1956), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT57), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n557), .A2(new_n1131), .A3(new_n562), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n557), .B2(new_n562), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1021), .A2(new_n1022), .A3(new_n987), .A4(new_n1135), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT121), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1027), .A2(new_n987), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1027), .B2(new_n987), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n832), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1348), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT122), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1141), .A2(new_n1146), .A3(new_n1143), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1145), .A2(new_n605), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1134), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1137), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1027), .A2(new_n987), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT121), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1027), .A2(new_n987), .A3(new_n1138), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1021), .A2(new_n1022), .A3(new_n990), .A4(new_n987), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n874), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1160), .B(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1147), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1146), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1164));
  OAI211_X1 g739(.A(KEYINPUT60), .B(new_n604), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1130), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1151), .A2(KEYINPUT61), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1134), .B1(new_n1130), .B2(new_n1136), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1137), .B2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1162), .A2(new_n1165), .A3(new_n1167), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT60), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1145), .A2(new_n1173), .A3(new_n1147), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1172), .A2(new_n1174), .A3(new_n605), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1153), .B1(new_n1171), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1128), .A2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g752(.A(KEYINPUT124), .B(new_n1020), .C1(new_n1117), .C2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1180));
  AOI211_X1 g755(.A(KEYINPUT59), .B(new_n874), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1170), .B(new_n1167), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g757(.A(new_n1173), .B(new_n605), .C1(new_n1145), .C2(new_n1147), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1172), .A2(new_n1174), .A3(new_n605), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1152), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1090), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1100), .A2(new_n1126), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT54), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1190), .A3(new_n1124), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1102), .B(new_n1116), .C1(new_n1186), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1020), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1179), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1017), .B1(new_n1178), .B2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NAND4_X1  g770(.A1(new_n686), .A2(new_n713), .A3(G319), .A4(new_n714), .ZN(new_n1197));
  AOI21_X1  g771(.A(new_n1197), .B1(new_n661), .B2(new_n665), .ZN(new_n1198));
  INV_X1    g772(.A(new_n923), .ZN(new_n1199));
  NOR2_X1   g773(.A1(new_n920), .A2(new_n921), .ZN(new_n1200));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g775(.A1(new_n979), .A2(new_n980), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n1201), .A2(new_n1202), .ZN(G308));
  OAI221_X1 g777(.A(new_n1198), .B1(new_n1199), .B2(new_n1200), .C1(new_n979), .C2(new_n980), .ZN(G225));
endmodule


