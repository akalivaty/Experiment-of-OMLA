//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n546, new_n547, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1109, new_n1110;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n452), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2106), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n458), .A2(new_n459), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  AND2_X1   g040(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT3), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(G137), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n470), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT67), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n475), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n474), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n468), .A2(new_n470), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n475), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  INV_X1    g059(.A(new_n482), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n475), .ZN(new_n486));
  INV_X1    g061(.A(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(new_n475), .B2(G112), .ZN(new_n489));
  OAI221_X1 g064(.A(new_n484), .B1(new_n486), .B2(new_n487), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n470), .A2(new_n476), .A3(G138), .A4(new_n475), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT4), .A2(G138), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n468), .A2(new_n475), .A3(new_n470), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n470), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT69), .Z(new_n511));
  OR2_X1    g086(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n507), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n516), .A2(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n511), .A2(new_n521), .ZN(G166));
  AOI22_X1  g097(.A1(new_n518), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(new_n514), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(G51), .B2(new_n509), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n509), .A2(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n519), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n517), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  INV_X1    g113(.A(new_n509), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n519), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G188));
  XNOR2_X1  g123(.A(KEYINPUT70), .B(KEYINPUT9), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n509), .A2(G53), .A3(new_n549), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI21_X1  g127(.A(KEYINPUT9), .B1(new_n539), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n519), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n514), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n556), .A2(G91), .B1(G651), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n555), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G171), .ZN(G301));
  XNOR2_X1  g137(.A(new_n528), .B(KEYINPUT72), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G286));
  INV_X1    g139(.A(G166), .ZN(G303));
  NAND2_X1  g140(.A1(new_n556), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n509), .A2(G49), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  AOI22_X1  g144(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n570), .A2(new_n517), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n509), .A2(G48), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n519), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n517), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n556), .A2(G85), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n509), .A2(G47), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(KEYINPUT73), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n556), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  AOI22_X1  g161(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(new_n517), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n509), .A2(KEYINPUT74), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(G54), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n586), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n563), .B2(new_n596), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n563), .B2(new_n596), .ZN(G280));
  XNOR2_X1  g174(.A(KEYINPUT75), .B(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(G860), .B2(new_n600), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n470), .A2(new_n476), .ZN(new_n606));
  NOR4_X1   g181(.A1(new_n606), .A2(G2105), .A3(new_n467), .A4(new_n466), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT12), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(G2100), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n483), .A2(G123), .ZN(new_n611));
  INV_X1    g186(.A(G135), .ZN(new_n612));
  NOR2_X1   g187(.A1(G99), .A2(G2105), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n614));
  OAI221_X1 g189(.A(new_n611), .B1(new_n486), .B2(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(G2096), .Z(new_n616));
  NAND2_X1  g191(.A1(new_n610), .A2(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2430), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2435), .ZN(new_n619));
  XOR2_X1   g194(.A(G2427), .B(G2438), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT14), .ZN(new_n622));
  XOR2_X1   g197(.A(G2451), .B(G2454), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n622), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n627), .B(new_n628), .Z(new_n629));
  AND2_X1   g204(.A1(new_n629), .A2(G14), .ZN(G401));
  XOR2_X1   g205(.A(G2072), .B(G2078), .Z(new_n631));
  XOR2_X1   g206(.A(G2067), .B(G2678), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2084), .B(G2090), .Z(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n631), .B1(new_n635), .B2(KEYINPUT18), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2100), .Z(new_n638));
  AND2_X1   g213(.A1(new_n635), .A2(KEYINPUT17), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n633), .A2(new_n634), .ZN(new_n640));
  AOI21_X1  g215(.A(KEYINPUT18), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(G227));
  XOR2_X1   g217(.A(G1956), .B(G2474), .Z(new_n643));
  XOR2_X1   g218(.A(G1961), .B(G1966), .Z(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1971), .B(G1976), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT19), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n643), .A2(new_n644), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n654));
  OAI211_X1 g229(.A(new_n653), .B(new_n654), .C1(new_n652), .C2(new_n651), .ZN(new_n655));
  XOR2_X1   g230(.A(G1991), .B(G1996), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT76), .B(G1986), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G1981), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n659), .B(new_n661), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G229));
  INV_X1    g238(.A(G16), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G4), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n593), .B2(new_n664), .ZN(new_n666));
  INV_X1    g241(.A(G1348), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G29), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G26), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT28), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n483), .A2(G128), .ZN(new_n672));
  NOR2_X1   g247(.A1(G104), .A2(G2105), .ZN(new_n673));
  OAI21_X1  g248(.A(G2104), .B1(new_n475), .B2(G116), .ZN(new_n674));
  INV_X1    g249(.A(G140), .ZN(new_n675));
  OAI221_X1 g250(.A(new_n672), .B1(new_n673), .B2(new_n674), .C1(new_n675), .C2(new_n486), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G29), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n677), .A2(KEYINPUT81), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(KEYINPUT81), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G2067), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(G16), .A2(G19), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n542), .B2(G16), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(G1341), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n668), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT82), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n664), .A2(KEYINPUT23), .A3(G20), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n689));
  INV_X1    g264(.A(G20), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G299), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n688), .B(new_n691), .C1(new_n692), .C2(new_n664), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1956), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n669), .A2(G33), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT25), .Z(new_n698));
  INV_X1    g273(.A(G139), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n486), .B2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT83), .Z(new_n701));
  NAND2_X1  g276(.A1(G115), .A2(G2104), .ZN(new_n702));
  INV_X1    g277(.A(G127), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n606), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(G2105), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n696), .B1(new_n705), .B2(new_n669), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(G2072), .Z(new_n707));
  NOR2_X1   g282(.A1(G29), .A2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n483), .A2(G129), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT86), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(G2105), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT88), .Z(new_n717));
  AOI21_X1  g292(.A(new_n708), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n615), .A2(new_n669), .ZN(new_n721));
  NAND2_X1  g296(.A1(G171), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G5), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G1961), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT84), .B(KEYINPUT24), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G34), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G29), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G160), .B2(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G2084), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT85), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(G1966), .ZN(new_n733));
  NAND2_X1  g308(.A1(G168), .A2(G16), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G16), .B2(G21), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n721), .B(new_n732), .C1(new_n733), .C2(new_n735), .ZN(new_n736));
  NAND4_X1  g311(.A1(new_n695), .A2(new_n707), .A3(new_n720), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n669), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n669), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G2078), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n740), .B1(G2084), .B2(new_n729), .C1(new_n735), .C2(new_n733), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n669), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n669), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT29), .Z(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n739), .A2(G2078), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT89), .B(G28), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(new_n669), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n746), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n741), .B(new_n751), .C1(new_n745), .C2(new_n744), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n730), .A2(new_n731), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n752), .B(new_n753), .C1(new_n724), .C2(new_n723), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT31), .B(G11), .Z(new_n755));
  NOR3_X1   g330(.A1(new_n737), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT90), .Z(new_n757));
  NOR2_X1   g332(.A1(G16), .A2(G23), .ZN(new_n758));
  INV_X1    g333(.A(G288), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT33), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1976), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n664), .A2(G6), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n575), .B2(new_n664), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT32), .B(G1981), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT78), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n764), .B(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G22), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G166), .B2(G16), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT79), .B(G1971), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n762), .A2(new_n767), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT34), .ZN(new_n773));
  MUX2_X1   g348(.A(G24), .B(G290), .S(G16), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT77), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G1986), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n483), .A2(G119), .ZN(new_n777));
  NOR2_X1   g352(.A1(G95), .A2(G2105), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n779));
  INV_X1    g354(.A(G131), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n777), .B1(new_n778), .B2(new_n779), .C1(new_n780), .C2(new_n486), .ZN(new_n781));
  MUX2_X1   g356(.A(G25), .B(new_n781), .S(G29), .Z(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT35), .B(G1991), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n775), .A2(G1986), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n776), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n773), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(KEYINPUT80), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT36), .Z(new_n791));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n788), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n757), .A2(new_n793), .ZN(G311));
  INV_X1    g369(.A(G311), .ZN(G150));
  NAND2_X1  g370(.A1(G80), .A2(G543), .ZN(new_n796));
  INV_X1    g371(.A(G67), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n514), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G651), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n556), .A2(G93), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n509), .A2(G55), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G860), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT37), .Z(new_n805));
  OR2_X1    g380(.A1(new_n803), .A2(KEYINPUT92), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n803), .A2(KEYINPUT92), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n542), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n806), .A2(new_n542), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n593), .A2(G559), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT93), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n815), .B2(KEYINPUT39), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n805), .B1(new_n817), .B2(new_n819), .ZN(G145));
  NAND2_X1  g395(.A1(new_n494), .A2(new_n496), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n501), .A2(KEYINPUT94), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n498), .A2(new_n823), .A3(new_n500), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n821), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n676), .B(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n717), .B(new_n826), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(new_n705), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n826), .B(new_n716), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n705), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  NOR2_X1   g408(.A1(G106), .A2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n486), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G130), .B2(new_n483), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n781), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n832), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n615), .B(G160), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n490), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT96), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n608), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n839), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g422(.A1(new_n803), .A2(new_n596), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n812), .B(KEYINPUT97), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n602), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n593), .A2(G299), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n592), .A2(new_n692), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT98), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT41), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  MUX2_X1   g432(.A(new_n852), .B(new_n853), .S(KEYINPUT99), .Z(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n858), .B2(new_n856), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n855), .B1(new_n850), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT42), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n575), .B(KEYINPUT100), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G166), .ZN(new_n863));
  XNOR2_X1  g438(.A(G290), .B(new_n759), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n861), .B(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n848), .B1(new_n868), .B2(new_n596), .ZN(G295));
  OAI21_X1  g444(.A(new_n848), .B1(new_n868), .B2(new_n596), .ZN(G331));
  NOR2_X1   g445(.A1(new_n528), .A2(G171), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(G286), .B2(G171), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n812), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n853), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(new_n865), .C1(new_n859), .C2(new_n874), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(new_n845), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n853), .A2(new_n856), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n873), .B(new_n878), .C1(new_n856), .C2(new_n858), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n865), .B(KEYINPUT102), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n879), .B(new_n880), .C1(new_n854), .C2(new_n873), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n877), .A2(KEYINPUT43), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n875), .B1(new_n859), .B2(new_n874), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n880), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT43), .B1(new_n877), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT44), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n877), .A2(new_n884), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT43), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n877), .A2(new_n881), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(KEYINPUT43), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n886), .B1(new_n891), .B2(KEYINPUT44), .ZN(G397));
  NOR2_X1   g467(.A1(new_n825), .A2(G1384), .ZN(new_n893));
  XOR2_X1   g468(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT104), .B1(G160), .B2(G40), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  INV_X1    g472(.A(G40), .ZN(new_n898));
  NOR4_X1   g473(.A1(new_n474), .A2(new_n480), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n895), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(G1996), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n717), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n904), .A2(KEYINPUT105), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n676), .B(new_n681), .ZN(new_n908));
  INV_X1    g483(.A(new_n716), .ZN(new_n909));
  INV_X1    g484(.A(G1996), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI211_X1 g486(.A(new_n905), .B(new_n906), .C1(new_n907), .C2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n781), .B(new_n783), .Z(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n901), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(G290), .B(G1986), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(G303), .A2(G8), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT55), .Z(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT107), .Z(new_n919));
  INV_X1    g494(.A(G8), .ZN(new_n920));
  NOR2_X1   g495(.A1(G164), .A2(G1384), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT50), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n900), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n825), .B2(G1384), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n498), .A2(new_n823), .A3(new_n500), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n823), .B1(new_n498), .B2(new_n500), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n497), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT50), .B1(new_n926), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n745), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n893), .A2(KEYINPUT45), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n900), .C1(new_n921), .C2(new_n894), .ZN(new_n938));
  INV_X1    g513(.A(G1971), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n920), .B1(new_n936), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n919), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n918), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n896), .B(new_n899), .C1(new_n921), .C2(new_n922), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n926), .A2(KEYINPUT50), .A3(new_n931), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n745), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n940), .A3(KEYINPUT111), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G8), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT111), .B1(new_n946), .B2(new_n940), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n943), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n930), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT106), .B1(new_n929), .B2(new_n930), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n900), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G8), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(G1976), .B2(new_n759), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n955), .B(new_n956), .C1(G1976), .C2(new_n759), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n575), .B(G1981), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT109), .B1(new_n959), .B2(KEYINPUT108), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT109), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n962), .B2(KEYINPUT49), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n960), .A2(KEYINPUT49), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n954), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n957), .A2(new_n958), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n942), .A2(new_n950), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n900), .A2(KEYINPUT45), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n953), .A2(KEYINPUT112), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n926), .A2(new_n931), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n971), .B(new_n900), .C1(new_n972), .C2(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n921), .A2(new_n894), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n733), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n923), .A2(new_n932), .A3(G2084), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT122), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(G168), .A2(new_n920), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT123), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n975), .B2(new_n733), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT122), .B1(new_n984), .B2(new_n920), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n981), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT51), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(KEYINPUT124), .A3(KEYINPUT51), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n984), .A2(new_n920), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n991), .A2(KEYINPUT51), .A3(new_n982), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n989), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n979), .A2(new_n982), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT121), .Z(new_n996));
  AND3_X1   g571(.A1(new_n994), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT125), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT62), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT125), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n986), .A2(KEYINPUT124), .A3(KEYINPUT51), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT124), .B1(new_n986), .B2(KEYINPUT51), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n992), .ZN(new_n1003));
  INV_X1    g578(.A(new_n996), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n994), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OR2_X1    g583(.A1(new_n938), .A2(G2078), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n1009), .A2(new_n1010), .B1(new_n724), .B2(new_n934), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(G2078), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n975), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n999), .A2(new_n1008), .A3(G171), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n944), .A2(new_n945), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT113), .B(G1956), .Z(new_n1019));
  AND2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT56), .B(G2072), .Z(new_n1021));
  NOR2_X1   g596(.A1(new_n938), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1017), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT57), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1024), .A2(KEYINPUT57), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n692), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(G299), .A2(new_n1024), .A3(KEYINPUT57), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n1020), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n935), .A2(G1348), .B1(G2067), .B2(new_n953), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n593), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n1020), .A2(new_n1029), .A3(new_n1022), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g612(.A1(new_n1034), .A2(KEYINPUT115), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1032), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1029), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT61), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1036), .C2(new_n1040), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT60), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1033), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n592), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n1048), .B2(new_n1034), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT61), .B(new_n1036), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1047), .A2(new_n1046), .A3(new_n593), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1045), .A2(new_n1050), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n938), .A2(G1996), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT58), .B(G1341), .Z(new_n1055));
  NAND2_X1  g630(.A1(new_n953), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n809), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT117), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1057), .B2(KEYINPUT117), .ZN(new_n1062));
  OR3_X1    g637(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT120), .B(new_n1039), .C1(new_n1053), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1051), .B(new_n1052), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1068), .A2(new_n1065), .A3(new_n1049), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1039), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(G171), .B(KEYINPUT54), .Z(new_n1072));
  NOR2_X1   g647(.A1(new_n895), .A2(new_n1013), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(G40), .A3(G160), .A4(new_n937), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1011), .B1(KEYINPUT126), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g650(.A(new_n1072), .B(new_n1075), .C1(KEYINPUT126), .C2(new_n1074), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1014), .B2(new_n1072), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1016), .A2(new_n1066), .A3(new_n1071), .A4(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n968), .B1(new_n1015), .B2(new_n1078), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n964), .A2(G1976), .A3(G288), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G305), .A2(G1981), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n965), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n967), .B(KEYINPUT110), .ZN(new_n1083));
  INV_X1    g658(.A(new_n968), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n984), .A2(new_n920), .A3(G286), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT63), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT63), .B1(new_n941), .B2(new_n918), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n942), .A2(new_n1085), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1083), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI221_X1 g664(.A(new_n1082), .B1(new_n942), .B2(new_n1083), .C1(new_n1086), .C2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n916), .B1(new_n1079), .B2(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n901), .A2(G1986), .A3(G290), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT48), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n914), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n781), .A2(new_n783), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n912), .A2(new_n1095), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n676), .A2(G2067), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n901), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(KEYINPUT46), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n902), .B(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n901), .B1(new_n909), .B2(new_n908), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1099), .B2(KEYINPUT46), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(new_n1104), .B(KEYINPUT47), .Z(new_n1105));
  NOR3_X1   g680(.A1(new_n1094), .A2(new_n1098), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1091), .A2(new_n1106), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g682(.A1(new_n891), .A2(new_n464), .ZN(new_n1109));
  NOR2_X1   g683(.A1(G401), .A2(G227), .ZN(new_n1110));
  NAND4_X1  g684(.A1(new_n846), .A2(new_n1109), .A3(new_n662), .A4(new_n1110), .ZN(G225));
  INV_X1    g685(.A(G225), .ZN(G308));
endmodule


