//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n562, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  OR2_X1    g031(.A1(new_n456), .A2(KEYINPUT66), .ZN(new_n457));
  AOI22_X1  g032(.A1(new_n456), .A2(KEYINPUT66), .B1(G567), .B2(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  AND3_X1   g037(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(new_n462), .B2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n461), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n461), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n474), .B1(new_n475), .B2(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT67), .B1(new_n476), .B2(new_n461), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  OAI21_X1  g054(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n473), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n472), .B1(new_n477), .B2(new_n483), .ZN(G160));
  INV_X1    g059(.A(KEYINPUT3), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n485), .B1(new_n467), .B2(KEYINPUT68), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n487));
  AOI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n461), .B1(new_n486), .B2(new_n487), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n489), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  OAI211_X1 g070(.A(G138), .B(new_n461), .C1(new_n478), .C2(new_n479), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT4), .A2(G138), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n461), .B(new_n499), .C1(new_n463), .C2(new_n464), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n503), .B1(new_n463), .B2(new_n464), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(G114), .B2(new_n461), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n501), .A2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  NAND2_X1  g086(.A1(G75), .A2(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT71), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n510), .A2(new_n515), .A3(G88), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(G50), .A3(G543), .ZN(new_n517));
  AND3_X1   g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT70), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT70), .B1(new_n516), .B2(new_n517), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n515), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G51), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n515), .A2(G89), .ZN(new_n528));
  AND2_X1   g103(.A1(G63), .A2(G651), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n510), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  XOR2_X1   g107(.A(KEYINPUT5), .B(G543), .Z(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  INV_X1    g109(.A(G77), .ZN(new_n535));
  INV_X1    g110(.A(G543), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n533), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n539), .B1(new_n535), .B2(new_n536), .C1(new_n533), .C2(new_n534), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(G651), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT73), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n538), .A2(new_n543), .A3(new_n540), .A4(G651), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n510), .A2(new_n515), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(G90), .A2(new_n546), .B1(new_n523), .B2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n542), .A2(new_n544), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  INV_X1    g124(.A(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n533), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n550), .B1(new_n553), .B2(KEYINPUT74), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(KEYINPUT74), .B2(new_n553), .ZN(new_n555));
  AOI22_X1  g130(.A1(G81), .A2(new_n546), .B1(new_n523), .B2(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT75), .ZN(G176));
  XOR2_X1   g136(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n562));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n533), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n568), .B2(new_n569), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n523), .A2(new_n574), .A3(G53), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT9), .B1(new_n522), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n575), .A2(new_n577), .B1(G91), .B2(new_n546), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n573), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n520), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n514), .B(KEYINPUT78), .C1(new_n518), .C2(new_n519), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n510), .A2(new_n515), .A3(G87), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n515), .A2(G49), .A3(G543), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  INV_X1    g163(.A(G48), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n545), .A2(new_n588), .B1(new_n522), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n510), .A2(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n550), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n550), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n599));
  AOI22_X1  g174(.A1(G85), .A2(new_n546), .B1(new_n523), .B2(G47), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(G290));
  AND3_X1   g176(.A1(new_n510), .A2(new_n515), .A3(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n523), .A2(KEYINPUT80), .ZN(new_n604));
  INV_X1    g179(.A(G54), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n522), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n533), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n604), .A2(new_n607), .B1(new_n610), .B2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G171), .B2(new_n613), .ZN(G284));
  OAI21_X1  g190(.A(new_n614), .B1(G171), .B2(new_n613), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(new_n578), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(new_n572), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n617), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n617), .B1(new_n619), .B2(G868), .ZN(G280));
  INV_X1    g196(.A(new_n612), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n557), .A2(new_n613), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n612), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n470), .A2(new_n475), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n488), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n461), .A2(G111), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n637));
  AND3_X1   g212(.A1(new_n490), .A2(new_n637), .A3(G123), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n490), .B2(G123), .ZN(new_n639));
  OAI221_X1 g214(.A(new_n634), .B1(new_n635), .B2(new_n636), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT82), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n641), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n633), .A2(new_n643), .A3(new_n645), .ZN(G156));
  XNOR2_X1  g221(.A(G2427), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2430), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT85), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n657), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n661), .ZN(new_n663));
  AND3_X1   g238(.A1(new_n662), .A2(G14), .A3(new_n663), .ZN(G401));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n632), .ZN(new_n672));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n668), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(new_n642), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(new_n687), .B(new_n686), .S(new_n679), .Z(new_n688));
  NOR2_X1   g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT87), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT88), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n691), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT89), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G229));
  NAND2_X1  g275(.A1(new_n490), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n488), .A2(G131), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n461), .A2(G107), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n701), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(G16), .A2(G24), .ZN(new_n710));
  INV_X1    g285(.A(G290), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G16), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n709), .B(new_n713), .C1(KEYINPUT90), .C2(KEYINPUT36), .ZN(new_n714));
  NOR2_X1   g289(.A1(G6), .A2(G16), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n594), .B2(G16), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT32), .ZN(new_n717));
  INV_X1    g292(.A(G1981), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(G166), .A2(G16), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G16), .B2(G22), .ZN(new_n721));
  INV_X1    g296(.A(G1971), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G16), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G23), .ZN(new_n726));
  INV_X1    g301(.A(G288), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT33), .B(G1976), .Z(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  NAND4_X1  g305(.A1(new_n719), .A2(new_n723), .A3(new_n724), .A4(new_n730), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT34), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n714), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT91), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n725), .A2(G19), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n558), .B2(new_n725), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1341), .Z(new_n740));
  INV_X1    g315(.A(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G26), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT28), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n490), .A2(G128), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n488), .A2(G140), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n461), .A2(G116), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT92), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n743), .B1(new_n749), .B2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2067), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n725), .A2(G4), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n622), .B2(new_n725), .ZN(new_n753));
  INV_X1    g328(.A(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n740), .A2(new_n751), .A3(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT93), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n741), .A2(G32), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n490), .A2(G129), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n488), .A2(G141), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT26), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n470), .A2(G105), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n759), .A2(new_n760), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n758), .B1(new_n765), .B2(new_n741), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT27), .ZN(new_n767));
  INV_X1    g342(.A(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G5), .A2(G16), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT96), .Z(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G301), .B2(new_n725), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n769), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n725), .A2(G21), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G168), .B2(new_n725), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT95), .Z(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n780), .A2(G1966), .B1(G29), .B2(new_n641), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT30), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n782), .A2(G28), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n741), .B1(new_n782), .B2(G28), .ZN(new_n784));
  AND2_X1   g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NOR2_X1   g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  OAI22_X1  g361(.A1(new_n783), .A2(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n741), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n741), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n787), .B1(new_n789), .B2(G2078), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n781), .B(new_n790), .C1(G2078), .C2(new_n789), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT25), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n475), .A2(G127), .ZN(new_n794));
  NAND2_X1  g369(.A1(G115), .A2(G2104), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n461), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI211_X1 g371(.A(new_n793), .B(new_n796), .C1(G139), .C2(new_n488), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT94), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n741), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n741), .B2(G33), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(G2072), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT98), .B(KEYINPUT23), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n725), .A2(G20), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  INV_X1    g383(.A(G2072), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n801), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G1966), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n779), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT24), .ZN(new_n813));
  INV_X1    g388(.A(G34), .ZN(new_n814));
  AOI21_X1  g389(.A(G29), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n813), .B2(new_n814), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G160), .B2(new_n741), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G2084), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n741), .A2(G35), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G162), .B2(new_n741), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G2090), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n817), .A2(G2084), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n812), .A2(new_n818), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n791), .A2(new_n803), .A3(new_n810), .A4(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n737), .A2(new_n757), .A3(new_n776), .A4(new_n826), .ZN(G150));
  INV_X1    g402(.A(G150), .ZN(G311));
  INV_X1    g403(.A(G93), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT100), .B(G55), .Z(new_n830));
  OAI22_X1  g405(.A1(new_n545), .A2(new_n829), .B1(new_n522), .B2(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(new_n550), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G860), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n557), .B1(new_n838), .B2(new_n834), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n834), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n557), .B(KEYINPUT101), .C1(new_n833), .C2(new_n831), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n612), .A2(new_n623), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n844));
  XOR2_X1   g419(.A(new_n843), .B(new_n844), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n842), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n835), .B1(new_n847), .B2(KEYINPUT39), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n837), .B1(new_n848), .B2(new_n849), .ZN(G145));
  XOR2_X1   g425(.A(new_n748), .B(KEYINPUT92), .Z(new_n851));
  AOI22_X1  g426(.A1(new_n488), .A2(new_n499), .B1(new_n496), .B2(new_n497), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n504), .A2(new_n853), .A3(new_n507), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n502), .B1(new_n486), .B2(new_n487), .ZN(new_n855));
  INV_X1    g430(.A(G114), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n505), .B1(new_n856), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT102), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n852), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n851), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n798), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n749), .B(new_n859), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(new_n799), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n764), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n630), .B(new_n705), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n488), .A2(G142), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n867), .B(KEYINPUT103), .Z(new_n868));
  NAND2_X1  g443(.A1(new_n490), .A2(G130), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT104), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n461), .A2(G118), .ZN(new_n871));
  OAI21_X1  g446(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n868), .B(new_n870), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n866), .B(new_n873), .Z(new_n874));
  NAND3_X1  g449(.A1(new_n861), .A2(new_n765), .A3(new_n863), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n865), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n874), .B1(new_n865), .B2(new_n875), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n865), .A2(KEYINPUT105), .A3(new_n874), .A4(new_n875), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n641), .B(new_n494), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G160), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n878), .A2(new_n880), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n876), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n883), .B1(new_n886), .B2(new_n879), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g465(.A(new_n842), .B(new_n626), .Z(new_n891));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(G299), .B2(new_n622), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n619), .A2(KEYINPUT106), .A3(new_n612), .ZN(new_n894));
  NAND2_X1  g469(.A1(G299), .A2(new_n622), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n891), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n842), .B(new_n626), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n900), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n893), .A2(new_n894), .A3(KEYINPUT41), .A4(new_n895), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(KEYINPUT107), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G290), .B(G166), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n594), .B(new_n727), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n909), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n897), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n910), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n910), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(G868), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g493(.A(new_n917), .B1(G868), .B2(new_n834), .ZN(G331));
  NAND2_X1  g494(.A1(G286), .A2(KEYINPUT109), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n921));
  NAND2_X1  g496(.A1(G168), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(G171), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(G301), .A2(KEYINPUT109), .A3(G286), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n842), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n840), .A2(new_n923), .A3(new_n841), .A4(new_n924), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(new_n901), .A3(new_n904), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(new_n896), .A3(new_n927), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n913), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n888), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n909), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT43), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n902), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n939));
  OR2_X1    g514(.A1(new_n903), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n896), .A2(KEYINPUT110), .A3(new_n900), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n903), .A2(new_n939), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n938), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n928), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n913), .B1(new_n944), .B2(new_n930), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n945), .A2(new_n932), .A3(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT44), .B1(new_n936), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n946), .B1(new_n933), .B2(new_n935), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n945), .A2(new_n932), .A3(KEYINPUT43), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n951), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g527(.A(G1384), .ZN(new_n953));
  OAI211_X1 g528(.A(KEYINPUT45), .B(new_n953), .C1(new_n501), .C2(new_n508), .ZN(new_n954));
  NAND3_X1  g529(.A1(G160), .A2(new_n954), .A3(G40), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT45), .B1(new_n859), .B2(new_n953), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n811), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G40), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n958), .B(new_n472), .C1(new_n477), .C2(new_n483), .ZN(new_n959));
  INV_X1    g534(.A(G2084), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n859), .A2(new_n961), .A3(new_n953), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n953), .B1(new_n501), .B2(new_n508), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT50), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n959), .A2(new_n960), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n957), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(G8), .A3(G286), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT120), .B(G8), .C1(new_n966), .C2(G286), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT121), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n969), .A3(KEYINPUT51), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT51), .ZN(new_n972));
  OAI21_X1  g547(.A(G8), .B1(new_n966), .B2(G286), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(new_n973), .B2(new_n969), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n967), .B(new_n970), .C1(new_n971), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1976), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(G288), .B2(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT115), .ZN(new_n978));
  NOR2_X1   g553(.A1(G288), .A2(new_n976), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT114), .ZN(new_n980));
  NAND4_X1  g555(.A1(G160), .A2(G40), .A3(new_n953), .A4(new_n859), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n978), .A2(new_n980), .A3(G8), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n477), .A2(new_n483), .ZN(new_n983));
  INV_X1    g558(.A(new_n472), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(G40), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n859), .A2(new_n953), .ZN(new_n986));
  OAI21_X1  g561(.A(G8), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT114), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n979), .B(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT49), .ZN(new_n991));
  OAI21_X1  g566(.A(G1981), .B1(new_n590), .B2(new_n593), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n590), .A2(new_n593), .A3(G1981), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n594), .A2(new_n718), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n992), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n995), .A2(new_n997), .A3(G8), .A4(new_n981), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n982), .A2(new_n990), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n581), .A2(G8), .A3(new_n582), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n581), .A2(KEYINPUT55), .A3(G8), .A4(new_n582), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n859), .A2(KEYINPUT45), .A3(new_n953), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n963), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n959), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n722), .ZN(new_n1009));
  INV_X1    g584(.A(G2090), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n959), .A2(new_n1010), .A3(new_n962), .A4(new_n964), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1004), .A2(new_n1012), .A3(G8), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(KEYINPUT116), .A3(new_n959), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n961), .B1(new_n859), .B2(new_n953), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1017), .B1(new_n1018), .B2(new_n985), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n855), .A2(new_n857), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n852), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n961), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1016), .A2(new_n1019), .A3(new_n1010), .A4(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1014), .B1(new_n1023), .B2(new_n1009), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n999), .B(new_n1013), .C1(new_n1024), .C2(new_n1004), .ZN(new_n1025));
  INV_X1    g600(.A(G2078), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n959), .A2(new_n1026), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n959), .A2(new_n962), .A3(new_n964), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n773), .ZN(new_n1031));
  INV_X1    g606(.A(new_n956), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(new_n959), .A3(new_n954), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1026), .A2(KEYINPUT53), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1029), .B(new_n1031), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G301), .A2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n542), .A2(KEYINPUT54), .A3(new_n544), .A4(new_n547), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1035), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n476), .A2(new_n461), .ZN(new_n1042));
  NOR4_X1   g617(.A1(new_n1042), .A2(new_n472), .A3(new_n958), .A4(new_n1034), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1032), .A2(new_n1005), .A3(new_n1043), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1039), .A2(new_n1029), .A3(new_n1031), .A4(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1041), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1025), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n975), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1016), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1049));
  INV_X1    g624(.A(G1956), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT56), .B(G2072), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n959), .A2(new_n1005), .A3(new_n1007), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n573), .A2(new_n1054), .A3(new_n578), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT57), .B1(new_n618), .B2(new_n572), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1051), .A2(new_n1053), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1018), .A2(new_n985), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1060), .A2(KEYINPUT116), .B1(new_n961), .B2(new_n1021), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1956), .B1(new_n1061), .B2(new_n1019), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1053), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1057), .B(KEYINPUT118), .ZN(new_n1065));
  OAI211_X1 g640(.A(KEYINPUT61), .B(new_n1059), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  AOI211_X1 g642(.A(new_n1063), .B(new_n1057), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1058), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G2067), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n959), .A2(new_n953), .A3(new_n1071), .A4(new_n859), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT117), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1030), .A2(new_n754), .ZN(new_n1074));
  INV_X1    g649(.A(new_n986), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n959), .A2(new_n1075), .A3(new_n1076), .A4(new_n1071), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1073), .A2(new_n1074), .A3(KEYINPUT60), .A4(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n612), .ZN(new_n1079));
  AOI22_X1  g654(.A1(KEYINPUT117), .A2(new_n1072), .B1(new_n1030), .B2(new_n754), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(KEYINPUT60), .A3(new_n622), .A4(new_n1077), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1073), .A2(new_n1074), .A3(new_n1077), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT60), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1079), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n1086));
  OR2_X1    g661(.A1(new_n1086), .A2(KEYINPUT59), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1088));
  NAND4_X1  g663(.A1(new_n959), .A2(new_n768), .A3(new_n1005), .A4(new_n1007), .ZN(new_n1089));
  XOR2_X1   g664(.A(KEYINPUT58), .B(G1341), .Z(new_n1090));
  NAND2_X1  g665(.A1(new_n981), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n557), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  MUX2_X1   g667(.A(new_n1087), .B(new_n1088), .S(new_n1092), .Z(new_n1093));
  NAND4_X1  g668(.A1(new_n1066), .A2(new_n1070), .A3(new_n1085), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1082), .A2(new_n622), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1064), .A2(new_n1065), .B1(new_n1068), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1048), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n966), .A2(G8), .A3(G168), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1099), .B1(new_n1025), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1012), .A2(G8), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1100), .A2(new_n1099), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n1013), .A4(new_n999), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n982), .A2(new_n990), .A3(new_n998), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1013), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n998), .A2(new_n976), .A3(new_n727), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n987), .B1(new_n1109), .B2(new_n996), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n1098), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1111), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1093), .A2(new_n1085), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1057), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT61), .B1(new_n1118), .B2(new_n1059), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1096), .B1(new_n1120), .B2(new_n1066), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1114), .B(new_n1116), .C1(new_n1121), .C2(new_n1048), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  INV_X1    g698(.A(new_n975), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n975), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1035), .A2(G171), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1025), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1126), .A2(new_n1127), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1113), .A2(new_n1122), .A3(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n749), .B(new_n1071), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1032), .A2(new_n985), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1136), .A2(KEYINPUT113), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(KEYINPUT113), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n764), .B(G1996), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1137), .A2(new_n1138), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n705), .A2(new_n708), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n705), .A2(new_n708), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1134), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1140), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(G1986), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n711), .A2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT112), .Z(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n1145), .B2(new_n711), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1144), .B1(new_n1134), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1132), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1134), .A2(new_n768), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT46), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT125), .Z(new_n1155));
  AOI21_X1  g730(.A(new_n1135), .B1(new_n1133), .B2(new_n765), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1147), .A2(new_n1134), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT48), .Z(new_n1162));
  OAI21_X1  g737(.A(new_n1160), .B1(new_n1144), .B2(new_n1162), .ZN(new_n1163));
  AOI22_X1  g738(.A1(new_n1140), .A2(new_n1142), .B1(new_n1071), .B2(new_n851), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1135), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1151), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g744(.A1(new_n459), .A2(G227), .ZN(new_n1171));
  XNOR2_X1  g745(.A(new_n1171), .B(KEYINPUT127), .ZN(new_n1172));
  NOR2_X1   g746(.A1(G401), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n699), .A2(new_n889), .A3(new_n1173), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n1174), .A2(new_n951), .ZN(G308));
  OR2_X1    g749(.A1(new_n1174), .A2(new_n951), .ZN(G225));
endmodule


