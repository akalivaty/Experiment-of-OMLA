//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1178, new_n1179,
    new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n452), .A2(G567), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT65), .Z(new_n456));
  AOI21_X1  g031(.A(new_n456), .B1(new_n451), .B2(G2106), .ZN(G319));
  INV_X1    g032(.A(G125), .ZN(new_n458));
  OR2_X1    g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G113), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(KEYINPUT67), .B(G2105), .C1(new_n461), .C2(new_n466), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT68), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n472), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n475), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n480), .C2(new_n481), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n491), .A2(new_n493), .A3(G2104), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n497), .B1(new_n480), .B2(new_n481), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n497), .B(new_n500), .C1(new_n481), .C2(new_n480), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n495), .B1(new_n499), .B2(new_n501), .ZN(G164));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT71), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(G543), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n506), .A2(KEYINPUT71), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n505), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  OAI211_X1 g088(.A(G50), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n517), .A2(KEYINPUT69), .A3(G50), .A4(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n513), .A2(G88), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n510), .B2(new_n512), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(G651), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT72), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(G166));
  NAND2_X1  g104(.A1(new_n510), .A2(new_n512), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n510), .A2(new_n532), .A3(new_n512), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g109(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n513), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n505), .A2(new_n511), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G51), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n535), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n534), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G651), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n513), .A2(G90), .B1(new_n539), .B2(G52), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n531), .B2(new_n533), .ZN(new_n550));
  AND2_X1   g125(.A1(G68), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT74), .B(G43), .Z(new_n553));
  AOI22_X1  g128(.A1(new_n513), .A2(G81), .B1(new_n539), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND3_X1  g137(.A1(new_n539), .A2(KEYINPUT76), .A3(G53), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n564), .A2(new_n565), .B1(G91), .B2(new_n513), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n530), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n544), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT72), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT72), .B1(new_n519), .B2(new_n524), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT77), .ZN(new_n576));
  AND2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G303));
  AOI22_X1  g152(.A1(new_n513), .A2(G87), .B1(new_n539), .B2(G49), .ZN(new_n578));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n531), .A2(new_n579), .A3(new_n533), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n580), .A2(new_n581), .A3(G651), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n581), .B1(new_n580), .B2(G651), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(G288));
  AOI22_X1  g160(.A1(new_n513), .A2(G86), .B1(new_n539), .B2(G48), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n510), .B2(new_n512), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n591), .A2(new_n592), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n586), .B1(new_n593), .B2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n534), .A2(G60), .ZN(new_n596));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n544), .B1(new_n598), .B2(KEYINPUT80), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(KEYINPUT80), .B2(new_n598), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n513), .A2(G85), .B1(new_n539), .B2(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n600), .A2(KEYINPUT81), .A3(new_n601), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(new_n513), .A2(G92), .ZN(new_n607));
  XOR2_X1   g182(.A(new_n607), .B(KEYINPUT10), .Z(new_n608));
  NAND2_X1  g183(.A1(new_n530), .A2(G66), .ZN(new_n609));
  INV_X1    g184(.A(G79), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n511), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n539), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(G171), .B2(new_n614), .ZN(G321));
  NAND2_X1  g192(.A1(G299), .A2(new_n614), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(new_n614), .B2(G168), .ZN(G297));
  OAI21_X1  g194(.A(new_n618), .B1(new_n614), .B2(G168), .ZN(G280));
  INV_X1    g195(.A(G860), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n613), .B1(G559), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g198(.A1(new_n555), .A2(new_n614), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n613), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g202(.A(KEYINPUT3), .B(G2104), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n472), .A2(G2104), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT83), .B(G2100), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n483), .A2(G123), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n475), .A2(G135), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n472), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(G2096), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n634), .A2(new_n635), .A3(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n653), .A2(new_n656), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(G401));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n664), .B2(new_n661), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n665), .B1(KEYINPUT85), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(KEYINPUT85), .B2(new_n667), .ZN(new_n669));
  INV_X1    g244(.A(new_n661), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n670), .A2(new_n666), .A3(new_n663), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n662), .A2(new_n666), .A3(new_n664), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(new_n641), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT86), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1971), .B(G1976), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n682), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  AOI211_X1 g261(.A(new_n684), .B(new_n686), .C1(new_n679), .C2(new_n683), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1981), .B(G1986), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT87), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n689), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G6), .ZN(new_n696));
  INV_X1    g271(.A(G305), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT32), .B(G1981), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n695), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(new_n578), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n580), .A2(G651), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(KEYINPUT78), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n703), .B1(new_n705), .B2(new_n582), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n702), .B1(new_n706), .B2(new_n695), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT90), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G16), .A2(G22), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G166), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1971), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n701), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n716));
  INV_X1    g291(.A(G290), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G16), .B2(G24), .ZN(new_n719));
  INV_X1    g294(.A(G1986), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n720), .B2(new_n719), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n715), .A2(KEYINPUT34), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT88), .B(G29), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G25), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n483), .A2(G119), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n475), .A2(G131), .ZN(new_n728));
  OR2_X1    g303(.A1(G95), .A2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n729), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n726), .B1(new_n732), .B2(new_n725), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT35), .B(G1991), .Z(new_n734));
  XOR2_X1   g309(.A(new_n733), .B(new_n734), .Z(new_n735));
  NOR3_X1   g310(.A1(new_n722), .A2(new_n723), .A3(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT36), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n695), .A2(G4), .ZN(new_n738));
  INV_X1    g313(.A(new_n613), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n695), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n695), .A2(G19), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n556), .B2(new_n695), .ZN(new_n744));
  INV_X1    g319(.A(G1341), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n724), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n483), .A2(G128), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n475), .A2(G140), .ZN(new_n750));
  OR2_X1    g325(.A1(G104), .A2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n753), .A2(KEYINPUT91), .A3(G29), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT91), .B1(new_n753), .B2(G29), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n748), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n742), .A2(new_n746), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(KEYINPUT92), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(KEYINPUT92), .ZN(new_n761));
  INV_X1    g336(.A(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G32), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT26), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n475), .A2(G141), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n629), .A2(G105), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n765), .B(new_n768), .C1(G129), .C2(new_n483), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n763), .B1(new_n769), .B2(new_n762), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT27), .B(G1996), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G162), .A2(new_n725), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G35), .B2(new_n725), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT29), .B(G2090), .Z(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n724), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n724), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2078), .ZN(new_n779));
  INV_X1    g354(.A(G28), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(KEYINPUT30), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(KEYINPUT30), .B2(new_n780), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT95), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n782), .B(new_n784), .C1(new_n640), .C2(new_n724), .ZN(new_n785));
  OR3_X1    g360(.A1(new_n776), .A2(new_n779), .A3(new_n785), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n772), .B(new_n786), .C1(new_n774), .C2(new_n775), .ZN(new_n787));
  NOR2_X1   g362(.A1(G168), .A2(new_n695), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n695), .B2(G21), .ZN(new_n789));
  INV_X1    g364(.A(G1966), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT25), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n475), .A2(G139), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT93), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n472), .B2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G33), .B(new_n799), .S(G29), .Z(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G2072), .ZN(new_n801));
  INV_X1    g376(.A(G2084), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT24), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(G34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(G34), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n724), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n478), .B2(new_n762), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n801), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n789), .A2(new_n790), .B1(new_n800), .B2(G2072), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n787), .A2(new_n791), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n695), .A2(G20), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT23), .Z(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G299), .B2(G16), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1956), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n807), .A2(new_n802), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(KEYINPUT94), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n815), .A2(KEYINPUT94), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n695), .A2(G5), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(G171), .B2(new_n695), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1961), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n810), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n737), .A2(new_n760), .A3(new_n761), .A4(new_n822), .ZN(G150));
  INV_X1    g398(.A(G150), .ZN(G311));
  NAND2_X1  g399(.A1(new_n739), .A2(G559), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n534), .A2(G67), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n544), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n513), .A2(G93), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n539), .A2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n556), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n555), .B1(new_n829), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n826), .B(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n621), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n833), .A2(new_n621), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n478), .B(new_n640), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n488), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n753), .B(G164), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n799), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n769), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n483), .A2(G130), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n472), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G142), .B2(new_n475), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(new_n631), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n731), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n850), .A2(new_n857), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n847), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT96), .Z(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n858), .B(new_n847), .C1(KEYINPUT97), .C2(new_n859), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n859), .A2(KEYINPUT97), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g442(.A(new_n613), .B(G299), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n868), .B(KEYINPUT41), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n836), .B(new_n625), .ZN(new_n871));
  MUX2_X1   g446(.A(new_n869), .B(new_n870), .S(new_n871), .Z(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT42), .Z(new_n873));
  XNOR2_X1  g448(.A(G288), .B(G166), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n876));
  NOR2_X1   g451(.A1(G290), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(G290), .A2(new_n876), .ZN(new_n879));
  AOI21_X1  g454(.A(G305), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n879), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n881), .A2(new_n697), .A3(new_n877), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n875), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n697), .B1(new_n881), .B2(new_n877), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n878), .A2(G305), .A3(new_n879), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n874), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n883), .A2(KEYINPUT99), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n873), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(G868), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(G868), .B2(new_n833), .ZN(G295));
  OAI21_X1  g465(.A(new_n889), .B1(G868), .B2(new_n833), .ZN(G331));
  NAND2_X1  g466(.A1(G301), .A2(G168), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT100), .Z(new_n893));
  NOR2_X1   g468(.A1(G301), .A2(G168), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT101), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n836), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n836), .B1(new_n893), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n870), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n869), .A3(new_n896), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(new_n883), .A3(new_n886), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(new_n862), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n902), .B1(new_n886), .B2(new_n883), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n883), .A2(new_n886), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(new_n899), .A3(new_n901), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n908), .A2(new_n909), .A3(new_n862), .A4(new_n903), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n911), .B(new_n912), .ZN(G397));
  INV_X1    g488(.A(KEYINPUT126), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n474), .A2(G40), .A3(new_n476), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n463), .B(new_n465), .C1(new_n482), .C2(new_n458), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT67), .B1(new_n916), .B2(G2105), .ZN(new_n917));
  INV_X1    g492(.A(new_n470), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G164), .B2(G1384), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR2_X1   g498(.A1(G290), .A2(G1986), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n769), .B(G1996), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n753), .B(new_n757), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n731), .B(new_n734), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT102), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n924), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G290), .A2(G1986), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G8), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT103), .B1(G164), .B2(G1384), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT103), .ZN(new_n936));
  INV_X1    g511(.A(G1384), .ZN(new_n937));
  INV_X1    g512(.A(new_n501), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n500), .B1(new_n628), .B2(new_n497), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n936), .B(new_n937), .C1(new_n940), .C2(new_n495), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n934), .A2(new_n935), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n474), .A2(new_n476), .A3(G40), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n943), .B1(new_n469), .B2(new_n470), .ZN(new_n944));
  NOR2_X1   g519(.A1(G164), .A2(G1384), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n935), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G2090), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n499), .A2(new_n501), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n490), .A2(new_n494), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n952), .A2(KEYINPUT45), .A3(new_n937), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n921), .A2(new_n944), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n713), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n933), .B1(new_n949), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT55), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n933), .B1(KEYINPUT104), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n575), .A2(new_n576), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n957), .A2(KEYINPUT104), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n962));
  INV_X1    g537(.A(new_n960), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n575), .A2(new_n576), .A3(new_n958), .A4(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n962), .B1(new_n961), .B2(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n956), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n934), .A2(new_n944), .A3(new_n941), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G8), .ZN(new_n969));
  INV_X1    g544(.A(G1981), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(new_n586), .C1(new_n593), .C2(new_n594), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(new_n586), .B2(new_n591), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(KEYINPUT106), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n974), .B(new_n970), .C1(new_n586), .C2(new_n591), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n971), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT49), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n972), .B(KEYINPUT106), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n982), .A2(KEYINPUT107), .A3(new_n977), .A4(new_n971), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n969), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n969), .B1(G1976), .B2(new_n706), .ZN(new_n985));
  INV_X1    g560(.A(G1976), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(G288), .B2(new_n986), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n968), .A2(G8), .ZN(new_n990));
  OAI211_X1 g565(.A(G1976), .B(new_n578), .C1(new_n583), .C2(new_n584), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n984), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n961), .A2(new_n964), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n936), .B1(new_n952), .B2(new_n937), .ZN(new_n995));
  AOI211_X1 g570(.A(KEYINPUT103), .B(G1384), .C1(new_n950), .C2(new_n951), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT109), .B(new_n944), .C1(new_n997), .C2(new_n935), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n935), .B1(new_n934), .B2(new_n941), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n999), .B1(new_n1000), .B2(new_n919), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n945), .A2(new_n935), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n998), .A2(new_n1001), .A3(new_n948), .A4(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(new_n955), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n994), .B1(new_n1004), .B2(new_n933), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n967), .A2(new_n993), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT121), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n934), .A2(new_n941), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n919), .B1(new_n1009), .B2(new_n920), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n953), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n952), .A2(KEYINPUT110), .A3(KEYINPUT45), .A4(new_n937), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G1966), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n934), .A2(new_n935), .A3(new_n941), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n944), .A3(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1018), .A2(G2084), .ZN(new_n1019));
  OAI21_X1  g594(.A(G8), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1008), .B1(new_n1020), .B2(KEYINPUT117), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n920), .B1(new_n995), .B2(new_n996), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n1022), .A3(new_n944), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n790), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n947), .A2(new_n802), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(G168), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G8), .ZN(new_n1027));
  OR2_X1    g602(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT62), .ZN(new_n1029));
  OAI21_X1  g604(.A(G286), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(new_n1026), .A3(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1021), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1028), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT121), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n967), .A2(new_n993), .A3(new_n1005), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G2078), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1014), .A2(new_n1022), .A3(new_n944), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1961), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n942), .B2(new_n946), .ZN(new_n1040));
  INV_X1    g615(.A(G2078), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n921), .A2(new_n944), .A3(new_n953), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1036), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1038), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G171), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1044), .A2(KEYINPUT118), .A3(G171), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1007), .A2(new_n1033), .A3(new_n1035), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT123), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n1021), .A2(new_n1031), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT62), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1050), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(KEYINPUT123), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  OAI211_X1 g637(.A(G8), .B(G168), .C1(new_n1015), .C2(new_n1019), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1062), .B1(new_n1006), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n956), .B1(new_n961), .B2(new_n964), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1065), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n967), .A3(new_n993), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n706), .A2(new_n986), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n981), .A2(new_n983), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n971), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(new_n990), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n981), .A2(new_n983), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n990), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n992), .B1(new_n985), .B2(new_n987), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n967), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT108), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT108), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1079), .B(new_n1072), .C1(new_n967), .C2(new_n1076), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1064), .A2(new_n1067), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1018), .A2(new_n1039), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1082));
  AOI211_X1 g657(.A(new_n1046), .B(G301), .C1(new_n1082), .C2(new_n1038), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT118), .B1(new_n1044), .B2(G171), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n943), .B1(G2105), .B2(new_n916), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n921), .A2(new_n1085), .A3(KEYINPUT119), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT119), .B1(new_n921), .B2(new_n1085), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n953), .B(new_n1037), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1082), .A2(G301), .A3(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1083), .A2(new_n1084), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT120), .B1(new_n1091), .B2(KEYINPUT54), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT54), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1093), .B(new_n1094), .C1(new_n1049), .C2(new_n1090), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT54), .B1(new_n1044), .B2(G171), .ZN(new_n1097));
  AOI21_X1  g672(.A(G301), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1096), .A2(new_n1007), .A3(new_n1035), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT116), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT56), .B(G2072), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT112), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n954), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1107));
  INV_X1    g682(.A(G1956), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT57), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(KEYINPUT111), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G299), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(KEYINPUT111), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1103), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1102), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1116), .B2(new_n1115), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT115), .B1(new_n1119), .B2(KEYINPUT114), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(KEYINPUT115), .B2(new_n1119), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(new_n745), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n968), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1996), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n921), .A2(new_n944), .A3(new_n953), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n555), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  MUX2_X1   g702(.A(new_n1120), .B(new_n1121), .S(new_n1127), .Z(new_n1128));
  NOR2_X1   g703(.A1(new_n968), .A2(G2067), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n741), .B2(new_n1018), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(KEYINPUT60), .A3(new_n739), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(KEYINPUT60), .B2(new_n1130), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n739), .B1(new_n1130), .B2(KEYINPUT60), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1128), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1109), .A2(new_n1114), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n1116), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1136), .B2(new_n1102), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n613), .B2(new_n1130), .ZN(new_n1138));
  AOI22_X1  g713(.A1(new_n1118), .A2(new_n1137), .B1(new_n1116), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1081), .B1(new_n1101), .B2(new_n1139), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1052), .A2(new_n1061), .B1(new_n1140), .B2(KEYINPUT122), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1081), .B(new_n1142), .C1(new_n1101), .C2(new_n1139), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n932), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n929), .A2(new_n927), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(new_n923), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n924), .A2(new_n922), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1148), .B2(KEYINPUT48), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(KEYINPUT48), .B2(new_n1148), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n732), .A2(new_n734), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n927), .A2(new_n1151), .B1(G2067), .B2(new_n753), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n922), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n1125), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT46), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n926), .A2(new_n769), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n923), .B2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT125), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT47), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1150), .A2(new_n1153), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n914), .B1(new_n1144), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1140), .A2(KEYINPUT122), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1060), .A2(KEYINPUT123), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1059), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1163), .A2(new_n1052), .A3(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1162), .A2(new_n1165), .A3(new_n1143), .ZN(new_n1166));
  INV_X1    g741(.A(new_n932), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1160), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT126), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1161), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g745(.A1(G229), .A2(G227), .ZN(new_n1172));
  OAI211_X1 g746(.A(new_n1172), .B(G319), .C1(new_n659), .C2(new_n658), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n866), .A2(new_n1173), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n911), .A2(KEYINPUT127), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g749(.A(KEYINPUT127), .B1(new_n911), .B2(new_n1174), .ZN(new_n1176));
  NOR2_X1   g750(.A1(new_n1175), .A2(new_n1176), .ZN(G308));
  NAND2_X1  g751(.A1(new_n911), .A2(new_n1174), .ZN(new_n1178));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n1179));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n911), .A2(new_n1174), .A3(KEYINPUT127), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1181), .ZN(G225));
endmodule


