//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:54 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(G952), .ZN(new_n187));
  AOI211_X1 g001(.A(G953), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT68), .A2(G953), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT68), .A2(G953), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G902), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n193), .B1(G234), .B2(G237), .ZN(new_n194));
  AND2_X1   g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT21), .B(G898), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n188), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G214), .B1(G237), .B2(G902), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT67), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n200));
  INV_X1    g014(.A(G113), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(KEYINPUT66), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n203), .B1(KEYINPUT2), .B2(G113), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT2), .A2(G113), .ZN(new_n206));
  XNOR2_X1  g020(.A(G116), .B(G119), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n205), .B2(new_n206), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n199), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  NOR3_X1   g024(.A1(new_n203), .A2(KEYINPUT2), .A3(G113), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT66), .B1(new_n200), .B2(new_n201), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n206), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n207), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(KEYINPUT67), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT4), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT77), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n220), .A2(KEYINPUT3), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n221), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(G107), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT77), .ZN(new_n228));
  INV_X1    g042(.A(G107), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G104), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n219), .B(G101), .C1(new_n225), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(G101), .B1(new_n225), .B2(new_n231), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n227), .A2(KEYINPUT77), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n228), .B1(new_n234), .B2(new_n230), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n221), .A2(new_n223), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n226), .A4(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n218), .A2(new_n232), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  OAI21_X1  g057(.A(G113), .B1(new_n243), .B2(KEYINPUT5), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n244), .B1(KEYINPUT5), .B2(new_n207), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n208), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT79), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n230), .A2(new_n226), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G101), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n238), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n238), .B2(new_n249), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n240), .A2(new_n241), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT6), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n241), .B1(new_n240), .B2(new_n252), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT84), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n240), .A2(new_n252), .ZN(new_n257));
  INV_X1    g071(.A(new_n241), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT6), .A4(new_n253), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G143), .B(G146), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT0), .B(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT85), .ZN(new_n272));
  INV_X1    g086(.A(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(KEYINPUT1), .ZN(new_n274));
  AND3_X1   g088(.A1(new_n274), .A2(new_n263), .A3(new_n265), .ZN(new_n275));
  OR2_X1    g089(.A1(KEYINPUT65), .A2(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT65), .A2(G128), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT1), .B1(new_n264), .B2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n268), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n272), .B1(new_n283), .B2(G125), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n271), .A2(KEYINPUT85), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G224), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G953), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n286), .B(new_n288), .Z(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n255), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n256), .A2(new_n261), .A3(new_n289), .A4(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G210), .B1(G237), .B2(G902), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT7), .B1(new_n287), .B2(G953), .ZN(new_n294));
  OR3_X1    g108(.A1(new_n284), .A2(new_n285), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n284), .B2(new_n285), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n295), .A2(new_n253), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n241), .B(KEYINPUT8), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n252), .A2(KEYINPUT86), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n238), .A2(new_n249), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n208), .B2(new_n245), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n301), .B1(new_n252), .B2(KEYINPUT86), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n298), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(G902), .B1(new_n297), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n292), .A2(new_n293), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n293), .B1(new_n292), .B2(new_n304), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n198), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n198), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n292), .A2(new_n304), .ZN(new_n312));
  INV_X1    g126(.A(new_n293), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n314), .B2(new_n305), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT87), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n197), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G113), .B(G122), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(new_n222), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G125), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G140), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(new_n262), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT68), .A2(G953), .ZN(new_n326));
  INV_X1    g140(.A(G237), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT68), .A2(G953), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n326), .A2(G214), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n264), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n191), .A2(G143), .A3(G214), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g146(.A1(KEYINPUT18), .A2(G131), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n325), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n332), .A2(new_n333), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G131), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n330), .A2(new_n331), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n338), .B1(new_n330), .B2(new_n331), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n321), .A2(new_n323), .A3(KEYINPUT16), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n262), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(G146), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(KEYINPUT72), .A3(new_n348), .ZN(new_n349));
  AOI211_X1 g163(.A(KEYINPUT72), .B(G146), .C1(new_n344), .C2(new_n345), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n349), .A2(new_n351), .B1(new_n340), .B2(KEYINPUT17), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n343), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n332), .A2(KEYINPUT17), .A3(G131), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(KEYINPUT72), .ZN(new_n356));
  AOI21_X1  g170(.A(G146), .B1(new_n344), .B2(new_n345), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n355), .B(new_n353), .C1(new_n358), .C2(new_n350), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n319), .B(new_n337), .C1(new_n354), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n355), .B1(new_n358), .B2(new_n350), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n363), .A2(KEYINPUT88), .B1(new_n342), .B2(new_n341), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n336), .B1(new_n364), .B2(new_n359), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT90), .B1(new_n365), .B2(new_n319), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n337), .B1(new_n354), .B2(new_n360), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT90), .ZN(new_n368));
  INV_X1    g182(.A(new_n319), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n362), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(G475), .B1(new_n371), .B2(G902), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n346), .A2(new_n262), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n324), .B(KEYINPUT19), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n373), .B(new_n341), .C1(new_n262), .C2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n369), .B1(new_n375), .B2(new_n336), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n361), .ZN(new_n377));
  NOR2_X1   g191(.A1(G475), .A2(G902), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(KEYINPUT89), .A3(new_n361), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n383), .A2(KEYINPUT20), .A3(new_n378), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n372), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT9), .B(G234), .ZN(new_n387));
  INV_X1    g201(.A(G217), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n387), .A2(new_n388), .A3(G953), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n391));
  INV_X1    g205(.A(G122), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(G116), .ZN(new_n393));
  INV_X1    g207(.A(G116), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(KEYINPUT91), .A3(G122), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n396), .A2(KEYINPUT14), .B1(G116), .B2(new_n392), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n397), .A2(KEYINPUT93), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n396), .A2(KEYINPUT14), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n397), .B2(KEYINPUT93), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n229), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n276), .A2(G143), .A3(new_n277), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n273), .A2(G143), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(G134), .ZN(new_n406));
  INV_X1    g220(.A(G134), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n402), .B2(new_n404), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n392), .A2(G116), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(new_n409), .ZN(new_n410));
  OAI22_X1  g224(.A1(new_n406), .A2(new_n408), .B1(G107), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n407), .B1(new_n413), .B2(new_n403), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n405), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(G134), .B2(new_n405), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n410), .B(new_n229), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n390), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  OAI221_X1 g233(.A(new_n389), .B1(new_n417), .B2(new_n416), .C1(new_n401), .C2(new_n411), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(G478), .B1(KEYINPUT94), .B2(KEYINPUT15), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(KEYINPUT94), .B2(KEYINPUT15), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n421), .A2(new_n424), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n386), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G221), .B1(new_n387), .B2(G902), .ZN(new_n430));
  NAND2_X1  g244(.A1(KEYINPUT80), .A2(KEYINPUT12), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT12), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n300), .A2(KEYINPUT79), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n238), .A2(new_n247), .A3(new_n249), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n282), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n279), .A2(KEYINPUT78), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT78), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n263), .A2(new_n438), .A3(KEYINPUT1), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(G128), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n275), .B1(new_n440), .B2(new_n281), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n441), .A2(new_n300), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT64), .ZN(new_n444));
  INV_X1    g258(.A(G137), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT64), .A2(G137), .ZN(new_n447));
  AND2_X1   g261(.A1(KEYINPUT11), .A2(G134), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(KEYINPUT11), .A2(G134), .ZN(new_n450));
  NOR2_X1   g264(.A1(KEYINPUT11), .A2(G134), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(G137), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G131), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n452), .A3(new_n338), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT80), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n433), .B1(new_n443), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n433), .ZN(new_n461));
  AOI211_X1 g275(.A(new_n461), .B(new_n458), .C1(new_n436), .C2(new_n442), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT10), .B(new_n283), .C1(new_n250), .C2(new_n251), .ZN(new_n464));
  INV_X1    g278(.A(new_n456), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT10), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n441), .B2(new_n300), .ZN(new_n467));
  INV_X1    g281(.A(new_n270), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n239), .A2(new_n468), .A3(new_n232), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n464), .A2(new_n465), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n191), .A2(G227), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G140), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n463), .A2(KEYINPUT82), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT82), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n250), .A2(new_n251), .A3(new_n283), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n441), .A2(new_n300), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n459), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n461), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n443), .A2(new_n433), .A3(new_n459), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n476), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n478), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n469), .A2(new_n467), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT10), .B1(new_n488), .B2(new_n275), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n489), .B1(new_n434), .B2(new_n435), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n456), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n470), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n493));
  INV_X1    g307(.A(new_n475), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n497));
  OAI22_X1  g311(.A1(new_n477), .A2(new_n486), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G469), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n193), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n485), .A2(new_n491), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n487), .A2(new_n490), .A3(new_n456), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n502), .B1(new_n482), .B2(new_n483), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n503), .B2(new_n475), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT81), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT81), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n501), .B(new_n506), .C1(new_n503), .C2(new_n475), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(G469), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n499), .A2(new_n193), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n500), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n429), .A2(new_n430), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n317), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n446), .A2(new_n407), .A3(new_n447), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n338), .B1(G134), .B2(G137), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n455), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n282), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n270), .B1(new_n454), .B2(new_n455), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n514), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n455), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n338), .B1(new_n449), .B2(new_n452), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n468), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n455), .B(new_n517), .C1(new_n488), .C2(new_n275), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(KEYINPUT30), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n521), .A2(new_n218), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n524), .A2(new_n210), .A3(new_n217), .A4(new_n525), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT31), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n326), .A2(G210), .A3(new_n327), .A4(new_n328), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT27), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT27), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n191), .A2(new_n533), .A3(G210), .A4(new_n327), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT26), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n532), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n236), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n532), .A2(new_n534), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT26), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(G101), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n529), .A2(new_n530), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n527), .A2(new_n528), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT31), .B1(new_n546), .B2(new_n543), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT28), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n528), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n524), .A2(new_n525), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n551), .A2(new_n218), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n548), .B1(new_n552), .B2(KEYINPUT69), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n218), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n528), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n550), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n545), .B(new_n547), .C1(new_n557), .C2(new_n544), .ZN(new_n558));
  NOR2_X1   g372(.A1(G472), .A2(G902), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT32), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT71), .ZN(new_n563));
  INV_X1    g377(.A(G472), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n544), .A2(new_n549), .A3(KEYINPUT29), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n548), .B1(new_n554), .B2(new_n528), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n193), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT29), .B1(new_n546), .B2(new_n543), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n543), .B1(new_n548), .B2(new_n528), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n554), .A2(new_n555), .A3(new_n528), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT28), .B1(new_n554), .B2(new_n555), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n567), .B1(new_n573), .B2(KEYINPUT70), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT70), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n568), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  AOI211_X1 g390(.A(new_n563), .B(new_n564), .C1(new_n574), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n573), .A2(KEYINPUT70), .ZN(new_n578));
  INV_X1    g392(.A(new_n567), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT71), .B1(new_n580), .B2(G472), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n562), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n583));
  XOR2_X1   g397(.A(new_n583), .B(KEYINPUT22), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G137), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n242), .A2(G128), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT23), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n242), .B2(G128), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n276), .A2(G119), .A3(new_n277), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n587), .B(new_n589), .C1(new_n590), .C2(new_n588), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n590), .A2(new_n587), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT24), .B(G110), .Z(new_n593));
  AOI22_X1  g407(.A1(G110), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n351), .A3(new_n349), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n591), .A2(G110), .B1(new_n592), .B2(new_n593), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n324), .A2(new_n262), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n348), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT73), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT73), .B1(new_n595), .B2(new_n598), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n586), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n585), .B1(new_n599), .B2(new_n600), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n193), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT25), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT25), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n603), .A2(new_n607), .A3(new_n193), .A4(new_n604), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n388), .B1(G234), .B2(new_n193), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n606), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n603), .A2(new_n604), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n609), .A2(G902), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n610), .A2(KEYINPUT74), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(KEYINPUT74), .B1(new_n610), .B2(new_n613), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n582), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n513), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  INV_X1    g433(.A(new_n430), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT82), .B1(new_n463), .B2(new_n476), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n484), .A2(new_n485), .A3(new_n478), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n492), .A2(new_n494), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n495), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n509), .B1(new_n627), .B2(new_n499), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n620), .B1(new_n628), .B2(new_n508), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n558), .A2(new_n193), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n630), .A2(G472), .B1(new_n558), .B2(new_n559), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n629), .A2(new_n616), .A3(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n197), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n315), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n420), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n420), .A2(new_n635), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(KEYINPUT33), .A3(new_n419), .A4(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n193), .A2(G478), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT33), .B1(new_n419), .B2(new_n420), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(KEYINPUT95), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT95), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n642), .B(KEYINPUT33), .C1(new_n419), .C2(new_n420), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n638), .B(new_n639), .C1(new_n641), .C2(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n421), .A2(G478), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n386), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n634), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n632), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT97), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT34), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G104), .ZN(G6));
  NAND2_X1  g466(.A1(new_n383), .A2(new_n384), .ZN(new_n653));
  INV_X1    g467(.A(new_n378), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n380), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(new_n428), .A3(new_n372), .A4(new_n385), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n634), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n632), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR2_X1   g474(.A1(new_n585), .A2(KEYINPUT36), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n599), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n612), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n610), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n631), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n513), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n629), .A2(new_n582), .A3(new_n315), .A4(new_n664), .ZN(new_n670));
  INV_X1    g484(.A(new_n188), .ZN(new_n671));
  INV_X1    g485(.A(new_n195), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n671), .B1(new_n672), .B2(G900), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT98), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n656), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n669), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n582), .A2(new_n664), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n511), .A2(new_n315), .A3(new_n430), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n675), .A4(KEYINPUT99), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  OAI21_X1  g496(.A(KEYINPUT100), .B1(new_n306), .B2(new_n307), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT100), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n314), .A2(new_n684), .A3(new_n305), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n683), .A2(KEYINPUT38), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT38), .B1(new_n683), .B2(new_n685), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n386), .A2(new_n428), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n610), .A2(new_n663), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n529), .A2(new_n543), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n543), .A2(new_n554), .A3(new_n528), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n193), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n562), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n689), .A2(new_n198), .A3(new_n690), .A4(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n688), .A2(KEYINPUT101), .A3(new_n696), .ZN(new_n700));
  XOR2_X1   g514(.A(new_n674), .B(KEYINPUT39), .Z(new_n701));
  NAND2_X1  g515(.A1(new_n629), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT40), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(new_n704), .B(KEYINPUT102), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n707));
  INV_X1    g521(.A(new_n674), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n386), .A2(new_n646), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n670), .B2(new_n709), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n386), .A2(new_n646), .A3(new_n708), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT103), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  AOI22_X1  g528(.A1(new_n621), .A2(new_n622), .B1(new_n625), .B2(new_n495), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(G902), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n430), .A3(new_n500), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT104), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n500), .A3(new_n719), .A4(new_n430), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n617), .A3(new_n648), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND3_X1  g538(.A1(new_n721), .A2(new_n617), .A3(new_n657), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  NAND4_X1  g540(.A1(new_n582), .A2(new_n429), .A3(new_n633), .A4(new_n664), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n718), .A2(new_n315), .A3(new_n720), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT105), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n718), .A2(new_n730), .A3(new_n315), .A4(new_n720), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n727), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n242), .ZN(G21));
  NAND2_X1  g547(.A1(new_n689), .A2(new_n315), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n610), .A2(new_n613), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n630), .A2(G472), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n543), .B1(new_n566), .B2(new_n550), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n545), .A2(new_n547), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n559), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n721), .A2(new_n633), .A3(new_n735), .A4(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G122), .ZN(G24));
  NAND2_X1  g559(.A1(new_n729), .A2(new_n731), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n664), .A2(new_n738), .A3(new_n741), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n709), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  AOI21_X1  g565(.A(new_n499), .B1(new_n504), .B2(new_n193), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n627), .B2(new_n499), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n620), .A2(new_n311), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n314), .A2(new_n305), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n711), .A2(new_n756), .A3(KEYINPUT42), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n582), .A2(new_n737), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n711), .A2(new_n756), .A3(new_n582), .A4(new_n616), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT42), .B1(new_n760), .B2(KEYINPUT106), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n617), .A2(new_n762), .A3(new_n711), .A4(new_n756), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n759), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n338), .ZN(G33));
  NAND3_X1  g579(.A1(new_n617), .A2(new_n675), .A3(new_n756), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT107), .B(G134), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G36));
  NAND4_X1  g582(.A1(new_n646), .A2(new_n372), .A3(new_n381), .A4(new_n385), .ZN(new_n769));
  AND2_X1   g583(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n770));
  NOR2_X1   g584(.A1(KEYINPUT108), .A2(KEYINPUT43), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n386), .ZN(new_n773));
  INV_X1    g587(.A(new_n771), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n646), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n690), .A2(new_n631), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT109), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT44), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT110), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n314), .A2(new_n198), .A3(new_n305), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n780), .B2(KEYINPUT44), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n505), .A2(new_n507), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n504), .A2(new_n787), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n499), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n509), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n500), .B1(new_n791), .B2(KEYINPUT46), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n790), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n793), .A2(KEYINPUT46), .A3(new_n510), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n430), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n701), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n785), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n782), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  XNOR2_X1  g614(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n795), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n430), .B(new_n801), .C1(new_n792), .C2(new_n794), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  OR4_X1    g619(.A1(new_n616), .A2(new_n582), .A3(new_n709), .A4(new_n783), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n320), .ZN(G42));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n809));
  NOR2_X1   g623(.A1(G952), .A2(G953), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n721), .B(new_n617), .C1(new_n648), .C2(new_n657), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n812));
  INV_X1    g626(.A(new_n427), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n813), .B2(new_n425), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n426), .A2(KEYINPUT113), .A3(new_n427), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n647), .B1(new_n386), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n632), .A2(new_n317), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n317), .B(new_n512), .C1(new_n617), .C2(new_n665), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n811), .A2(new_n744), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n749), .A2(new_n756), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n816), .A2(new_n664), .A3(new_n708), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n655), .A2(new_n385), .A3(new_n372), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(new_n823), .A3(new_n783), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n582), .A3(new_n629), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n766), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  NOR4_X1   g640(.A1(new_n820), .A2(new_n764), .A3(new_n732), .A4(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n746), .A2(new_n749), .B1(new_n677), .B2(new_n680), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n664), .A2(new_n620), .A3(new_n674), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n695), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n734), .A2(new_n830), .A3(new_n753), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n710), .B2(new_n712), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(KEYINPUT52), .A2(new_n832), .A3(new_n750), .A4(new_n681), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n827), .B(KEYINPUT53), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n832), .A2(new_n750), .A3(new_n681), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n828), .A2(KEYINPUT52), .A3(new_n832), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT53), .B1(new_n841), .B2(new_n827), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n836), .A2(new_n842), .A3(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n836), .B2(new_n842), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n841), .A2(new_n827), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT114), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n845), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n850), .B2(KEYINPUT54), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n721), .A2(new_n688), .A3(new_n311), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n671), .B(new_n742), .C1(new_n772), .C2(new_n775), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT50), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n721), .A2(new_n688), .A3(new_n311), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n671), .B1(new_n772), .B2(new_n775), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n743), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT115), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n718), .A2(new_n720), .A3(new_n784), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n747), .A3(new_n857), .ZN(new_n863));
  INV_X1    g677(.A(new_n561), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n558), .A2(KEYINPUT32), .A3(new_n559), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n188), .A4(new_n694), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n614), .A3(new_n615), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n718), .A3(new_n720), .A4(new_n784), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n386), .A2(new_n646), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n716), .A2(new_n500), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n620), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n803), .A2(new_n804), .A3(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n858), .A2(new_n783), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n853), .A2(KEYINPUT50), .A3(new_n854), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n859), .B1(new_n856), .B2(new_n858), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n861), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n758), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n862), .A2(new_n884), .A3(new_n857), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT48), .ZN(new_n886));
  INV_X1    g700(.A(G953), .ZN(new_n887));
  OAI211_X1 g701(.A(G952), .B(new_n887), .C1(new_n868), .C2(new_n647), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n746), .B2(new_n854), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n889), .A3(KEYINPUT116), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n882), .B1(new_n877), .B2(new_n879), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n876), .A2(new_n895), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n852), .A2(new_n883), .A3(new_n894), .A4(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n892), .A2(new_n893), .B1(new_n876), .B2(new_n895), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n852), .B1(new_n898), .B2(new_n883), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n810), .B1(new_n851), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT49), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n737), .A2(new_n754), .ZN(new_n903));
  OAI22_X1  g717(.A1(new_n872), .A2(new_n902), .B1(new_n903), .B2(KEYINPUT112), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(KEYINPUT112), .B2(new_n903), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n769), .B(new_n695), .C1(new_n872), .C2(new_n902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n688), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n809), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n848), .A2(new_n910), .A3(new_n835), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n842), .A2(new_n844), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n848), .A2(new_n835), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n844), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n900), .B(new_n911), .C1(new_n914), .C2(new_n910), .ZN(new_n915));
  INV_X1    g729(.A(new_n810), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n917), .A2(KEYINPUT118), .A3(new_n907), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n909), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n191), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n913), .A2(G902), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT56), .B1(new_n923), .B2(G210), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n256), .A2(new_n261), .A3(new_n291), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(new_n289), .Z(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT55), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n921), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n924), .B2(new_n928), .ZN(G51));
  NAND2_X1  g744(.A1(new_n913), .A2(KEYINPUT54), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(KEYINPUT119), .A3(new_n911), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n913), .A2(new_n933), .A3(KEYINPUT54), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n509), .B(KEYINPUT57), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n498), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n793), .B(KEYINPUT120), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n923), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n920), .B1(new_n937), .B2(new_n939), .ZN(G54));
  NAND2_X1  g754(.A1(KEYINPUT58), .A2(G475), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n922), .A2(new_n653), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n653), .B1(new_n922), .B2(new_n941), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n921), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n942), .A2(new_n946), .A3(new_n921), .A4(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(G60));
  OR2_X1    g762(.A1(new_n641), .A2(new_n643), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(new_n638), .ZN(new_n950));
  INV_X1    g764(.A(new_n851), .ZN(new_n951));
  XNOR2_X1  g765(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n952));
  NAND2_X1  g766(.A1(G478), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  AND4_X1   g769(.A1(new_n950), .A2(new_n932), .A3(new_n934), .A4(new_n954), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n955), .A2(new_n956), .A3(new_n920), .ZN(G63));
  NAND2_X1  g771(.A1(G217), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT60), .Z(new_n959));
  AOI21_X1  g773(.A(new_n611), .B1(new_n913), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT124), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n921), .B1(new_n961), .B2(KEYINPUT61), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n913), .A2(new_n964), .A3(new_n662), .A4(new_n959), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n913), .A2(new_n662), .A3(new_n959), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT123), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n961), .A2(KEYINPUT61), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G66));
  INV_X1    g784(.A(new_n196), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n887), .B1(new_n971), .B2(G224), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n820), .A2(new_n732), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n974), .B2(new_n191), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n925), .B1(G898), .B2(new_n191), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT125), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  AND2_X1   g792(.A1(new_n521), .A2(new_n526), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(new_n374), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n828), .A2(new_n713), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n705), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  INV_X1    g798(.A(new_n807), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n705), .A2(new_n986), .A3(new_n982), .ZN(new_n987));
  INV_X1    g801(.A(new_n702), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(new_n617), .A3(new_n784), .A4(new_n817), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n799), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n990), .A2(new_n192), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n192), .A2(G227), .A3(G900), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n980), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n995));
  INV_X1    g809(.A(G227), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n996), .A3(G900), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n192), .B(new_n997), .C1(new_n995), .C2(G900), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n980), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n799), .A2(new_n982), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n734), .A2(new_n758), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n766), .B1(new_n797), .B2(new_n1002), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n1000), .A2(new_n764), .A3(new_n807), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n999), .B1(new_n1004), .B2(new_n191), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n994), .A2(new_n1005), .ZN(G72));
  NOR2_X1   g820(.A1(new_n990), .A2(new_n974), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  AOI211_X1 g824(.A(new_n543), .B(new_n529), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n546), .A2(new_n544), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1010), .ZN(new_n1013));
  NOR4_X1   g827(.A1(new_n914), .A2(new_n691), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1004), .A2(new_n973), .ZN(new_n1015));
  AOI211_X1 g829(.A(new_n544), .B(new_n546), .C1(new_n1015), .C2(new_n1010), .ZN(new_n1016));
  NOR4_X1   g830(.A1(new_n1011), .A2(new_n1014), .A3(new_n1016), .A4(new_n920), .ZN(G57));
endmodule


