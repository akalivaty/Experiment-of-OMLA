//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  AOI22_X1  g002(.A1(new_n202), .A2(new_n203), .B1(G211gat), .B2(G218gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(new_n202), .B2(new_n203), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n208), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(new_n205), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n218), .B2(new_n214), .ZN(new_n219));
  NOR2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(KEYINPUT64), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G169gat), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT23), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT25), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n223), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n220), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n219), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n231), .B1(new_n237), .B2(new_n230), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n232), .A3(KEYINPUT65), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT27), .B(G183gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n217), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n218), .B1(new_n242), .B2(KEYINPUT28), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n216), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT27), .B1(new_n216), .B2(KEYINPUT66), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT28), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n217), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n248));
  OAI22_X1  g047(.A1(new_n248), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT26), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n249), .A2(KEYINPUT67), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(KEYINPUT67), .B2(new_n250), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n229), .ZN(new_n253));
  OAI221_X1 g052(.A(new_n243), .B1(new_n244), .B2(new_n247), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G226gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n240), .B(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n255), .A2(new_n256), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n259), .A2(KEYINPUT29), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n240), .B2(new_n254), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n213), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n212), .A3(new_n257), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT74), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n263), .A2(KEYINPUT74), .A3(new_n212), .A4(new_n257), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n269), .A2(KEYINPUT37), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT37), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G8gat), .B(G36gat), .Z(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT76), .ZN(new_n276));
  XNOR2_X1  g075(.A(G64gat), .B(G92gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n274), .A2(KEYINPUT38), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n273), .B1(new_n262), .B2(new_n264), .ZN(new_n281));
  AOI211_X1 g080(.A(new_n278), .B(new_n281), .C1(new_n268), .C2(new_n273), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n272), .A2(new_n280), .B1(new_n282), .B2(KEYINPUT38), .ZN(new_n283));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT0), .ZN(new_n285));
  XOR2_X1   g084(.A(G57gat), .B(G85gat), .Z(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n288));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n291));
  INV_X1    g090(.A(G113gat), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(G113gat), .B2(G120gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n289), .B(KEYINPUT68), .C1(new_n294), .C2(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G141gat), .B(G148gat), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n305), .B1(new_n307), .B2(KEYINPUT2), .ZN(new_n308));
  XNOR2_X1  g107(.A(G141gat), .B(G148gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT78), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n305), .B1(new_n306), .B2(KEYINPUT77), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n313));
  OAI221_X1 g112(.A(new_n312), .B1(KEYINPUT77), .B2(new_n305), .C1(new_n309), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT79), .B1(new_n301), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n315), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT79), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n300), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n315), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n288), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n300), .B1(KEYINPUT3), .B2(new_n315), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n323), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n301), .A2(new_n315), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n316), .A2(new_n319), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n328), .B(new_n330), .C1(new_n331), .C2(KEYINPUT4), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n331), .B2(KEYINPUT4), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n328), .A2(new_n288), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n287), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT6), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n268), .A2(new_n278), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(new_n337), .A3(new_n287), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT6), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n339), .B(new_n340), .C1(new_n343), .C2(new_n338), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n283), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347));
  INV_X1    g146(.A(G50gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT29), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n315), .B2(KEYINPUT3), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n212), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n355), .B2(new_n354), .ZN(new_n357));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n326), .B1(new_n213), .B2(KEYINPUT29), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n315), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n354), .A2(new_n213), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n211), .A2(KEYINPUT82), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n363), .A2(KEYINPUT29), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n209), .A2(KEYINPUT82), .A3(new_n211), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT3), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n362), .B1(new_n366), .B2(new_n317), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n358), .ZN(new_n368));
  INV_X1    g167(.A(G22gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n361), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n361), .B2(new_n368), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n352), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n361), .A2(new_n368), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G22gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n375), .A2(new_n370), .A3(new_n351), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT40), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n325), .A2(new_n327), .ZN(new_n381));
  INV_X1    g180(.A(new_n334), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  XOR2_X1   g182(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n323), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n287), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT39), .B1(new_n321), .B2(new_n323), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(new_n383), .B2(new_n323), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n379), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n388), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n390), .A2(KEYINPUT40), .A3(new_n287), .A4(new_n385), .ZN(new_n391));
  INV_X1    g190(.A(new_n338), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n269), .A2(new_n279), .A3(new_n271), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT30), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n395), .B(new_n279), .C1(new_n266), .C2(new_n267), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n340), .A2(new_n395), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n378), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n338), .A2(new_n401), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n324), .A2(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT80), .B1(new_n403), .B2(new_n287), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n402), .A2(new_n404), .A3(new_n342), .A4(new_n341), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n339), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT30), .B1(new_n268), .B2(new_n278), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(new_n396), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n394), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n377), .B(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n346), .A2(new_n400), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n240), .A2(new_n254), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT69), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT69), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n240), .A2(new_n416), .A3(new_n254), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n300), .A3(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n240), .A2(new_n416), .A3(new_n301), .A4(new_n254), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(G227gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(new_n256), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n413), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n413), .ZN(new_n425));
  AOI211_X1 g224(.A(new_n422), .B(new_n425), .C1(new_n418), .C2(new_n419), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT72), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT72), .B1(new_n424), .B2(new_n426), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n418), .A2(new_n422), .A3(new_n419), .ZN(new_n432));
  XNOR2_X1  g231(.A(G15gat), .B(G43gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT33), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(KEYINPUT32), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT70), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n432), .A2(new_n440), .A3(KEYINPUT32), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n432), .A2(new_n436), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n435), .B1(new_n432), .B2(KEYINPUT32), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n439), .A2(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n431), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(new_n441), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n443), .A2(new_n442), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n446), .A2(new_n447), .A3(new_n427), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT36), .B1(new_n445), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n447), .ZN(new_n450));
  INV_X1    g249(.A(new_n427), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT36), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n444), .A2(new_n427), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n412), .A2(new_n449), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT35), .B1(new_n373), .B2(new_n376), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n339), .B1(new_n343), .B2(new_n338), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(new_n399), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n427), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(new_n448), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n452), .A2(new_n454), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n408), .A2(new_n457), .A3(new_n394), .A4(new_n458), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT86), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n450), .A2(new_n430), .A3(new_n429), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n377), .A3(new_n454), .ZN(new_n470));
  OAI21_X1  g269(.A(KEYINPUT35), .B1(new_n470), .B2(new_n409), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT17), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n480));
  INV_X1    g279(.A(G36gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT91), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT91), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n480), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT92), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT92), .ZN(new_n488));
  NOR4_X1   g287(.A1(KEYINPUT91), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n484), .B1(new_n480), .B2(new_n481), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n491), .B2(new_n479), .ZN(new_n492));
  AND2_X1   g291(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(KEYINPUT89), .A2(G29gat), .ZN(new_n494));
  OAI21_X1  g293(.A(G36gat), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT90), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT89), .B(G29gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT90), .A3(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(G43gat), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n348), .ZN(new_n501));
  NAND2_X1  g300(.A1(G43gat), .A2(G50gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT15), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n501), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n497), .A2(new_n499), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NOR3_X1   g306(.A1(new_n487), .A2(new_n492), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n497), .A2(new_n499), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n479), .A2(new_n482), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n474), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(G8gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT93), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n515), .A2(G1gat), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT16), .B1(new_n515), .B2(G1gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n518), .B2(KEYINPUT94), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n518), .B1(G1gat), .B2(new_n514), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n509), .A2(new_n510), .ZN(new_n523));
  INV_X1    g322(.A(new_n504), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n486), .A2(KEYINPUT92), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n491), .A2(new_n488), .A3(new_n479), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n504), .A2(new_n506), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n526), .A2(new_n509), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(KEYINPUT17), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n512), .A2(new_n522), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT95), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n521), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n531), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n535), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n534), .B(new_n521), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n533), .B(KEYINPUT13), .Z(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n536), .A2(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n539), .A3(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n473), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT96), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT96), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n473), .A2(new_n557), .A3(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560));
  INV_X1    g359(.A(G57gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(G64gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(G57gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n562), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(G71gat), .ZN(new_n568));
  INV_X1    g367(.A(G78gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AND3_X1   g369(.A1(new_n570), .A2(KEYINPUT97), .A3(new_n566), .ZN(new_n571));
  AOI21_X1  g370(.A(KEYINPUT97), .B1(new_n570), .B2(new_n566), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n560), .B(new_n567), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n566), .A2(new_n565), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n563), .A2(G57gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n561), .A2(G64gat), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n566), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n570), .A2(KEYINPUT97), .A3(new_n566), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(KEYINPUT98), .B1(new_n567), .B2(new_n578), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n521), .B1(KEYINPUT21), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n586));
  AND2_X1   g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G127gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n588), .A2(G127gat), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  INV_X1    g392(.A(new_n585), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n594), .A3(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G155gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n592), .A2(new_n595), .A3(new_n600), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G85gat), .A2(G92gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT7), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT7), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G99gat), .B(G106gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n613), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n512), .A2(new_n530), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G190gat), .B(G218gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT99), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n617), .A2(new_n618), .ZN(new_n624));
  AND2_X1   g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n534), .A2(new_n624), .B1(KEYINPUT41), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n625), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n623), .B1(new_n620), .B2(new_n626), .ZN(new_n633));
  OR3_X1    g432(.A1(new_n628), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n628), .B2(new_n633), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n604), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n584), .A2(new_n624), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  INV_X1    g439(.A(new_n578), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n560), .B1(new_n577), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(new_n619), .A3(new_n573), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n584), .A2(KEYINPUT10), .A3(new_n624), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(G230gat), .A2(G233gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n639), .A2(new_n645), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n650), .B1(new_n651), .B2(new_n649), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT101), .ZN(new_n656));
  XNOR2_X1  g455(.A(G176gat), .B(G204gat), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT101), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n655), .B(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n657), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g464(.A(new_n650), .B(new_n663), .C1(new_n651), .C2(new_n649), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(KEYINPUT102), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n652), .A2(new_n668), .A3(new_n664), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n638), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n559), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n406), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n399), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT16), .B(G8gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n513), .B1(new_n673), .B2(new_n399), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT42), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n677), .B2(new_n678), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(G1325gat));
  INV_X1    g483(.A(new_n673), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n685), .A2(G15gat), .A3(new_n465), .ZN(new_n686));
  INV_X1    g485(.A(new_n455), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n453), .B1(new_n469), .B2(new_n454), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT103), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n449), .A2(new_n690), .A3(new_n455), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G15gat), .B1(new_n685), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n686), .A2(new_n694), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n673), .A2(new_n411), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(new_n604), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n636), .A3(new_n670), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n556), .B2(new_n558), .ZN(new_n701));
  INV_X1    g500(.A(new_n498), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n674), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n636), .A2(KEYINPUT44), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n456), .B2(new_n472), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n670), .B(KEYINPUT104), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n699), .A2(new_n709), .A3(new_n554), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n689), .A2(new_n412), .A3(new_n691), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n463), .B1(new_n460), .B2(new_n462), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT86), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n471), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n468), .B2(new_n471), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n636), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n708), .B(new_n710), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(new_n674), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n705), .B(new_n706), .C1(new_n702), .C2(new_n721), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n701), .A2(new_n481), .A3(new_n399), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(KEYINPUT46), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(KEYINPUT46), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n720), .A2(new_n399), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n724), .B(new_n725), .C1(new_n481), .C2(new_n726), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n701), .A2(new_n500), .A3(new_n462), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n720), .A2(new_n692), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(new_n500), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT47), .B(new_n728), .C1(new_n729), .C2(new_n500), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1330gat));
  AOI21_X1  g533(.A(new_n348), .B1(new_n720), .B2(new_n378), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n701), .A2(new_n348), .A3(new_n411), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737));
  OR3_X1    g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n718), .A2(new_n719), .ZN(new_n739));
  INV_X1    g538(.A(new_n708), .ZN(new_n740));
  INV_X1    g539(.A(new_n710), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n739), .A2(new_n411), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n742), .A2(KEYINPUT106), .A3(G50gat), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT106), .B1(new_n742), .B2(G50gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n743), .A2(new_n744), .A3(new_n736), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n738), .B1(new_n745), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g545(.A(new_n717), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n715), .A3(new_n711), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n638), .A2(new_n709), .A3(new_n554), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(KEYINPUT107), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n406), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n561), .ZN(G1332gat));
  INV_X1    g555(.A(new_n399), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n754), .B2(new_n693), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n752), .A2(new_n568), .A3(new_n462), .A4(new_n753), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(G1334gat));
  INV_X1    g567(.A(new_n411), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(new_n569), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n604), .A2(new_n554), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n671), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n739), .A2(new_n740), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT109), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n739), .A2(new_n777), .A3(new_n740), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n406), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n748), .A2(new_n781), .A3(new_n636), .A4(new_n772), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n636), .B(new_n772), .C1(new_n716), .C2(new_n717), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT51), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n674), .A2(new_n611), .A3(new_n671), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(G1336gat));
  OAI21_X1  g586(.A(G92gat), .B1(new_n775), .B2(new_n757), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n757), .A2(new_n709), .A3(G92gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n782), .A2(new_n784), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n779), .B2(new_n757), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n781), .A2(KEYINPUT111), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n783), .B(new_n794), .Z(new_n795));
  XOR2_X1   g594(.A(new_n789), .B(KEYINPUT110), .Z(new_n796));
  AOI21_X1  g595(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n791), .B1(new_n792), .B2(new_n797), .ZN(G1337gat));
  XOR2_X1   g597(.A(KEYINPUT112), .B(G99gat), .Z(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n779), .B2(new_n693), .ZN(new_n800));
  OR3_X1    g599(.A1(new_n465), .A2(new_n670), .A3(new_n799), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n785), .B2(new_n801), .ZN(G1338gat));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803));
  INV_X1    g602(.A(G106gat), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n708), .B(new_n773), .C1(new_n718), .C2(new_n719), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n378), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n709), .A2(G106gat), .A3(new_n377), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n782), .A2(new_n784), .A3(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n803), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G106gat), .B1(new_n775), .B2(new_n377), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(KEYINPUT113), .A3(new_n809), .A4(new_n808), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n776), .A2(new_n411), .A3(new_n778), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n815), .A2(G106gat), .B1(new_n795), .B2(new_n807), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n814), .B1(new_n816), .B2(new_n809), .ZN(G1339gat));
  NOR2_X1   g616(.A1(new_n540), .A2(new_n541), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n533), .B1(new_n531), .B2(new_n535), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n548), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n667), .A2(new_n553), .A3(new_n669), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n649), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n646), .A2(new_n647), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n822), .B1(new_n646), .B2(new_n647), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n663), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n824), .A2(new_n827), .A3(KEYINPUT114), .A4(KEYINPUT55), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(new_n824), .B2(new_n827), .ZN(new_n833));
  INV_X1    g632(.A(new_n666), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AND4_X1   g635(.A1(new_n539), .A2(new_n538), .A3(new_n542), .A4(new_n549), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n549), .B1(new_n552), .B2(new_n539), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n821), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(KEYINPUT115), .B(new_n821), .C1(new_n836), .C2(new_n839), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n637), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n836), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n845), .A2(new_n553), .A3(new_n636), .A4(new_n820), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n604), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n638), .A2(new_n554), .A3(new_n671), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n843), .A2(new_n637), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n554), .A2(new_n832), .A3(new_n835), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT115), .B1(new_n851), .B2(new_n821), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n846), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n699), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  INV_X1    g654(.A(new_n848), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n406), .A2(new_n399), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n769), .A2(new_n462), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n292), .B1(new_n862), .B2(new_n554), .ZN(new_n863));
  XOR2_X1   g662(.A(new_n863), .B(KEYINPUT117), .Z(new_n864));
  INV_X1    g663(.A(new_n470), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n857), .A3(new_n674), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n866), .A2(new_n867), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n757), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n554), .A2(new_n292), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(G1340gat));
  NAND2_X1  g671(.A1(new_n671), .A2(new_n293), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875));
  INV_X1    g674(.A(new_n862), .ZN(new_n876));
  OAI21_X1  g675(.A(G120gat), .B1(new_n876), .B2(new_n709), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n874), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n875), .B1(new_n874), .B2(new_n877), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n876), .B2(new_n699), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n699), .A2(G127gat), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n870), .B2(new_n882), .ZN(G1342gat));
  NOR3_X1   g682(.A1(new_n399), .A2(G134gat), .A3(new_n637), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n855), .B1(new_n854), .B2(new_n856), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT116), .B(new_n848), .C1(new_n853), .C2(new_n699), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n674), .A4(new_n865), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n866), .A2(new_n867), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n862), .A2(new_n636), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n891), .A2(new_n892), .B1(G134gat), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n884), .B1(new_n868), .B2(new_n869), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(KEYINPUT56), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n891), .A2(KEYINPUT120), .A3(new_n892), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT121), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n901), .B(new_n894), .C1(new_n897), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1343gat));
  NOR2_X1   g702(.A1(new_n858), .A2(new_n377), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n693), .A2(new_n859), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n840), .A2(new_n637), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n604), .B1(new_n908), .B2(new_n846), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n411), .B1(new_n909), .B2(new_n848), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(KEYINPUT57), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n839), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n692), .A2(new_n377), .ZN(new_n914));
  AND4_X1   g713(.A1(new_n674), .A2(new_n888), .A3(new_n757), .A4(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n839), .A2(G141gat), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n915), .A2(new_n916), .B1(KEYINPUT122), .B2(KEYINPUT58), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g717(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1344gat));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(G148gat), .C1(new_n912), .C2(new_n670), .ZN(new_n922));
  INV_X1    g721(.A(G148gat), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n910), .A2(new_n905), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n907), .A2(new_n670), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n922), .B1(new_n928), .B2(new_n921), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n915), .A2(new_n923), .A3(new_n671), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1345gat));
  AOI21_X1  g730(.A(G155gat), .B1(new_n915), .B2(new_n604), .ZN(new_n932));
  INV_X1    g731(.A(new_n912), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n604), .A2(G155gat), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT123), .Z(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n933), .B2(new_n935), .ZN(G1346gat));
  AND3_X1   g735(.A1(new_n933), .A2(G162gat), .A3(new_n636), .ZN(new_n937));
  AOI21_X1  g736(.A(G162gat), .B1(new_n915), .B2(new_n636), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n937), .A2(new_n938), .ZN(G1347gat));
  NOR2_X1   g738(.A1(new_n674), .A2(new_n757), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT124), .Z(new_n941));
  NAND4_X1  g740(.A1(new_n888), .A2(new_n769), .A3(new_n462), .A4(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(new_n224), .A3(new_n839), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n858), .A2(new_n674), .A3(new_n757), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n865), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(new_n554), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n947), .B2(new_n224), .ZN(G1348gat));
  OAI21_X1  g747(.A(G176gat), .B1(new_n942), .B2(new_n709), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n671), .A2(new_n225), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n945), .B2(new_n950), .ZN(G1349gat));
  OAI21_X1  g750(.A(G183gat), .B1(new_n942), .B2(new_n699), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n604), .A2(new_n241), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n945), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n942), .B2(new_n637), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n958));
  OR2_X1    g757(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g758(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n217), .A3(new_n636), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n957), .A2(new_n958), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n961), .B(new_n962), .C1(new_n963), .C2(new_n959), .ZN(G1351gat));
  NAND2_X1  g763(.A1(new_n944), .A2(new_n914), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(G197gat), .B1(new_n966), .B2(new_n554), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n941), .A2(new_n693), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n968), .B1(new_n924), .B2(new_n925), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n554), .A2(G197gat), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1352gat));
  NOR3_X1   g770(.A1(new_n965), .A2(G204gat), .A3(new_n670), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT62), .ZN(new_n973));
  INV_X1    g772(.A(new_n969), .ZN(new_n974));
  OAI21_X1  g773(.A(G204gat), .B1(new_n974), .B2(new_n709), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(G1353gat));
  OR3_X1    g775(.A1(new_n965), .A2(G211gat), .A3(new_n699), .ZN(new_n977));
  OAI21_X1  g776(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n978), .B1(new_n969), .B2(new_n604), .ZN(new_n979));
  AND2_X1   g778(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  OAI21_X1  g782(.A(G218gat), .B1(new_n974), .B2(new_n637), .ZN(new_n984));
  OR3_X1    g783(.A1(new_n965), .A2(G218gat), .A3(new_n637), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1355gat));
endmodule


