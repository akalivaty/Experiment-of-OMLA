//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n540, new_n541, new_n542, new_n545,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n564, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n599, new_n600, new_n601, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(G137), .A3(new_n459), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n463), .A2(new_n466), .ZN(G160));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G136), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT66), .Z(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT67), .ZN(new_n476));
  OR2_X1    g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n459), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n476), .B1(G124), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n484), .B1(new_n468), .B2(new_n469), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n484), .B(new_n487), .C1(new_n469), .C2(new_n468), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  OR2_X1    g065(.A1(new_n459), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  AOI22_X1  g068(.A1(new_n479), .A2(G126), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n489), .B2(new_n494), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n495), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g075(.A(KEYINPUT69), .B(G651), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n498), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G50), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G88), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  OR2_X1    g083(.A1(new_n508), .A2(new_n501), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(G303));
  INV_X1    g085(.A(G303), .ZN(G166));
  XNOR2_X1  g086(.A(KEYINPUT70), .B(G51), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n502), .A2(G543), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n514), .A2(KEYINPUT7), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(KEYINPUT7), .ZN(new_n516));
  AND2_X1   g091(.A1(G63), .A2(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(new_n516), .B1(new_n505), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n502), .A2(new_n505), .ZN(new_n519));
  INV_X1    g094(.A(G89), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n513), .B(new_n518), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G168));
  NAND2_X1  g097(.A1(G77), .A2(G543), .ZN(new_n523));
  XOR2_X1   g098(.A(KEYINPUT5), .B(G543), .Z(new_n524));
  INV_X1    g099(.A(G64), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n501), .ZN(new_n529));
  OAI211_X1 g104(.A(KEYINPUT71), .B(new_n523), .C1(new_n524), .C2(new_n525), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT72), .ZN(new_n532));
  AOI22_X1  g107(.A1(G52), .A2(new_n503), .B1(new_n506), .B2(G90), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n528), .A2(new_n534), .A3(new_n529), .A4(new_n530), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  NAND2_X1  g112(.A1(new_n503), .A2(G43), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n502), .A2(G81), .A3(new_n505), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n501), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT73), .Z(G188));
  AOI22_X1  g123(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n499), .ZN(new_n550));
  INV_X1    g125(.A(G91), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT75), .B1(new_n519), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT75), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n502), .A2(new_n553), .A3(G91), .A4(new_n505), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n503), .A2(G53), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n502), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n555), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n521), .B(new_n564), .ZN(G286));
  NAND3_X1  g140(.A1(new_n502), .A2(G49), .A3(G543), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n502), .A2(G87), .A3(new_n505), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND3_X1  g144(.A1(new_n502), .A2(G86), .A3(new_n505), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT78), .ZN(new_n571));
  NAND2_X1  g146(.A1(G73), .A2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G61), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n524), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n574), .A2(KEYINPUT77), .A3(new_n529), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n577), .B2(new_n501), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n575), .A2(new_n578), .B1(new_n503), .B2(G48), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n571), .A2(new_n579), .ZN(G305));
  NAND2_X1  g155(.A1(new_n506), .A2(G85), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n503), .A2(G47), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n581), .B(new_n582), .C1(new_n501), .C2(new_n583), .ZN(G290));
  NAND3_X1  g159(.A1(new_n502), .A2(G92), .A3(new_n505), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n524), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n503), .A2(G54), .B1(G651), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G171), .B2(new_n593), .ZN(G284));
  OAI21_X1  g170(.A(new_n594), .B1(G171), .B2(new_n593), .ZN(G321));
  XNOR2_X1  g171(.A(new_n521), .B(KEYINPUT76), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n593), .ZN(new_n598));
  AOI211_X1 g173(.A(KEYINPUT79), .B(new_n598), .C1(new_n593), .C2(G299), .ZN(new_n599));
  AND2_X1   g174(.A1(new_n598), .A2(KEYINPUT79), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT80), .ZN(G297));
  XNOR2_X1  g177(.A(new_n601), .B(KEYINPUT81), .ZN(G280));
  AND2_X1   g178(.A1(new_n587), .A2(new_n591), .ZN(new_n604));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G860), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g182(.A1(new_n604), .A2(new_n605), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n479), .A2(G123), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n459), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  INV_X1    g189(.A(G135), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n460), .A2(new_n459), .ZN(new_n616));
  OAI221_X1 g191(.A(new_n612), .B1(new_n613), .B2(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2096), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n619), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT83), .Z(G156));
  XOR2_X1   g202(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n628));
  XOR2_X1   g203(.A(KEYINPUT15), .B(G2435), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n630), .B2(new_n631), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n633), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  XNOR2_X1  g219(.A(G2067), .B(G2678), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(new_n623), .ZN(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n646), .B2(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(new_n618), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1991), .B(G1996), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1971), .B(G1976), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  MUX2_X1   g241(.A(new_n666), .B(new_n665), .S(new_n658), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G1981), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1986), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n671), .A2(new_n673), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n656), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n671), .A2(new_n673), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n673), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n677), .A2(new_n655), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G35), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G162), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2090), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NOR2_X1   g262(.A1(G168), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n687), .B2(G21), .ZN(new_n689));
  INV_X1    g264(.A(G1966), .ZN(new_n690));
  NOR2_X1   g265(.A1(G16), .A2(G19), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n542), .B2(G16), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n689), .A2(new_n690), .B1(G1341), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G2078), .ZN(new_n694));
  NOR2_X1   g269(.A1(G164), .A2(new_n681), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G27), .B2(new_n681), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n686), .B(new_n693), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n687), .A2(G20), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT23), .Z(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G299), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1956), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n681), .A2(G33), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT94), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT25), .ZN(new_n706));
  NAND2_X1  g281(.A1(G115), .A2(G2104), .ZN(new_n707));
  INV_X1    g282(.A(G127), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n470), .B2(new_n708), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n709), .A2(G2105), .B1(new_n471), .B2(G139), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n703), .B1(new_n713), .B2(new_n681), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2072), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n681), .A2(G32), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n471), .A2(G141), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT96), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT26), .Z(new_n720));
  NAND2_X1  g295(.A1(new_n479), .A2(G129), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n718), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n716), .B1(new_n724), .B2(new_n681), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT30), .B(G28), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT31), .A2(G11), .ZN(new_n729));
  NAND2_X1  g304(.A1(KEYINPUT31), .A2(G11), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n728), .A2(new_n681), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n617), .B2(new_n681), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n681), .B1(new_n733), .B2(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n733), .B2(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G160), .B2(G29), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n732), .B1(new_n736), .B2(G2084), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n727), .B(new_n737), .C1(G2084), .C2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n696), .A2(new_n694), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G1341), .B2(new_n692), .ZN(new_n740));
  OR4_X1    g315(.A1(new_n702), .A2(new_n715), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n742));
  INV_X1    g317(.A(G116), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G2105), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT92), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G140), .B2(new_n471), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n479), .A2(G128), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT91), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G29), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT93), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n681), .A2(G26), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT28), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G171), .A2(new_n687), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G5), .B2(new_n687), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G4), .A2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT90), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n592), .B2(new_n687), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1348), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n756), .A2(new_n760), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n689), .A2(new_n690), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(new_n759), .B2(new_n758), .ZN(new_n768));
  NOR4_X1   g343(.A1(new_n697), .A2(new_n741), .A3(new_n765), .A4(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  MUX2_X1   g345(.A(G6), .B(G305), .S(G16), .Z(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT32), .B(G1981), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n773), .A2(KEYINPUT87), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(KEYINPUT87), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n687), .A2(G22), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G166), .B2(new_n687), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1971), .Z(new_n778));
  NAND3_X1  g353(.A1(new_n774), .A2(new_n775), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT88), .ZN(new_n780));
  NAND2_X1  g355(.A1(G288), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT88), .A4(new_n568), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G23), .B(new_n783), .S(G16), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G1976), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(KEYINPUT34), .B1(new_n779), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n775), .A2(new_n778), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n786), .B(G1976), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT34), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n790), .A2(new_n791), .A3(new_n792), .A4(new_n774), .ZN(new_n793));
  MUX2_X1   g368(.A(G24), .B(G290), .S(G16), .Z(new_n794));
  XOR2_X1   g369(.A(KEYINPUT86), .B(G1986), .Z(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n681), .A2(G25), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n471), .A2(G131), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n479), .A2(G119), .ZN(new_n799));
  OR2_X1    g374(.A1(G95), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n681), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT35), .B(G1991), .Z(new_n805));
  XOR2_X1   g380(.A(new_n804), .B(new_n805), .Z(new_n806));
  OR2_X1    g381(.A1(new_n796), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n794), .B2(new_n795), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n789), .A2(new_n793), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n770), .B1(new_n810), .B2(new_n811), .ZN(G311));
  INV_X1    g387(.A(new_n810), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n769), .B1(new_n813), .B2(new_n814), .ZN(G150));
  NOR2_X1   g390(.A1(new_n592), .A2(new_n605), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT38), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(new_n501), .ZN(new_n819));
  INV_X1    g394(.A(G55), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT99), .B(G93), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n819), .B1(new_n559), .B2(new_n820), .C1(new_n519), .C2(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n542), .B(new_n822), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n817), .B(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(KEYINPUT39), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n825), .A2(new_n826), .A3(G860), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n822), .A2(G860), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n827), .A2(new_n829), .ZN(G145));
  INV_X1    g405(.A(G37), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n479), .A2(G130), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n459), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G142), .B2(new_n471), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n621), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n802), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n724), .A2(new_n749), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n489), .A2(new_n494), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n724), .A2(new_n749), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n842), .ZN(new_n845));
  INV_X1    g420(.A(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n846), .B2(new_n840), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n711), .B(KEYINPUT95), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n844), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n713), .A2(new_n852), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n844), .A2(new_n847), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n832), .B(new_n839), .C1(new_n851), .C2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n839), .A2(new_n832), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n844), .A2(new_n847), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n849), .A2(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n839), .A2(new_n832), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n856), .A2(new_n859), .A3(new_n860), .A4(new_n850), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n617), .B(G160), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n481), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n855), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n863), .B1(new_n855), .B2(new_n861), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT102), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  AOI211_X1 g442(.A(new_n867), .B(new_n863), .C1(new_n855), .C2(new_n861), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n831), .B(new_n864), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g445(.A(G305), .B(new_n783), .Z(new_n871));
  XNOR2_X1  g446(.A(G290), .B(G303), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n542), .B(new_n822), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n608), .ZN(new_n877));
  INV_X1    g452(.A(G299), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n592), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n604), .A2(G299), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT41), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n880), .A3(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n877), .B2(new_n887), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n874), .B(new_n875), .C1(new_n888), .C2(KEYINPUT103), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(KEYINPUT103), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n888), .A2(new_n875), .A3(KEYINPUT103), .A4(new_n874), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  MUX2_X1   g468(.A(new_n822), .B(new_n893), .S(G868), .Z(G295));
  MUX2_X1   g469(.A(new_n822), .B(new_n893), .S(G868), .Z(G331));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n896));
  NAND2_X1  g471(.A1(G301), .A2(new_n521), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(G301), .B2(G286), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n823), .A2(new_n898), .A3(KEYINPUT106), .ZN(new_n899));
  NAND2_X1  g474(.A1(G171), .A2(new_n597), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n876), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n823), .A2(new_n898), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(new_n902), .A2(new_n905), .B1(new_n886), .B2(new_n885), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n881), .A3(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT108), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n903), .A2(new_n909), .A3(new_n901), .A4(new_n881), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n873), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n901), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n876), .B1(new_n897), .B2(new_n900), .ZN(new_n914));
  INV_X1    g489(.A(new_n886), .ZN(new_n915));
  AOI21_X1  g490(.A(KEYINPUT41), .B1(new_n879), .B2(new_n880), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n913), .A2(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n887), .B(KEYINPUT105), .C1(new_n914), .C2(new_n913), .ZN(new_n920));
  INV_X1    g495(.A(new_n873), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n905), .A2(new_n881), .A3(new_n899), .A4(new_n901), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n912), .A2(new_n831), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT43), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(new_n922), .A3(new_n920), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n873), .A2(KEYINPUT107), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G37), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n919), .A2(new_n927), .A3(new_n922), .A4(new_n920), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n896), .B1(new_n925), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n930), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n924), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n930), .B1(new_n929), .B2(new_n931), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n933), .B1(new_n896), .B2(new_n937), .ZN(G397));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n842), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n941));
  INV_X1    g516(.A(G40), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n463), .A2(new_n466), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n749), .B(new_n755), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n724), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT125), .B(KEYINPUT46), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT125), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT46), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n944), .A2(G1996), .ZN(new_n951));
  MUX2_X1   g526(.A(new_n948), .B(new_n950), .S(new_n951), .Z(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(KEYINPUT47), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n724), .B(G1996), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n944), .B1(new_n957), .B2(new_n945), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT110), .ZN(new_n959));
  INV_X1    g534(.A(new_n944), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n802), .B(new_n805), .Z(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OR3_X1    g537(.A1(new_n944), .A2(G290), .A3(G1986), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT48), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n803), .A2(new_n805), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n959), .A2(new_n965), .B1(G2067), .B2(new_n749), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n962), .A2(new_n964), .B1(new_n966), .B2(new_n960), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n956), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT47), .B1(new_n954), .B2(new_n955), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n489), .B2(new_n494), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n488), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n487), .B1(new_n460), .B2(new_n484), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n479), .A2(G126), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n491), .A2(new_n493), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT68), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n982));
  AOI21_X1  g557(.A(G1384), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n974), .B1(new_n983), .B2(KEYINPUT45), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n939), .B1(new_n495), .B2(new_n496), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n973), .A3(new_n941), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n984), .A2(new_n694), .A3(new_n986), .A4(new_n943), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT122), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n988), .A2(G2078), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n972), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n943), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G125), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n462), .B1(new_n470), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G2105), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(G40), .A3(new_n465), .A4(new_n464), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n998), .B1(new_n940), .B2(new_n941), .ZN(new_n999));
  INV_X1    g574(.A(new_n991), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n1000), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(KEYINPUT122), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n998), .B1(new_n1003), .B2(new_n971), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n983), .B2(new_n1003), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT121), .B(G1961), .Z(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n994), .A2(new_n1002), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n989), .A2(G301), .A3(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n999), .B(new_n991), .C1(new_n985), .C2(new_n941), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1003), .B(new_n939), .C1(new_n977), .C2(new_n980), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n943), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1013), .B2(new_n1006), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n988), .B2(new_n987), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1009), .B1(new_n1015), .B2(G301), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n999), .B1(new_n985), .B2(new_n941), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n690), .ZN(new_n1019));
  INV_X1    g594(.A(G2084), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1020), .B(new_n1004), .C1(new_n983), .C2(new_n1003), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(G168), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(G8), .ZN(new_n1023));
  AOI21_X1  g598(.A(G168), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT51), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1026), .A3(G8), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1016), .A2(new_n1017), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G303), .A2(G8), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT55), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1003), .B(new_n939), .C1(new_n495), .C2(new_n496), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n998), .B1(new_n940), .B2(KEYINPUT50), .ZN(new_n1032));
  XOR2_X1   g607(.A(KEYINPUT113), .B(G2090), .Z(new_n1033));
  AND3_X1   g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n984), .A2(new_n986), .A3(new_n943), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT112), .B(G1971), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1034), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G8), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1030), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1030), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n985), .A2(new_n941), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n998), .B1(new_n1042), .B2(new_n974), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1036), .B1(new_n1043), .B2(new_n986), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1013), .A2(new_n1033), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(G8), .B(new_n1041), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT49), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n571), .A2(new_n669), .A3(new_n579), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n669), .B1(new_n579), .B2(new_n570), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n579), .A2(new_n570), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G1981), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n571), .A2(new_n669), .A3(new_n579), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(KEYINPUT49), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1039), .B1(new_n943), .B2(new_n971), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1051), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n781), .A2(G1976), .A3(new_n782), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n1056), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1059), .A2(new_n1056), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n787), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1040), .A2(new_n1047), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT123), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT124), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n992), .A2(new_n993), .A3(new_n990), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT122), .B1(new_n999), .B2(new_n1001), .ZN(new_n1069));
  OAI22_X1  g644(.A1(new_n1068), .A2(new_n1069), .B1(new_n1013), .B2(new_n1006), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(new_n988), .B2(new_n987), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1067), .B1(new_n1071), .B2(G301), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n989), .A2(new_n1008), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1073), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1017), .B1(new_n1015), .B2(G301), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1040), .A2(new_n1047), .A3(new_n1064), .A4(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1028), .A2(new_n1066), .A3(new_n1076), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n701), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1082), .B(KEYINPUT118), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1081), .B1(new_n1035), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n562), .B1(new_n555), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g663(.A(KEYINPUT116), .B(new_n550), .C1(new_n552), .C2(new_n554), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT117), .B(new_n1086), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1085), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n940), .A2(new_n998), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1013), .A2(G1348), .B1(G2067), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g675(.A(KEYINPUT119), .B1(G2067), .B2(new_n1097), .C1(new_n1013), .C2(G1348), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1095), .B1(new_n592), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1043), .A2(new_n986), .A3(new_n1083), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1094), .A2(new_n1093), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1081), .B(new_n1104), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n592), .B1(new_n1102), .B2(KEYINPUT60), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n1110), .B(new_n604), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1109), .A2(new_n1111), .B1(KEYINPUT60), .B2(new_n1102), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT120), .B(G1996), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1035), .A2(new_n1113), .B1(new_n1096), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n542), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT59), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1107), .A2(new_n1095), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1107), .A2(new_n1095), .A3(KEYINPUT61), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1112), .A2(new_n1117), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1079), .B1(new_n1108), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1065), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1020), .A2(new_n1013), .B1(new_n1018), .B2(new_n690), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1125), .A2(new_n1039), .A3(G286), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT63), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1047), .A2(new_n1126), .A3(KEYINPUT63), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT114), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1035), .A2(new_n1037), .B1(new_n1033), .B2(new_n1013), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n1039), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT114), .B(G8), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1030), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1064), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1128), .B1(new_n1134), .B2(KEYINPUT115), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT115), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1136), .A3(new_n1064), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1127), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1047), .ZN(new_n1139));
  INV_X1    g714(.A(G288), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1057), .A2(new_n787), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1054), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1139), .A2(new_n1064), .B1(new_n1142), .B2(new_n1056), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT62), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1015), .A2(G301), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1025), .A2(new_n1147), .A3(new_n1027), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1066), .A2(new_n1078), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1143), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1123), .A2(new_n1138), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n960), .A2(G1986), .A3(G290), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n963), .A2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT109), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n962), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n970), .B1(new_n1152), .B2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g732(.A1(G401), .A2(new_n457), .A3(G227), .ZN(new_n1159));
  AND3_X1   g733(.A1(new_n676), .A2(new_n679), .A3(new_n1159), .ZN(new_n1160));
  OAI211_X1 g734(.A(new_n1160), .B(new_n869), .C1(new_n936), .C2(new_n935), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


