//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR3_X1   g0012(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G116), .ZN(new_n217));
  INV_X1    g0017(.A(G270), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n220), .B1(new_n201), .B2(new_n221), .C1(new_n203), .C2(new_n222), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n219), .B(new_n223), .C1(G97), .C2(G257), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(G1), .B2(G20), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT1), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n227), .A2(new_n212), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n202), .A2(new_n203), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n215), .B(new_n226), .C1(new_n228), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT14), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT66), .A2(G45), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT66), .A2(G45), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(new_n211), .A3(G274), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G238), .A3(new_n258), .ZN(new_n259));
  OR2_X1    g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G232), .A2(G1698), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n221), .B2(G1698), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n262), .A2(new_n264), .B1(G33), .B2(G97), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n255), .B(new_n259), .C1(new_n265), .C2(new_n257), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT73), .B1(new_n266), .B2(KEYINPUT13), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(new_n264), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n257), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n253), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT66), .A2(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G41), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n211), .A2(G274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n259), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT73), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n271), .A2(new_n277), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(KEYINPUT74), .B(KEYINPUT13), .C1(new_n270), .C2(new_n276), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT74), .B1(new_n266), .B2(KEYINPUT13), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n267), .B(new_n280), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n250), .B1(new_n284), .B2(G169), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n271), .A2(new_n277), .A3(new_n279), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n266), .A2(KEYINPUT13), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G179), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n284), .A2(new_n250), .A3(G169), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n286), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n227), .ZN(new_n294));
  INV_X1    g0094(.A(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G77), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n297), .A2(new_n298), .B1(new_n201), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n212), .A2(G68), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT11), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n294), .B1(new_n211), .B2(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  OAI22_X1  g0106(.A1(new_n303), .A2(new_n304), .B1(new_n203), .B2(new_n306), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n303), .A2(new_n304), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n302), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT12), .Z(new_n312));
  OR3_X1    g0112(.A1(new_n307), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n292), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G223), .A2(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G1698), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G222), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n262), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n257), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n320), .C1(G77), .C2(new_n262), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n257), .A2(new_n258), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G226), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n321), .A2(new_n255), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n204), .A2(G20), .ZN(new_n329));
  INV_X1    g0129(.A(G150), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n329), .B1(new_n330), .B2(new_n300), .C1(new_n331), .C2(new_n297), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n310), .A2(G20), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n332), .A2(new_n294), .B1(new_n201), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n305), .A2(G50), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n325), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n328), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT67), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n287), .A2(new_n288), .A3(G190), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n313), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n284), .A2(G200), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n333), .A2(G77), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n306), .A2(new_n298), .ZN(new_n351));
  OR2_X1    g0151(.A1(KEYINPUT15), .A2(G87), .ZN(new_n352));
  NAND2_X1  g0152(.A1(KEYINPUT15), .A2(G87), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(KEYINPUT70), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT70), .ZN(new_n355));
  AND2_X1   g0155(.A1(KEYINPUT15), .A2(G87), .ZN(new_n356));
  NOR2_X1   g0156(.A1(KEYINPUT15), .A2(G87), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT71), .B1(new_n359), .B2(new_n297), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G20), .A2(G77), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT71), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n354), .A2(new_n358), .A3(new_n362), .A4(new_n296), .ZN(new_n363));
  INV_X1    g0163(.A(new_n331), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n299), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n360), .A2(new_n361), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  AOI211_X1 g0166(.A(new_n350), .B(new_n351), .C1(new_n366), .C2(new_n294), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n234), .A2(G1698), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n222), .A2(new_n317), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n262), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(KEYINPUT68), .A2(G107), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT68), .A2(G107), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  NOR2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT69), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n370), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n379), .B1(new_n370), .B2(new_n378), .ZN(new_n382));
  NOR3_X1   g0182(.A1(new_n381), .A2(new_n382), .A3(new_n257), .ZN(new_n383));
  INV_X1    g0183(.A(G244), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n255), .B1(new_n384), .B2(new_n322), .ZN(new_n385));
  OAI21_X1  g0185(.A(G200), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n382), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n320), .A3(new_n380), .ZN(new_n388));
  INV_X1    g0188(.A(new_n385), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G190), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n367), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n343), .A2(new_n349), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(G169), .B1(new_n388), .B2(new_n389), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT72), .B1(new_n367), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(new_n327), .A3(new_n389), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n366), .A2(new_n294), .ZN(new_n396));
  INV_X1    g0196(.A(new_n350), .ZN(new_n397));
  INV_X1    g0197(.A(new_n351), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n338), .B1(new_n383), .B2(new_n385), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT72), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n394), .A2(new_n395), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n315), .A2(new_n392), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n337), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT9), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT9), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n337), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n325), .A2(G200), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n326), .A2(G190), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n407), .A2(new_n409), .A3(new_n410), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT10), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n406), .A2(KEYINPUT9), .B1(G190), .B2(new_n326), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT10), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n414), .A2(new_n415), .A3(new_n410), .A4(new_n409), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT16), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G58), .A2(G68), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n212), .B1(new_n229), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n260), .A2(new_n212), .A3(new_n261), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n261), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n421), .B1(new_n426), .B2(G68), .ZN(new_n427));
  INV_X1    g0227(.A(G159), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n300), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n419), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n203), .B1(new_n424), .B2(new_n425), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n432), .A2(KEYINPUT16), .A3(new_n429), .A4(new_n421), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n294), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n364), .A2(new_n333), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n305), .A2(new_n364), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n221), .A2(G1698), .ZN(new_n439));
  OAI221_X1 g0239(.A(new_n439), .B1(G223), .B2(G1698), .C1(new_n375), .C2(new_n376), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G87), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n320), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT76), .B1(new_n322), .B2(new_n234), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n257), .A2(new_n258), .A3(new_n445), .A4(G232), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n447), .A3(new_n255), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G179), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n449), .B1(new_n338), .B2(new_n448), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n438), .A2(KEYINPUT18), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT18), .B1(new_n438), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G200), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(G190), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n443), .A2(new_n447), .A3(new_n456), .A4(new_n255), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n434), .A2(new_n436), .A3(new_n458), .A4(new_n437), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NOR3_X1   g0261(.A1(new_n418), .A2(new_n453), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n405), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(G250), .A2(G1698), .ZN(new_n464));
  OAI221_X1 g0264(.A(new_n464), .B1(G257), .B2(new_n317), .C1(new_n375), .C2(new_n376), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT84), .B(G294), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G33), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n257), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n473), .A2(G264), .A3(new_n257), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n470), .B(G274), .C1(new_n472), .C2(new_n471), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n468), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G179), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n338), .B2(new_n477), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n212), .B(G87), .C1(new_n375), .C2(new_n376), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT22), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT22), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n262), .A2(new_n483), .A3(new_n212), .A4(G87), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT24), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT68), .B(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT23), .A3(G20), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT23), .B1(new_n207), .B2(G20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(G20), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n486), .B1(new_n485), .B2(new_n492), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n294), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n294), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n211), .A2(G33), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n496), .A2(new_n333), .A3(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G107), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n310), .A2(G20), .A3(new_n207), .ZN(new_n501));
  XNOR2_X1  g0301(.A(new_n501), .B(KEYINPUT82), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT25), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n495), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT83), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n495), .A2(KEYINPUT83), .A3(new_n500), .A4(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n480), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n509), .B(new_n212), .C1(G33), .C2(new_n206), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT80), .ZN(new_n511));
  AOI21_X1  g0311(.A(G20), .B1(new_n295), .B2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT80), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n509), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n217), .A2(G20), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n294), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n515), .A2(new_n517), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n516), .A2(G1), .A3(new_n309), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n499), .B2(G116), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n517), .A2(new_n511), .A3(new_n514), .A4(new_n519), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n520), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n522), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n473), .A2(new_n257), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G270), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n317), .A2(G257), .ZN(new_n530));
  NAND2_X1  g0330(.A1(G264), .A2(G1698), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n262), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  XOR2_X1   g0332(.A(KEYINPUT79), .B(G303), .Z(new_n533));
  OAI211_X1 g0333(.A(new_n532), .B(new_n320), .C1(new_n262), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n529), .A2(new_n534), .A3(new_n475), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n527), .A2(new_n536), .A3(G179), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n527), .A2(G169), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n527), .A2(new_n541), .A3(G169), .A4(new_n535), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n535), .A2(G200), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n456), .B2(new_n535), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n543), .B1(new_n527), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n333), .B1(new_n354), .B2(new_n358), .ZN(new_n547));
  INV_X1    g0347(.A(G87), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n498), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT78), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n206), .ZN(new_n551));
  INV_X1    g0351(.A(new_n373), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n551), .B1(new_n552), .B2(new_n371), .ZN(new_n553));
  NAND3_X1  g0353(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n212), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n550), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n262), .A2(new_n212), .A3(G68), .ZN(new_n558));
  OAI211_X1 g0358(.A(KEYINPUT78), .B(new_n555), .C1(new_n374), .C2(new_n551), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n297), .B2(new_n206), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  AOI211_X1 g0362(.A(new_n547), .B(new_n549), .C1(new_n562), .C2(new_n294), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n222), .A2(new_n317), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n384), .A2(G1698), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n375), .C2(new_n376), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n490), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT77), .B1(new_n566), .B2(new_n490), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n567), .A2(new_n568), .A3(new_n257), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n257), .B(G250), .C1(G1), .C2(new_n469), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n470), .A2(G274), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n569), .A2(G190), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n568), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n490), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n320), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n572), .ZN(new_n577));
  AOI21_X1  g0377(.A(G200), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n563), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n562), .A2(new_n294), .ZN(new_n580));
  INV_X1    g0380(.A(new_n547), .ZN(new_n581));
  INV_X1    g0381(.A(new_n359), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n499), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(new_n577), .A3(new_n327), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n338), .B1(new_n569), .B2(new_n572), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n579), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n485), .A2(new_n492), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT24), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n485), .A2(new_n486), .A3(new_n492), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n294), .B1(G107), .B2(new_n499), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n465), .A2(new_n467), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n320), .ZN(new_n595));
  INV_X1    g0395(.A(new_n474), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n595), .A2(new_n475), .A3(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(new_n456), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(G200), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n593), .A2(new_n503), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT4), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n262), .B2(G250), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(new_n317), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n602), .A2(G1698), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n605), .B(G244), .C1(new_n376), .C2(new_n375), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n384), .B1(new_n260), .B2(new_n261), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n606), .B(new_n509), .C1(new_n607), .C2(KEYINPUT4), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n320), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n528), .A2(G257), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n475), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n338), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n334), .A2(new_n206), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n499), .A2(G97), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n487), .B1(new_n424), .B2(new_n425), .ZN(new_n615));
  XNOR2_X1  g0415(.A(G97), .B(G107), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT6), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n212), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n300), .A2(new_n298), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n615), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n613), .B(new_n614), .C1(new_n622), .C2(new_n496), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n609), .A2(new_n327), .A3(new_n475), .A4(new_n610), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n612), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n622), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n294), .B1(new_n206), .B2(new_n334), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n611), .A2(G200), .ZN(new_n628));
  OAI21_X1  g0428(.A(G244), .B1(new_n375), .B2(new_n376), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n602), .B1(G33), .B2(G283), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n606), .C1(new_n317), .C2(new_n603), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(new_n320), .B1(G257), .B2(new_n528), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(G190), .A3(new_n475), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n627), .A2(new_n628), .A3(new_n633), .A4(new_n614), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n588), .A2(new_n601), .A3(new_n625), .A4(new_n634), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n463), .A2(new_n508), .A3(new_n546), .A4(new_n635), .ZN(G372));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n625), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n495), .A2(new_n500), .A3(new_n503), .A4(new_n600), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n587), .B(new_n579), .C1(new_n638), .C2(new_n598), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n504), .A2(new_n479), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n543), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n587), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n579), .A2(new_n587), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n625), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n612), .A2(new_n624), .A3(new_n623), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(KEYINPUT26), .A3(new_n587), .A4(new_n579), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n463), .B1(new_n643), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n349), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n314), .B1(new_n652), .B2(new_n403), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n459), .B(KEYINPUT17), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n453), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n343), .B1(new_n655), .B2(new_n418), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n651), .A2(new_n656), .ZN(G369));
  NOR2_X1   g0457(.A1(new_n309), .A2(G20), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n211), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n546), .B1(new_n527), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n540), .A2(new_n542), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n537), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n667), .A2(new_n527), .A3(new_n664), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G330), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n506), .A2(new_n507), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n479), .B2(new_n664), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n601), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n508), .A2(new_n664), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n543), .A2(new_n664), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n673), .A2(new_n601), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n664), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n504), .A2(new_n479), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n677), .A2(new_n683), .ZN(G399));
  NAND2_X1  g0484(.A1(new_n553), .A2(new_n217), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  INV_X1    g0486(.A(new_n213), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n686), .A2(new_n211), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(new_n231), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  INV_X1    g0491(.A(new_n639), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n634), .A2(new_n625), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n692), .B(new_n693), .C1(new_n508), .C2(new_n667), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n650), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n680), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT86), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(KEYINPUT86), .A3(new_n680), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(KEYINPUT29), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n664), .B1(new_n643), .B2(new_n650), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n632), .A2(G179), .A3(new_n475), .A4(new_n477), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n576), .A2(new_n577), .A3(new_n529), .A4(new_n534), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n477), .A2(G179), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n576), .A2(new_n577), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n611), .A3(new_n535), .A4(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n707), .ZN(new_n712));
  INV_X1    g0512(.A(new_n611), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n597), .A2(new_n327), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT30), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n708), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n664), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n719), .A3(new_n664), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n545), .A2(new_n527), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n667), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n508), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n640), .A3(new_n724), .A4(new_n680), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n704), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n691), .B1(new_n729), .B2(G1), .ZN(G364));
  NAND2_X1  g0530(.A1(new_n669), .A2(new_n670), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT87), .Z(new_n732));
  INV_X1    g0532(.A(new_n671), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n211), .B1(new_n658), .B2(G45), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n688), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n732), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n669), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n687), .A2(new_n262), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n272), .A2(new_n273), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n743), .B1(new_n230), .B2(new_n745), .C1(new_n245), .C2(new_n469), .ZN(new_n746));
  NAND3_X1  g0546(.A1(G355), .A2(new_n213), .A3(new_n262), .ZN(new_n747));
  OAI211_X1 g0547(.A(new_n746), .B(new_n747), .C1(G116), .C2(new_n213), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n227), .B1(G20), .B2(new_n338), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n741), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n212), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT89), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT89), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(G20), .A2(G179), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT88), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n756), .A2(new_n548), .B1(new_n201), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n752), .A2(new_n456), .A3(G200), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(G107), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G190), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n758), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n456), .A2(G200), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n758), .A2(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G77), .A2(new_n766), .B1(new_n768), .B2(G58), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n456), .A2(G179), .A3(G200), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n212), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n206), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n758), .A2(new_n456), .A3(G200), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n377), .B(new_n772), .C1(new_n773), .C2(G68), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n752), .A2(new_n764), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n428), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT32), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n763), .A2(new_n769), .A3(new_n774), .A4(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n262), .B1(new_n766), .B2(G311), .ZN(new_n779));
  INV_X1    g0579(.A(G322), .ZN(new_n780));
  INV_X1    g0580(.A(new_n768), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n771), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(new_n466), .B2(new_n783), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n759), .B(KEYINPUT90), .Z(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G326), .ZN(new_n787));
  INV_X1    g0587(.A(G283), .ZN(new_n788));
  INV_X1    g0588(.A(G329), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n761), .A2(new_n788), .B1(new_n775), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT91), .ZN(new_n791));
  XNOR2_X1  g0591(.A(KEYINPUT33), .B(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n773), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n784), .A2(new_n787), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G303), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n756), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n778), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n737), .B1(new_n797), .B2(new_n749), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n742), .A2(new_n751), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n738), .A2(new_n799), .ZN(G396));
  INV_X1    g0600(.A(G294), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n781), .A2(new_n801), .B1(new_n217), .B2(new_n765), .ZN(new_n802));
  INV_X1    g0602(.A(new_n775), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n772), .B(new_n802), .C1(G311), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n756), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n262), .B1(new_n805), .B2(G107), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n806), .A2(KEYINPUT93), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT92), .B(G283), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n773), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n795), .B2(new_n759), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(G87), .B2(new_n762), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n806), .A2(KEYINPUT93), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n804), .A2(new_n807), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n773), .A2(G150), .B1(new_n768), .B2(G143), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n815), .B2(new_n759), .C1(new_n428), .C2(new_n765), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n818), .B1(new_n202), .B2(new_n771), .C1(new_n203), .C2(new_n761), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n377), .B1(new_n803), .B2(G132), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n820), .B1(new_n201), .B2(new_n756), .C1(new_n816), .C2(new_n817), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n813), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n737), .B1(new_n822), .B2(new_n749), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n749), .A2(new_n739), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n399), .A2(new_n664), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n391), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n403), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n394), .A2(new_n402), .A3(new_n395), .A4(new_n826), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n823), .B1(G77), .B2(new_n825), .C1(new_n740), .C2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n701), .B(new_n830), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(new_n727), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(new_n736), .ZN(G384));
  NAND2_X1  g0634(.A1(new_n647), .A2(new_n649), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n587), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n666), .A2(new_n537), .A3(new_n641), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n635), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n830), .B(new_n680), .C1(new_n836), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n403), .A2(new_n664), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n313), .A2(new_n664), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n349), .A2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n284), .A2(new_n250), .A3(G169), .ZN(new_n845));
  INV_X1    g0645(.A(new_n290), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n845), .A2(new_n285), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT95), .ZN(new_n848));
  INV_X1    g0648(.A(new_n313), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT95), .B1(new_n292), .B2(new_n313), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n844), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n314), .A2(new_n680), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n839), .A2(new_n841), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT38), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT37), .ZN(new_n857));
  INV_X1    g0657(.A(new_n662), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n438), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n857), .B1(new_n859), .B2(KEYINPUT96), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT7), .B1(new_n377), .B2(new_n212), .ZN(new_n861));
  NOR4_X1   g0661(.A1(new_n375), .A2(new_n376), .A3(new_n423), .A4(G20), .ZN(new_n862));
  OAI21_X1  g0662(.A(G68), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n421), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n430), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT16), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n427), .A2(new_n419), .A3(new_n430), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n435), .B1(new_n868), .B2(new_n294), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n662), .B1(new_n869), .B2(new_n437), .ZN(new_n870));
  AND4_X1   g0670(.A1(new_n434), .A2(new_n436), .A3(new_n458), .A4(new_n437), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n438), .A2(new_n450), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n860), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT96), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n859), .A3(new_n459), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT18), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n873), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n438), .A2(KEYINPUT18), .A3(new_n450), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n859), .B1(new_n883), .B2(new_n654), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n856), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n870), .B1(new_n453), .B2(new_n461), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n878), .A4(new_n874), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n855), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n883), .A2(new_n858), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT97), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n857), .B1(new_n859), .B2(KEYINPUT98), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n872), .A3(new_n873), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT98), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT37), .B1(new_n870), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n877), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n856), .B1(new_n899), .B2(new_n884), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n887), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT39), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n850), .A2(new_n851), .A3(new_n664), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n887), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT97), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n889), .A2(new_n907), .A3(new_n891), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n893), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n700), .A2(new_n703), .ZN(new_n910));
  INV_X1    g0710(.A(new_n463), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n656), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n909), .B(new_n912), .Z(new_n913));
  INV_X1    g0713(.A(new_n830), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n852), .B2(new_n854), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n888), .A2(new_n915), .A3(new_n726), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n292), .A2(KEYINPUT95), .A3(new_n313), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n843), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n726), .B(new_n830), .C1(new_n920), .C2(new_n853), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n917), .B1(new_n900), .B2(new_n887), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n916), .A2(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n911), .A2(new_n726), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n924), .B(new_n925), .Z(new_n926));
  NOR2_X1   g0726(.A1(new_n926), .A2(new_n670), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n913), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n211), .B2(new_n658), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n618), .A2(new_n619), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT35), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G116), .A3(new_n228), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT94), .Z(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n931), .B2(new_n930), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n420), .A2(G77), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n230), .A2(new_n937), .B1(G50), .B2(new_n203), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(G1), .A3(new_n309), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n929), .A2(new_n936), .A3(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n623), .A2(new_n664), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n693), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n679), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n625), .B1(new_n942), .B2(new_n724), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n680), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n944), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n948), .A2(KEYINPUT99), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(KEYINPUT99), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n563), .A2(new_n680), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n644), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n646), .B2(new_n952), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n648), .A2(new_n664), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n942), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n954), .B(KEYINPUT43), .Z(new_n960));
  OAI221_X1 g0760(.A(new_n956), .B1(new_n677), .B2(new_n959), .C1(new_n951), .C2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n956), .B1(new_n951), .B2(new_n960), .ZN(new_n962));
  INV_X1    g0762(.A(new_n677), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n963), .A3(new_n958), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n688), .B(KEYINPUT41), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n679), .B1(new_n676), .B2(new_n678), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n671), .B(new_n967), .Z(new_n968));
  OR2_X1    g0768(.A1(new_n728), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT101), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n728), .A2(new_n970), .A3(new_n968), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n683), .A2(KEYINPUT44), .A3(new_n958), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n682), .B2(new_n959), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n683), .A2(KEYINPUT45), .A3(new_n958), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n682), .B2(new_n959), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(new_n677), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT100), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n677), .B1(new_n976), .B2(new_n980), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n971), .B(new_n972), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n966), .B1(new_n986), .B2(new_n729), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n961), .B(new_n964), .C1(new_n987), .C2(new_n735), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n262), .B1(new_n775), .B2(new_n815), .C1(new_n298), .C2(new_n761), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n783), .A2(G68), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n201), .B2(new_n765), .C1(new_n781), .C2(new_n330), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n989), .B(new_n991), .C1(G58), .C2(new_n805), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n786), .A2(G143), .ZN(new_n993));
  INV_X1    g0793(.A(new_n773), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n992), .B(new_n993), .C1(new_n428), .C2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT104), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT102), .B1(new_n805), .B2(G116), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT46), .Z(new_n998));
  INV_X1    g0798(.A(G311), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n785), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n762), .A2(G97), .ZN(new_n1001));
  INV_X1    g0801(.A(G317), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n377), .C1(new_n1002), .C2(new_n775), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT103), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1003), .A2(new_n1004), .B1(new_n466), .B2(new_n773), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n783), .A2(new_n374), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n768), .A2(new_n533), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n766), .A2(new_n808), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n998), .A2(new_n1000), .A3(new_n1005), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n996), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT47), .Z(new_n1013));
  AND2_X1   g0813(.A1(new_n1013), .A2(new_n749), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n743), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n750), .B1(new_n213), .B2(new_n359), .C1(new_n240), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n741), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n736), .B(new_n1016), .C1(new_n954), .C2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n988), .A2(new_n1020), .ZN(G387));
  INV_X1    g0821(.A(new_n688), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n728), .B2(new_n968), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n969), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n766), .A2(new_n533), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n773), .A2(G311), .B1(new_n768), .B2(G317), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n785), .C2(new_n780), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n783), .A2(new_n808), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n805), .A2(new_n466), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT107), .Z(new_n1032));
  AND2_X1   g0832(.A1(new_n1032), .A2(KEYINPUT49), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1032), .A2(KEYINPUT49), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n803), .A2(G326), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n377), .B1(new_n761), .B2(new_n217), .ZN(new_n1036));
  NOR4_X1   g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n805), .A2(G77), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n331), .B2(new_n994), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n759), .A2(new_n428), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n765), .A2(new_n203), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n768), .A2(G50), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n582), .A2(new_n783), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(KEYINPUT106), .B(G150), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n377), .B1(new_n803), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1001), .A4(new_n1045), .ZN(new_n1046));
  NOR4_X1   g0846(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n749), .B1(new_n1037), .B2(new_n1047), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n331), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1049));
  OAI21_X1  g0849(.A(KEYINPUT50), .B1(new_n331), .B2(G50), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n469), .A3(new_n1050), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n1051), .B(new_n686), .C1(G68), .C2(G77), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n237), .A2(new_n745), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT105), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n743), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n686), .A2(new_n213), .A3(new_n262), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n213), .A2(G107), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n750), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n674), .A2(new_n675), .A3(new_n741), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1048), .A2(new_n736), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1024), .B(new_n1061), .C1(new_n734), .C2(new_n968), .ZN(G393));
  INV_X1    g0862(.A(new_n983), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n981), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n969), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n986), .A2(new_n688), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n735), .A3(new_n981), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n771), .A2(new_n298), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n377), .B(new_n1068), .C1(G143), .C2(new_n803), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1069), .B1(new_n548), .B2(new_n761), .C1(new_n331), .C2(new_n765), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G68), .B2(new_n805), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n781), .A2(new_n428), .B1(new_n330), .B2(new_n759), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1071), .B(new_n1073), .C1(new_n201), .C2(new_n994), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT108), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n783), .A2(G116), .B1(new_n762), .B2(G107), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n262), .B1(new_n803), .B2(G322), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n765), .C2(new_n801), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n533), .B2(new_n773), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n781), .A2(new_n999), .B1(new_n1002), .B2(new_n759), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT52), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n805), .A2(new_n808), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1075), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n737), .B1(new_n1086), .B2(new_n749), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n750), .B1(new_n206), .B2(new_n213), .C1(new_n248), .C2(new_n1015), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n1017), .C2(new_n958), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n1067), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1066), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT109), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1066), .A2(KEYINPUT109), .A3(new_n1090), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(G390));
  INV_X1    g0895(.A(KEYINPUT110), .ZN(new_n1096));
  AND4_X1   g0896(.A1(G330), .A2(new_n405), .A3(new_n462), .A4(new_n726), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(new_n912), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n840), .B1(new_n701), .B2(new_n830), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n726), .A2(G330), .A3(new_n830), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n920), .A2(new_n853), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1100), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT86), .B1(new_n695), .B2(new_n680), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n697), .B(new_n664), .C1(new_n694), .C2(new_n650), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n830), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n841), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1105), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n463), .B1(new_n700), .B2(new_n703), .ZN(new_n1113));
  NOR4_X1   g0913(.A1(new_n1113), .A2(KEYINPUT110), .A3(new_n1097), .A4(new_n656), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1099), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1103), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n904), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n901), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n852), .A2(new_n854), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1118), .B1(new_n1109), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n839), .A2(new_n841), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n904), .B1(new_n1121), .B2(new_n1119), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n903), .B2(new_n905), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n905), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT39), .B1(new_n900), .B2(new_n887), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1125), .A2(new_n1126), .B1(new_n904), .B2(new_n855), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1102), .B1(new_n1108), .B2(new_n841), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1127), .B(new_n1103), .C1(new_n1128), .C2(new_n1118), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1022), .B1(new_n1115), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1099), .A2(new_n1114), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1112), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1130), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1131), .A2(new_n735), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n739), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n805), .A2(new_n1044), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT53), .Z(new_n1141));
  OAI21_X1  g0941(.A(new_n262), .B1(new_n761), .B2(new_n201), .ZN(new_n1142));
  INV_X1    g0942(.A(G132), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT54), .B(G143), .Z(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT111), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n781), .A2(new_n1143), .B1(new_n1145), .B2(new_n765), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1142), .B(new_n1146), .C1(G159), .C2(new_n783), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n803), .A2(G125), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n759), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G128), .A2(new_n1149), .B1(new_n773), .B2(G137), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1141), .A2(new_n1147), .A3(new_n1148), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n759), .A2(new_n788), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n781), .A2(new_n217), .B1(new_n206), .B2(new_n765), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(new_n1068), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n377), .B1(new_n775), .B2(new_n801), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G68), .B2(new_n762), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n805), .A2(G87), .B1(new_n374), .B2(new_n773), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1151), .B1(new_n1152), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n737), .B1(new_n1159), .B2(new_n749), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1139), .B(new_n1160), .C1(new_n364), .C2(new_n825), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1137), .A2(new_n1138), .A3(new_n1161), .ZN(G378));
  INV_X1    g0962(.A(KEYINPUT55), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n417), .B2(new_n340), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n340), .ZN(new_n1165));
  AOI211_X1 g0965(.A(KEYINPUT55), .B(new_n1165), .C1(new_n413), .C2(new_n416), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1164), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n337), .A2(new_n858), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT56), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1169), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n924), .B2(G330), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n885), .A2(new_n887), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n917), .B1(new_n1175), .B2(new_n921), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n922), .A2(new_n923), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1170), .A2(KEYINPUT114), .A3(new_n1172), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT114), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AND4_X1   g0980(.A1(G330), .A2(new_n1176), .A3(new_n1177), .A4(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n909), .B1(new_n1174), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n921), .B1(new_n887), .B2(new_n885), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1177), .B(G330), .C1(new_n1183), .C2(KEYINPUT40), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1173), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n907), .B1(new_n889), .B2(new_n891), .ZN(new_n1187));
  AOI211_X1 g0987(.A(KEYINPUT97), .B(new_n890), .C1(new_n855), .C2(new_n888), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1176), .A2(new_n1180), .A3(G330), .A4(new_n1177), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1186), .A2(new_n1189), .A3(new_n906), .A4(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1182), .A2(KEYINPUT115), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT115), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n909), .C1(new_n1174), .C2(new_n1181), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1133), .B1(new_n1130), .B2(new_n1112), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1197), .B1(new_n1182), .B2(new_n1191), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1022), .B1(new_n1199), .B2(new_n1195), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1192), .A2(new_n735), .A3(new_n1194), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n773), .A2(G97), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1149), .A2(G116), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1038), .A2(new_n990), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n768), .A2(G107), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT112), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n262), .B1(new_n803), .B2(G283), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1208), .B1(new_n202), .B2(new_n761), .C1(new_n765), .C2(new_n359), .ZN(new_n1209));
  NOR4_X1   g1009(.A1(new_n1205), .A2(new_n1207), .A3(G41), .A4(new_n1209), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT58), .Z(new_n1211));
  OAI21_X1  g1011(.A(new_n201), .B1(new_n375), .B2(G41), .ZN(new_n1212));
  AOI21_X1  g1012(.A(G33), .B1(new_n803), .B2(G124), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1213), .B(new_n251), .C1(new_n428), .C2(new_n761), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n994), .A2(new_n1143), .B1(new_n756), .B2(new_n1145), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G137), .A2(new_n766), .B1(new_n768), .B2(G128), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n330), .B2(new_n771), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G125), .C2(new_n1149), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(KEYINPUT113), .B(KEYINPUT59), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1218), .B(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1211), .B(new_n1212), .C1(new_n1214), .C2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n737), .B1(new_n1221), .B2(new_n749), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(G50), .B2(new_n825), .C1(new_n1180), .C2(new_n740), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1202), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1201), .A2(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT116), .Z(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(G375));
  OAI22_X1  g1027(.A1(new_n994), .A2(new_n217), .B1(new_n801), .B2(new_n759), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n766), .A2(new_n374), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n768), .A2(G283), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n377), .B1(new_n775), .B2(new_n795), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G77), .B2(new_n762), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1232), .A4(new_n1043), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1228), .B(new_n1233), .C1(G97), .C2(new_n805), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n768), .A2(G137), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1235), .B1(new_n1143), .B2(new_n759), .C1(new_n994), .C2(new_n1145), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT117), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n262), .B1(new_n761), .B2(new_n202), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT118), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n756), .A2(new_n428), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n765), .A2(new_n330), .B1(new_n201), .B2(new_n771), .ZN(new_n1242));
  NOR4_X1   g1042(.A1(new_n1237), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n803), .A2(G128), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1234), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT119), .Z(new_n1246));
  AOI21_X1  g1046(.A(new_n737), .B1(new_n1246), .B2(new_n749), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n740), .B2(new_n1119), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n203), .B2(new_n824), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(new_n1134), .B2(new_n735), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1112), .B1(new_n1099), .B2(new_n1114), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n965), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1250), .B1(new_n1252), .B2(new_n1115), .ZN(G381));
  NOR2_X1   g1053(.A1(G375), .A2(G378), .ZN(new_n1254));
  AND4_X1   g1054(.A1(new_n1020), .A2(new_n1093), .A3(new_n988), .A4(new_n1094), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(G393), .A2(G396), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(G381), .A2(G384), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(G407));
  NAND2_X1  g1058(.A1(new_n1138), .A2(new_n1161), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1226), .A2(G213), .A3(new_n663), .A4(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT120), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(G407), .A2(new_n1263), .A3(G213), .A4(new_n1264), .ZN(G409));
  NAND3_X1  g1065(.A1(new_n1201), .A2(G378), .A3(new_n1224), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1182), .A2(new_n1191), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n735), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1223), .B(new_n1268), .C1(new_n1196), .C2(new_n966), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1260), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT121), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n663), .A2(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT60), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1251), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1135), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n688), .B1(new_n1251), .B2(new_n1275), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1250), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G384), .A2(KEYINPUT122), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G384), .B(KEYINPUT122), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1250), .B(new_n1282), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1266), .A2(new_n1270), .A3(KEYINPUT121), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1273), .A2(new_n1274), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AND4_X1   g1089(.A1(KEYINPUT62), .A2(new_n1271), .A3(new_n1274), .A4(new_n1285), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1295));
  AND3_X1   g1095(.A1(new_n663), .A2(G213), .A3(G2897), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1284), .B(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1292), .A2(new_n1293), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n964), .A2(new_n961), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n986), .A2(new_n729), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n965), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1301), .B1(new_n1303), .B2(new_n734), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1094), .ZN(new_n1305));
  AOI21_X1  g1105(.A(KEYINPUT109), .B1(new_n1066), .B2(new_n1090), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n1304), .A2(new_n1019), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1093), .A2(new_n988), .A3(new_n1020), .A4(new_n1094), .ZN(new_n1308));
  AND2_X1   g1108(.A1(G393), .A2(G396), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT123), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1309), .A2(new_n1256), .A3(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1310), .B1(new_n1309), .B2(new_n1256), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AND3_X1   g1114(.A1(new_n1307), .A2(new_n1308), .A3(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1311), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1315), .A2(new_n1316), .A3(KEYINPUT126), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT126), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1093), .A2(new_n1094), .B1(new_n988), .B2(new_n1020), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1312), .B1(new_n1255), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1307), .A2(new_n1314), .A3(new_n1308), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1318), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1317), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1290), .B1(new_n1287), .B2(new_n1288), .ZN(new_n1324));
  OAI21_X1  g1124(.A(KEYINPUT125), .B1(new_n1324), .B2(new_n1298), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1300), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1295), .A2(KEYINPUT63), .A3(new_n1285), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1273), .A2(new_n1274), .A3(new_n1286), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1297), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1329), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1287), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1327), .B(new_n1328), .C1(new_n1332), .C2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1326), .A2(new_n1334), .ZN(G405));
  OAI21_X1  g1135(.A(KEYINPUT126), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1320), .A2(new_n1321), .A3(new_n1318), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1284), .A2(KEYINPUT127), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1336), .A2(new_n1337), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1339), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1266), .B1(new_n1226), .B2(G378), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1340), .A2(new_n1341), .A3(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1342), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1338), .B1(new_n1317), .B2(new_n1322), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1336), .A2(new_n1337), .A3(new_n1339), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1344), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1343), .A2(new_n1347), .ZN(G402));
endmodule


