

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589;

  XNOR2_X1 U321 ( .A(n460), .B(n459), .ZN(n545) );
  XNOR2_X1 U322 ( .A(n393), .B(n392), .ZN(n570) );
  XNOR2_X1 U323 ( .A(n391), .B(KEYINPUT121), .ZN(n392) );
  XNOR2_X1 U324 ( .A(n478), .B(n477), .ZN(n503) );
  XOR2_X1 U325 ( .A(KEYINPUT93), .B(n465), .Z(n569) );
  XOR2_X1 U326 ( .A(G36GAT), .B(G218GAT), .Z(n289) );
  NAND2_X1 U327 ( .A1(n569), .A2(n469), .ZN(n290) );
  XNOR2_X1 U328 ( .A(n325), .B(KEYINPUT111), .ZN(n326) );
  XNOR2_X1 U329 ( .A(n327), .B(n326), .ZN(n343) );
  XNOR2_X1 U330 ( .A(KEYINPUT98), .B(KEYINPUT97), .ZN(n456) );
  XNOR2_X1 U331 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U332 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U333 ( .A(n423), .B(n422), .ZN(n428) );
  XOR2_X1 U334 ( .A(G197GAT), .B(KEYINPUT21), .Z(n419) );
  XNOR2_X1 U335 ( .A(KEYINPUT26), .B(KEYINPUT95), .ZN(n459) );
  XNOR2_X1 U336 ( .A(n419), .B(n289), .ZN(n386) );
  XNOR2_X1 U337 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U338 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U339 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U340 ( .A(KEYINPUT38), .B(KEYINPUT106), .ZN(n477) );
  INV_X1 U341 ( .A(G43GAT), .ZN(n479) );
  XNOR2_X1 U342 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U343 ( .A(n479), .B(KEYINPUT40), .ZN(n480) );
  XNOR2_X1 U344 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  INV_X1 U346 ( .A(KEYINPUT112), .ZN(n345) );
  XOR2_X1 U347 ( .A(KEYINPUT71), .B(KEYINPUT73), .Z(n292) );
  XNOR2_X1 U348 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n291) );
  XNOR2_X1 U349 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U350 ( .A(G43GAT), .B(G50GAT), .Z(n294) );
  XOR2_X1 U351 ( .A(G15GAT), .B(G22GAT), .Z(n333) );
  XNOR2_X1 U352 ( .A(n333), .B(KEYINPUT68), .ZN(n293) );
  XNOR2_X1 U353 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U354 ( .A(n296), .B(n295), .Z(n298) );
  NAND2_X1 U355 ( .A1(G229GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U356 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U357 ( .A(G141GAT), .B(G197GAT), .Z(n300) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G113GAT), .ZN(n299) );
  XNOR2_X1 U359 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U360 ( .A(n302), .B(n301), .Z(n310) );
  XOR2_X1 U361 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n304) );
  XNOR2_X1 U362 ( .A(G36GAT), .B(G29GAT), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U364 ( .A(KEYINPUT72), .B(n305), .Z(n365) );
  XOR2_X1 U365 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n307) );
  XNOR2_X1 U366 ( .A(G1GAT), .B(G8GAT), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n365), .B(n308), .ZN(n309) );
  XOR2_X1 U369 ( .A(n310), .B(n309), .Z(n505) );
  INV_X1 U370 ( .A(n505), .ZN(n574) );
  XOR2_X1 U371 ( .A(G106GAT), .B(G78GAT), .Z(n418) );
  XOR2_X1 U372 ( .A(G99GAT), .B(G85GAT), .Z(n361) );
  XNOR2_X1 U373 ( .A(n418), .B(n361), .ZN(n324) );
  XOR2_X1 U374 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n312) );
  NAND2_X1 U375 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U377 ( .A(n313), .B(KEYINPUT33), .Z(n318) );
  XOR2_X1 U378 ( .A(G64GAT), .B(KEYINPUT75), .Z(n315) );
  XNOR2_X1 U379 ( .A(G204GAT), .B(G92GAT), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n315), .B(n314), .ZN(n381) );
  XNOR2_X1 U381 ( .A(G71GAT), .B(G57GAT), .ZN(n316) );
  XOR2_X1 U382 ( .A(n316), .B(KEYINPUT13), .Z(n341) );
  XOR2_X1 U383 ( .A(n381), .B(n341), .Z(n317) );
  XNOR2_X1 U384 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U385 ( .A(G120GAT), .B(G148GAT), .Z(n408) );
  XNOR2_X1 U386 ( .A(G176GAT), .B(n408), .ZN(n320) );
  INV_X1 U387 ( .A(KEYINPUT32), .ZN(n319) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n578) );
  XNOR2_X1 U389 ( .A(KEYINPUT41), .B(n578), .ZN(n559) );
  NOR2_X1 U390 ( .A1(n574), .A2(n559), .ZN(n327) );
  INV_X1 U391 ( .A(KEYINPUT46), .ZN(n325) );
  XOR2_X1 U392 ( .A(G211GAT), .B(KEYINPUT81), .Z(n329) );
  XNOR2_X1 U393 ( .A(G8GAT), .B(G183GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n383) );
  XOR2_X1 U395 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n331) );
  XNOR2_X1 U396 ( .A(G78GAT), .B(G64GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U398 ( .A(n333), .B(n332), .Z(n335) );
  NAND2_X1 U399 ( .A1(G231GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U401 ( .A(n336), .B(KEYINPUT15), .Z(n339) );
  XNOR2_X1 U402 ( .A(G1GAT), .B(G127GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n337), .B(G155GAT), .ZN(n410) );
  XNOR2_X1 U404 ( .A(n410), .B(KEYINPUT82), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U406 ( .A(n383), .B(n340), .ZN(n342) );
  XOR2_X1 U407 ( .A(n342), .B(n341), .Z(n552) );
  XOR2_X1 U408 ( .A(KEYINPUT110), .B(n552), .Z(n564) );
  NOR2_X1 U409 ( .A1(n343), .A2(n564), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n366) );
  XOR2_X1 U411 ( .A(KEYINPUT64), .B(KEYINPUT79), .Z(n347) );
  XNOR2_X1 U412 ( .A(KEYINPUT67), .B(KEYINPUT80), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U414 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n349) );
  XNOR2_X1 U415 ( .A(G190GAT), .B(G162GAT), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U417 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U418 ( .A(G50GAT), .B(G218GAT), .Z(n417) );
  XOR2_X1 U419 ( .A(G92GAT), .B(G106GAT), .Z(n353) );
  NAND2_X1 U420 ( .A1(G232GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n417), .B(n354), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT66), .B(KEYINPUT9), .Z(n358) );
  XNOR2_X1 U425 ( .A(KEYINPUT77), .B(KEYINPUT10), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U427 ( .A(n360), .B(n359), .Z(n363) );
  XOR2_X1 U428 ( .A(G43GAT), .B(G134GAT), .Z(n437) );
  XNOR2_X1 U429 ( .A(n437), .B(n361), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U431 ( .A(n365), .B(n364), .Z(n555) );
  INV_X1 U432 ( .A(n555), .ZN(n540) );
  NOR2_X1 U433 ( .A1(n366), .A2(n540), .ZN(n367) );
  XNOR2_X1 U434 ( .A(KEYINPUT47), .B(n367), .ZN(n375) );
  XOR2_X1 U435 ( .A(KEYINPUT36), .B(n555), .Z(n584) );
  INV_X1 U436 ( .A(n552), .ZN(n581) );
  NAND2_X1 U437 ( .A1(n584), .A2(n581), .ZN(n370) );
  XOR2_X1 U438 ( .A(KEYINPUT113), .B(KEYINPUT45), .Z(n368) );
  XNOR2_X1 U439 ( .A(KEYINPUT65), .B(n368), .ZN(n369) );
  XNOR2_X1 U440 ( .A(n370), .B(n369), .ZN(n371) );
  NAND2_X1 U441 ( .A1(n371), .A2(n574), .ZN(n372) );
  NOR2_X1 U442 ( .A1(n578), .A2(n372), .ZN(n373) );
  XOR2_X1 U443 ( .A(KEYINPUT114), .B(n373), .Z(n374) );
  NAND2_X1 U444 ( .A1(n375), .A2(n374), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n376), .B(KEYINPUT48), .ZN(n526) );
  XOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n378) );
  XNOR2_X1 U447 ( .A(G169GAT), .B(G176GAT), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n378), .B(n377), .ZN(n380) );
  XOR2_X1 U449 ( .A(G190GAT), .B(KEYINPUT19), .Z(n379) );
  XOR2_X1 U450 ( .A(n380), .B(n379), .Z(n447) );
  INV_X1 U451 ( .A(n447), .ZN(n382) );
  XOR2_X1 U452 ( .A(n382), .B(n381), .Z(n389) );
  XNOR2_X1 U453 ( .A(KEYINPUT94), .B(n383), .ZN(n385) );
  AND2_X1 U454 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U455 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U456 ( .A(n389), .B(n388), .Z(n390) );
  INV_X1 U457 ( .A(n390), .ZN(n454) );
  NAND2_X1 U458 ( .A1(n526), .A2(n454), .ZN(n393) );
  XOR2_X1 U459 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n391) );
  XOR2_X1 U460 ( .A(KEYINPUT2), .B(G162GAT), .Z(n395) );
  XNOR2_X1 U461 ( .A(KEYINPUT3), .B(KEYINPUT87), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U463 ( .A(G141GAT), .B(n396), .Z(n432) );
  XOR2_X1 U464 ( .A(KEYINPUT91), .B(G85GAT), .Z(n398) );
  XNOR2_X1 U465 ( .A(G29GAT), .B(G134GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U467 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n400) );
  XNOR2_X1 U468 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U470 ( .A(n402), .B(n401), .Z(n407) );
  XOR2_X1 U471 ( .A(KEYINPUT90), .B(G57GAT), .Z(n404) );
  NAND2_X1 U472 ( .A1(G225GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U474 ( .A(KEYINPUT92), .B(n405), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n409) );
  XOR2_X1 U476 ( .A(n409), .B(n408), .Z(n412) );
  XOR2_X1 U477 ( .A(G113GAT), .B(KEYINPUT0), .Z(n434) );
  XNOR2_X1 U478 ( .A(n434), .B(n410), .ZN(n411) );
  XNOR2_X1 U479 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n432), .B(n413), .ZN(n465) );
  XOR2_X1 U481 ( .A(G22GAT), .B(G148GAT), .Z(n415) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U486 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n421) );
  INV_X1 U487 ( .A(KEYINPUT24), .ZN(n420) );
  XOR2_X1 U488 ( .A(G155GAT), .B(G204GAT), .Z(n425) );
  XNOR2_X1 U489 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n424) );
  XNOR2_X1 U490 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U491 ( .A(n426), .B(KEYINPUT88), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n469) );
  OR2_X1 U495 ( .A1(n570), .A2(n290), .ZN(n433) );
  XNOR2_X1 U496 ( .A(n433), .B(KEYINPUT55), .ZN(n449) );
  XOR2_X1 U497 ( .A(n434), .B(G71GAT), .Z(n436) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U500 ( .A(n438), .B(n437), .Z(n446) );
  XOR2_X1 U501 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n440) );
  XNOR2_X1 U502 ( .A(G99GAT), .B(G183GAT), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U504 ( .A(G120GAT), .B(G127GAT), .Z(n442) );
  XNOR2_X1 U505 ( .A(G15GAT), .B(KEYINPUT85), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U507 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U508 ( .A(n446), .B(n445), .Z(n448) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n529) );
  NAND2_X1 U510 ( .A1(n449), .A2(n529), .ZN(n560) );
  INV_X1 U511 ( .A(n560), .ZN(n565) );
  NAND2_X1 U512 ( .A1(n565), .A2(n540), .ZN(n452) );
  XOR2_X1 U513 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n450) );
  INV_X1 U514 ( .A(n529), .ZN(n521) );
  NOR2_X1 U515 ( .A1(n578), .A2(n574), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n453), .B(KEYINPUT76), .ZN(n492) );
  NAND2_X1 U517 ( .A1(n454), .A2(n529), .ZN(n455) );
  NAND2_X1 U518 ( .A1(n455), .A2(n469), .ZN(n457) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT25), .ZN(n464) );
  INV_X1 U520 ( .A(KEYINPUT96), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n390), .B(KEYINPUT27), .ZN(n468) );
  NOR2_X1 U522 ( .A1(n529), .A2(n469), .ZN(n460) );
  NOR2_X1 U523 ( .A1(n468), .A2(n545), .ZN(n461) );
  XNOR2_X1 U524 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U525 ( .A1(n464), .A2(n463), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT99), .ZN(n473) );
  XOR2_X1 U528 ( .A(n521), .B(KEYINPUT86), .Z(n471) );
  NOR2_X1 U529 ( .A1(n468), .A2(n569), .ZN(n527) );
  XNOR2_X1 U530 ( .A(KEYINPUT28), .B(n469), .ZN(n532) );
  NAND2_X1 U531 ( .A1(n527), .A2(n532), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT100), .B(n474), .Z(n490) );
  AND2_X1 U535 ( .A1(n584), .A2(n552), .ZN(n475) );
  AND2_X1 U536 ( .A1(n490), .A2(n475), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT37), .B(n476), .Z(n517) );
  NAND2_X1 U538 ( .A1(n492), .A2(n517), .ZN(n478) );
  NOR2_X1 U539 ( .A1(n521), .A2(n503), .ZN(n481) );
  NOR2_X1 U540 ( .A1(n569), .A2(n503), .ZN(n485) );
  XNOR2_X1 U541 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n483) );
  INV_X1 U542 ( .A(G29GAT), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(G1328GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT102), .B(KEYINPUT34), .Z(n487) );
  XNOR2_X1 U546 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n494) );
  NAND2_X1 U548 ( .A1(n581), .A2(n555), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(KEYINPUT83), .ZN(n489) );
  XNOR2_X1 U550 ( .A(KEYINPUT16), .B(n489), .ZN(n491) );
  AND2_X1 U551 ( .A1(n491), .A2(n490), .ZN(n507) );
  NAND2_X1 U552 ( .A1(n507), .A2(n492), .ZN(n500) );
  NOR2_X1 U553 ( .A1(n569), .A2(n500), .ZN(n493) );
  XOR2_X1 U554 ( .A(n494), .B(n493), .Z(G1324GAT) );
  NOR2_X1 U555 ( .A1(n390), .A2(n500), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1325GAT) );
  NOR2_X1 U558 ( .A1(n521), .A2(n500), .ZN(n498) );
  XNOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G15GAT), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U562 ( .A1(n532), .A2(n500), .ZN(n501) );
  XOR2_X1 U563 ( .A(G22GAT), .B(n501), .Z(G1327GAT) );
  NOR2_X1 U564 ( .A1(n503), .A2(n390), .ZN(n502) );
  XOR2_X1 U565 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U566 ( .A1(n532), .A2(n503), .ZN(n504) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  NOR2_X1 U568 ( .A1(n559), .A2(n505), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n506), .B(KEYINPUT108), .ZN(n516) );
  NAND2_X1 U570 ( .A1(n507), .A2(n516), .ZN(n513) );
  NOR2_X1 U571 ( .A1(n569), .A2(n513), .ZN(n509) );
  XNOR2_X1 U572 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n390), .A2(n513), .ZN(n511) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n521), .A2(n513), .ZN(n512) );
  XOR2_X1 U578 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U579 ( .A1(n532), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U582 ( .A1(n517), .A2(n516), .ZN(n523) );
  NOR2_X1 U583 ( .A1(n569), .A2(n523), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NOR2_X1 U586 ( .A1(n390), .A2(n523), .ZN(n520) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n523), .ZN(n522) );
  XOR2_X1 U589 ( .A(G99GAT), .B(n522), .Z(G1338GAT) );
  NOR2_X1 U590 ( .A1(n532), .A2(n523), .ZN(n524) );
  XOR2_X1 U591 ( .A(KEYINPUT44), .B(n524), .Z(n525) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  NAND2_X1 U593 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(KEYINPUT115), .ZN(n546) );
  NAND2_X1 U595 ( .A1(n529), .A2(n546), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(n530), .Z(n531) );
  NAND2_X1 U597 ( .A1(n532), .A2(n531), .ZN(n537) );
  NOR2_X1 U598 ( .A1(n574), .A2(n537), .ZN(n533) );
  XOR2_X1 U599 ( .A(G113GAT), .B(n533), .Z(G1340GAT) );
  NOR2_X1 U600 ( .A1(n559), .A2(n537), .ZN(n535) );
  XNOR2_X1 U601 ( .A(KEYINPUT49), .B(KEYINPUT117), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U603 ( .A(G120GAT), .B(n536), .Z(G1341GAT) );
  INV_X1 U604 ( .A(n537), .ZN(n541) );
  NAND2_X1 U605 ( .A1(n541), .A2(n564), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n538), .B(KEYINPUT50), .ZN(n539) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U609 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  INV_X1 U612 ( .A(n545), .ZN(n572) );
  NAND2_X1 U613 ( .A1(n572), .A2(n546), .ZN(n547) );
  XOR2_X1 U614 ( .A(KEYINPUT119), .B(n547), .Z(n554) );
  NOR2_X1 U615 ( .A1(n574), .A2(n554), .ZN(n548) );
  XOR2_X1 U616 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  NOR2_X1 U617 ( .A1(n559), .A2(n554), .ZN(n550) );
  XNOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NOR2_X1 U621 ( .A1(n552), .A2(n554), .ZN(n553) );
  XOR2_X1 U622 ( .A(G155GAT), .B(n553), .Z(G1346GAT) );
  NOR2_X1 U623 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U624 ( .A(G162GAT), .B(n556), .Z(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT120), .B(n557), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n574), .ZN(n558) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n558), .Z(G1348GAT) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n576) );
  INV_X1 U637 ( .A(n569), .ZN(n571) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n577) );
  NOR2_X1 U640 ( .A1(n574), .A2(n577), .ZN(n575) );
  XOR2_X1 U641 ( .A(n576), .B(n575), .Z(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  INV_X1 U643 ( .A(n577), .ZN(n585) );
  NAND2_X1 U644 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  XOR2_X1 U646 ( .A(G211GAT), .B(KEYINPUT125), .Z(n583) );
  NAND2_X1 U647 ( .A1(n585), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n589) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(G1355GAT) );
endmodule

