//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n989, new_n990;
  XNOR2_X1  g000(.A(KEYINPUT14), .B(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT14), .ZN(new_n205));
  NOR3_X1   g004(.A1(new_n205), .A2(new_n203), .A3(G29gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT15), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT84), .ZN(new_n209));
  INV_X1    g008(.A(G43gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G50gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n204), .A2(new_n207), .B1(new_n208), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n208), .ZN(new_n215));
  INV_X1    g014(.A(G29gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n218));
  AOI21_X1  g017(.A(G36gat), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n215), .B(new_n213), .C1(new_n219), .C2(new_n206), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n208), .A3(new_n207), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n214), .A2(KEYINPUT17), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n212), .B2(new_n213), .ZN(new_n224));
  INV_X1    g023(.A(new_n220), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G15gat), .B(G22gat), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n228), .A2(G1gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT16), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n230), .B2(G1gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(KEYINPUT85), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G8gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n228), .A2(G1gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT85), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT86), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n239), .A3(new_n236), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n229), .A2(new_n233), .A3(new_n231), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT87), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT87), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n229), .A2(new_n243), .A3(new_n233), .A4(new_n231), .ZN(new_n244));
  AOI22_X1  g043(.A1(new_n238), .A2(new_n240), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(G229gat), .A2(G233gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n242), .A2(new_n244), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n232), .A2(new_n239), .A3(new_n236), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n239), .B1(new_n232), .B2(new_n236), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n224), .A2(new_n225), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n246), .A2(new_n247), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT18), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n251), .B(new_n252), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n247), .B(KEYINPUT13), .Z(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n246), .A2(KEYINPUT18), .A3(new_n247), .A4(new_n253), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G141gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT83), .B(G197gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT11), .B(G169gat), .Z(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT12), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n256), .A2(new_n259), .A3(new_n260), .A4(new_n267), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G99gat), .B(G106gat), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n273), .A2(KEYINPUT92), .ZN(new_n274));
  NAND3_X1  g073(.A1(KEYINPUT91), .A2(G85gat), .A3(G92gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT7), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g076(.A1(KEYINPUT91), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G99gat), .A2(G106gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT8), .ZN(new_n280));
  INV_X1    g079(.A(G85gat), .ZN(new_n281));
  INV_X1    g080(.A(G92gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n277), .A2(new_n278), .A3(new_n280), .A4(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n273), .A2(KEYINPUT92), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n274), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NOR3_X1   g085(.A1(new_n284), .A2(KEYINPUT92), .A3(new_n273), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n288), .A2(new_n224), .A3(new_n225), .ZN(new_n289));
  AND2_X1   g088(.A1(G232gat), .A2(G233gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(KEYINPUT41), .B2(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n227), .A2(KEYINPUT93), .A3(new_n288), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT93), .B1(new_n227), .B2(new_n288), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G190gat), .B(G218gat), .Z(new_n295));
  OR2_X1    g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n290), .A2(KEYINPUT41), .ZN(new_n297));
  XNOR2_X1  g096(.A(G134gat), .B(G162gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n295), .ZN(new_n300));
  AND3_X1   g099(.A1(new_n296), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n296), .B2(new_n300), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(KEYINPUT88), .A2(G64gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(KEYINPUT88), .A2(G64gat), .ZN(new_n307));
  OAI21_X1  g106(.A(G57gat), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n309));
  INV_X1    g108(.A(G57gat), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n310), .B2(G64gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G71gat), .A2(G78gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT9), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(KEYINPUT90), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n314), .ZN(new_n317));
  INV_X1    g116(.A(G71gat), .ZN(new_n318));
  INV_X1    g117(.A(G78gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n316), .A2(new_n317), .B1(new_n320), .B2(new_n313), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n309), .B(G57gat), .C1(new_n306), .C2(new_n307), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n312), .A2(new_n315), .A3(new_n321), .A4(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G57gat), .B(G64gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n313), .B(new_n320), .C1(new_n324), .C2(new_n314), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT21), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G231gat), .A2(G233gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G127gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n245), .B1(new_n327), .B2(new_n326), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(G183gat), .B(G211gat), .Z(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n339), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n326), .B1(new_n287), .B2(new_n286), .ZN(new_n343));
  NAND2_X1  g142(.A1(G230gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n284), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n273), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n284), .A2(new_n346), .A3(new_n273), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n323), .A3(new_n325), .A4(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n352), .A2(KEYINPUT96), .ZN(new_n353));
  XOR2_X1   g152(.A(KEYINPUT95), .B(KEYINPUT10), .Z(new_n354));
  AOI21_X1  g153(.A(new_n354), .B1(new_n343), .B2(new_n351), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n323), .A2(KEYINPUT10), .A3(new_n325), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n288), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n344), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(KEYINPUT96), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G120gat), .B(G148gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(G176gat), .B(G204gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n353), .A2(new_n358), .A3(new_n363), .A4(new_n359), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n304), .A2(new_n342), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G141gat), .B(G148gat), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT2), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n375), .B1(G155gat), .B2(G162gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n373), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G141gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G148gat), .ZN(new_n379));
  INV_X1    g178(.A(G148gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G141gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G155gat), .B(G162gat), .ZN(new_n383));
  INV_X1    g182(.A(G162gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT2), .B1(new_n335), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n377), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(KEYINPUT75), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n377), .A2(new_n386), .A3(new_n390), .A4(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n386), .ZN(new_n393));
  XOR2_X1   g192(.A(G113gat), .B(G120gat), .Z(new_n394));
  INV_X1    g193(.A(KEYINPUT1), .ZN(new_n395));
  XNOR2_X1  g194(.A(G127gat), .B(G134gat), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(G127gat), .B(G134gat), .Z(new_n398));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(KEYINPUT1), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n393), .A2(KEYINPUT3), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n392), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n400), .A2(new_n397), .A3(new_n377), .A4(new_n386), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n370), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT39), .ZN(new_n408));
  INV_X1    g207(.A(new_n393), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n400), .A2(new_n397), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n409), .B(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n411), .B2(new_n369), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n404), .B(KEYINPUT4), .ZN(new_n414));
  AOI211_X1 g213(.A(KEYINPUT39), .B(new_n369), .C1(new_n414), .C2(new_n402), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n416));
  XOR2_X1   g215(.A(G1gat), .B(G29gat), .Z(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n415), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n408), .B(new_n370), .C1(new_n403), .C2(new_n406), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT80), .B1(new_n424), .B2(new_n421), .ZN(new_n425));
  OAI211_X1 g224(.A(KEYINPUT40), .B(new_n413), .C1(new_n423), .C2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n416), .B1(new_n415), .B2(new_n422), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n421), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n431), .A2(KEYINPUT81), .A3(KEYINPUT40), .A4(new_n413), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT40), .B1(new_n431), .B2(new_n413), .ZN(new_n434));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n435), .B(KEYINPUT73), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT74), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT27), .B(G183gat), .ZN(new_n440));
  INV_X1    g239(.A(G190gat), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT65), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n443));
  NOR2_X1   g242(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(G183gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT27), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(G183gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n450), .A3(new_n441), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT65), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n445), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT26), .ZN(new_n457));
  NAND2_X1  g256(.A1(G183gat), .A2(G190gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(G169gat), .A2(G176gat), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT26), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n457), .B(new_n458), .C1(new_n461), .C2(new_n456), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n455), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT25), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT24), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n441), .ZN(new_n468));
  NAND3_X1  g267(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G169gat), .ZN(new_n471));
  INV_X1    g270(.A(G176gat), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT23), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G169gat), .B2(G176gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n475), .A3(new_n459), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n465), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  AND4_X1   g276(.A1(KEYINPUT25), .A2(new_n473), .A3(new_n475), .A4(new_n459), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT64), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n458), .B1(new_n479), .B2(KEYINPUT24), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n466), .A2(KEYINPUT64), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n468), .B(new_n469), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G226gat), .A2(G233gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(G197gat), .A2(G204gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(G197gat), .A2(G204gat), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT69), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT70), .ZN(new_n494));
  AND2_X1   g293(.A1(G211gat), .A2(G218gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(G211gat), .A2(G218gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(G211gat), .ZN(new_n498));
  INV_X1    g297(.A(G218gat), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G211gat), .A2(G218gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(KEYINPUT70), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G197gat), .B(G204gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT69), .ZN(new_n505));
  INV_X1    g304(.A(new_n492), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n493), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n500), .A2(new_n501), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n504), .A3(new_n506), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT71), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n493), .A2(new_n503), .A3(new_n512), .A4(new_n507), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT29), .B1(new_n464), .B2(new_n484), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n488), .B(new_n514), .C1(new_n487), .C2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n462), .B1(new_n442), .B2(new_n445), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n518), .A2(new_n455), .B1(new_n477), .B2(new_n483), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n486), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n514), .B1(new_n522), .B2(new_n488), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n439), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n488), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n513), .A2(new_n511), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n437), .B(new_n438), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n529), .A2(new_n516), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(new_n531), .A3(KEYINPUT30), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT5), .B1(new_n411), .B2(new_n369), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n414), .A2(new_n402), .A3(new_n369), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n414), .A2(new_n402), .A3(KEYINPUT5), .A4(new_n369), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n422), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n529), .A2(new_n538), .A3(new_n516), .A4(new_n530), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n532), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n434), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT78), .A2(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G228gat), .ZN(new_n544));
  INV_X1    g343(.A(G233gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n521), .B1(new_n389), .B2(new_n391), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n514), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n526), .B2(new_n527), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n387), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n393), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n495), .A2(new_n496), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n491), .B2(new_n492), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(new_n511), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n393), .A3(new_n520), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT77), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n556), .B2(new_n558), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n392), .A2(new_n520), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n528), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n546), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n543), .B1(new_n552), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G78gat), .B(G106gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G50gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n556), .A2(new_n558), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT77), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n547), .A2(new_n514), .ZN(new_n574));
  OAI22_X1  g373(.A1(new_n573), .A2(new_n574), .B1(new_n544), .B2(new_n545), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT3), .B1(new_n514), .B2(new_n549), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n563), .B(new_n546), .C1(new_n576), .C2(new_n409), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n577), .A3(new_n542), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n565), .A2(new_n569), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT79), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT79), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n565), .A2(new_n581), .A3(new_n578), .A4(new_n569), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G22gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n552), .B2(new_n564), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n575), .A2(new_n577), .A3(G22gat), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n585), .A2(new_n586), .A3(new_n568), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n433), .A2(new_n541), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n529), .A2(new_n590), .A3(new_n516), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT82), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n529), .A2(KEYINPUT82), .A3(new_n590), .A4(new_n516), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT37), .B1(new_n517), .B2(new_n523), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n439), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT38), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n535), .A2(new_n536), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT6), .B1(new_n599), .B2(new_n421), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n537), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n535), .A2(KEYINPUT6), .A3(new_n422), .A4(new_n536), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  MUX2_X1   g403(.A(new_n519), .B(new_n515), .S(new_n486), .Z(new_n605));
  AOI21_X1  g404(.A(new_n590), .B1(new_n605), .B2(new_n528), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n525), .A2(new_n514), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT38), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n595), .A2(new_n439), .A3(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n598), .A2(new_n604), .A3(new_n531), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n532), .A2(new_n539), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n587), .B1(new_n580), .B2(new_n582), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n589), .A2(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n451), .A2(new_n452), .A3(new_n445), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n445), .B1(new_n451), .B2(new_n452), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n615), .A2(new_n616), .A3(new_n462), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n618), .A2(new_n473), .A3(new_n459), .A4(new_n475), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n619), .A2(new_n465), .B1(new_n478), .B2(new_n482), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n410), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n410), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n464), .A2(new_n484), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G227gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT67), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT67), .ZN(new_n628));
  AOI211_X1 g427(.A(new_n628), .B(new_n625), .C1(new_n621), .C2(new_n623), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT32), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n627), .B2(new_n629), .ZN(new_n632));
  XOR2_X1   g431(.A(G15gat), .B(G43gat), .Z(new_n633));
  XNOR2_X1  g432(.A(G71gat), .B(G99gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n630), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n625), .A3(new_n623), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT34), .Z(new_n638));
  INV_X1    g437(.A(new_n635), .ZN(new_n639));
  OAI221_X1 g438(.A(KEYINPUT32), .B1(new_n631), .B2(new_n639), .C1(new_n627), .C2(new_n629), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n638), .B1(new_n636), .B2(new_n640), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT36), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT36), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n636), .A2(new_n640), .ZN(new_n647));
  INV_X1    g446(.A(new_n638), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT68), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n650), .A3(new_n641), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n643), .A2(KEYINPUT68), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n646), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n614), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n601), .A2(new_n602), .B1(new_n539), .B2(new_n532), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n583), .A2(new_n588), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT68), .ZN(new_n657));
  INV_X1    g456(.A(new_n652), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n655), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT35), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT35), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n656), .A2(new_n661), .A3(new_n655), .A4(new_n644), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n272), .B(new_n368), .C1(new_n654), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n604), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g465(.A(KEYINPUT97), .B(KEYINPUT42), .ZN(new_n667));
  INV_X1    g466(.A(new_n611), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT98), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(G8gat), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n672), .B(new_n673), .C1(new_n669), .C2(new_n675), .ZN(G1325gat));
  AOI21_X1  g475(.A(G15gat), .B1(new_n664), .B2(new_n644), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT36), .B1(new_n657), .B2(new_n658), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n649), .A2(new_n641), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n646), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT99), .B1(new_n653), .B2(new_n645), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G15gat), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT100), .Z(new_n686));
  AOI21_X1  g485(.A(new_n677), .B1(new_n686), .B2(new_n664), .ZN(G1326gat));
  NAND2_X1  g486(.A1(new_n664), .A2(new_n613), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  AOI21_X1  g489(.A(new_n272), .B1(new_n654), .B2(new_n663), .ZN(new_n691));
  INV_X1    g490(.A(new_n342), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n367), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n304), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n603), .A2(G29gat), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT102), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT101), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n702), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n656), .B2(new_n655), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n613), .A2(new_n612), .A3(KEYINPUT103), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n708), .A2(new_n709), .B1(new_n589), .B2(new_n610), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n682), .A3(new_n683), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n613), .B1(new_n651), .B2(new_n652), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n661), .B1(new_n713), .B2(new_n655), .ZN(new_n714));
  INV_X1    g513(.A(new_n662), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n660), .A2(new_n662), .A3(KEYINPUT104), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n711), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n303), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n654), .A2(new_n663), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(KEYINPUT44), .A3(new_n303), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n693), .A2(new_n272), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n724), .A2(new_n603), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n727), .A2(KEYINPUT105), .ZN(new_n728));
  OAI21_X1  g527(.A(G29gat), .B1(new_n727), .B2(KEYINPUT105), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n705), .B(new_n706), .C1(new_n728), .C2(new_n729), .ZN(G1328gat));
  AND2_X1   g529(.A1(new_n691), .A2(new_n694), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n203), .A3(new_n668), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT46), .Z(new_n733));
  NOR3_X1   g532(.A1(new_n724), .A2(new_n611), .A3(new_n726), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n203), .B2(new_n734), .ZN(G1329gat));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n210), .A3(new_n644), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(KEYINPUT47), .ZN(new_n737));
  AND4_X1   g536(.A1(new_n684), .A2(new_n721), .A3(new_n723), .A4(new_n725), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G43gat), .B1(new_n738), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n737), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n736), .B1(new_n738), .B2(new_n210), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n742), .A2(new_n745), .ZN(G1330gat));
  INV_X1    g545(.A(G50gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n747), .A3(new_n613), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n724), .A2(new_n656), .A3(new_n726), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n747), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT107), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT48), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  OAI221_X1 g552(.A(new_n748), .B1(new_n751), .B2(KEYINPUT48), .C1(new_n749), .C2(new_n747), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1331gat));
  NOR4_X1   g554(.A1(new_n692), .A2(new_n271), .A3(new_n303), .A4(new_n367), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n718), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n718), .A2(KEYINPUT108), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n603), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(new_n310), .ZN(G1332gat));
  INV_X1    g562(.A(KEYINPUT49), .ZN(new_n764));
  INV_X1    g563(.A(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n668), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT109), .Z(new_n767));
  OAI21_X1  g566(.A(KEYINPUT110), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n769));
  INV_X1    g568(.A(new_n767), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n759), .A2(new_n769), .A3(new_n760), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n764), .A2(new_n765), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1333gat));
  INV_X1    g573(.A(new_n684), .ZN(new_n775));
  OAI21_X1  g574(.A(G71gat), .B1(new_n761), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n644), .A2(new_n318), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n761), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n761), .A2(new_n656), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(new_n319), .ZN(G1335gat));
  NOR3_X1   g581(.A1(new_n342), .A2(new_n271), .A3(new_n367), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n721), .A2(new_n723), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784), .B2(new_n603), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n342), .A2(new_n271), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n718), .A2(new_n303), .A3(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n718), .A2(KEYINPUT51), .A3(new_n303), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n367), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n604), .A2(new_n281), .A3(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n785), .B1(new_n792), .B2(new_n794), .ZN(G1336gat));
  OAI21_X1  g594(.A(G92gat), .B1(new_n784), .B2(new_n611), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n791), .A2(new_n282), .A3(new_n668), .A4(new_n793), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT52), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n796), .A2(new_n797), .A3(new_n798), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1337gat));
  OAI21_X1  g602(.A(G99gat), .B1(new_n784), .B2(new_n775), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n680), .A2(G99gat), .A3(new_n367), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT112), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n792), .B2(new_n806), .ZN(G1338gat));
  NOR3_X1   g606(.A1(new_n656), .A2(G106gat), .A3(new_n367), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT53), .B1(new_n791), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n721), .A2(new_n613), .A3(new_n723), .A4(new_n783), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(G106gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n809), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n810), .A2(new_n812), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n791), .A2(new_n808), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n819), .B2(KEYINPUT53), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT114), .B(new_n821), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n815), .B1(new_n820), .B2(new_n822), .ZN(G1339gat));
  NOR2_X1   g622(.A1(new_n368), .A2(new_n271), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(new_n344), .C1(new_n355), .C2(new_n357), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n355), .A2(new_n357), .A3(new_n344), .ZN(new_n827));
  OAI211_X1 g626(.A(KEYINPUT54), .B(new_n358), .C1(new_n827), .C2(KEYINPUT116), .ZN(new_n828));
  INV_X1    g627(.A(new_n355), .ZN(new_n829));
  INV_X1    g628(.A(new_n357), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n345), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n364), .B(new_n826), .C1(new_n828), .C2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n301), .A3(new_n302), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n364), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(KEYINPUT117), .C1(new_n828), .C2(new_n833), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n366), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n831), .A2(new_n832), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT116), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n842), .A2(new_n843), .A3(KEYINPUT54), .A4(new_n358), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT117), .B1(new_n844), .B2(new_n839), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n257), .A2(new_n258), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n247), .B1(new_n246), .B2(new_n253), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n266), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n270), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT118), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(KEYINPUT118), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n838), .A2(new_n846), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n850), .A2(new_n367), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n269), .A2(new_n270), .B1(new_n834), .B2(new_n835), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n846), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n304), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n854), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n839), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n366), .A3(new_n840), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n271), .A2(new_n836), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n859), .B(new_n857), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n853), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n824), .B1(new_n867), .B2(new_n692), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n680), .A3(new_n613), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n603), .A2(new_n668), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n272), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n868), .A2(new_n603), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n713), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT120), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n873), .A2(KEYINPUT120), .A3(new_n713), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n611), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n272), .A2(G113gat), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT121), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n872), .B1(new_n879), .B2(new_n881), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n871), .A2(new_n883), .A3(new_n367), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n878), .A2(new_n611), .A3(new_n793), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n883), .ZN(G1341gat));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n692), .A2(G127gat), .ZN(new_n888));
  AOI211_X1 g687(.A(new_n668), .B(new_n888), .C1(new_n876), .C2(new_n877), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n869), .A2(new_n342), .A3(new_n870), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G127gat), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g692(.A(KEYINPUT122), .B(new_n891), .C1(new_n879), .C2(new_n888), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1342gat));
  INV_X1    g694(.A(G134gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n304), .A2(new_n668), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n878), .A2(new_n900), .A3(new_n896), .A4(new_n897), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n871), .B2(new_n304), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(G1343gat));
  NOR2_X1   g702(.A1(new_n868), .A2(new_n656), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n775), .A2(new_n870), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n856), .A2(new_n303), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n342), .B1(new_n908), .B2(new_n853), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n613), .B1(new_n909), .B2(new_n824), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(G141gat), .B1(new_n912), .B2(new_n272), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n684), .A2(new_n656), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n873), .A2(new_n611), .A3(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n378), .A3(new_n271), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1344gat));
  NOR3_X1   g719(.A1(new_n915), .A2(G148gat), .A3(new_n367), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT124), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT59), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT57), .B1(new_n868), .B2(new_n656), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n905), .B(new_n613), .C1(new_n909), .C2(new_n824), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR3_X1    g725(.A1(new_n926), .A2(new_n367), .A3(new_n907), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n923), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n367), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(KEYINPUT59), .A3(new_n380), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n922), .B1(new_n928), .B2(new_n930), .ZN(G1345gat));
  OAI21_X1  g730(.A(G155gat), .B1(new_n912), .B2(new_n692), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n335), .A3(new_n342), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n912), .B2(new_n304), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n873), .A2(new_n384), .A3(new_n897), .A4(new_n914), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n868), .A2(new_n604), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n713), .A2(new_n668), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n271), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n604), .A2(new_n611), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n869), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n944), .A2(new_n471), .A3(new_n272), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n942), .A2(new_n945), .ZN(G1348gat));
  NAND3_X1  g745(.A1(new_n941), .A2(new_n472), .A3(new_n793), .ZN(new_n947));
  OAI21_X1  g746(.A(G176gat), .B1(new_n944), .B2(new_n367), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(G1349gat));
  OAI21_X1  g748(.A(G183gat), .B1(new_n944), .B2(new_n692), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n342), .A2(new_n440), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n940), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n941), .A2(new_n441), .A3(new_n303), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n869), .A2(new_n303), .A3(new_n943), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(G190gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n955), .B2(G190gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(G1351gat));
  NOR3_X1   g758(.A1(new_n684), .A2(new_n611), .A3(new_n656), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n938), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n271), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n684), .A2(new_n604), .A3(new_n611), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n926), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n271), .A2(G197gat), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1352gat));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n793), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n968), .A2(G204gat), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n367), .A2(G204gat), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n961), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n973), .B1(new_n972), .B2(new_n970), .ZN(new_n974));
  AND4_X1   g773(.A1(new_n973), .A2(new_n961), .A3(new_n970), .A4(new_n971), .ZN(new_n975));
  OAI221_X1 g774(.A(new_n969), .B1(new_n970), .B2(new_n972), .C1(new_n974), .C2(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n498), .A3(new_n342), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n924), .A2(new_n342), .A3(new_n925), .A4(new_n963), .ZN(new_n978));
  OAI21_X1  g777(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n981));
  AND3_X1   g780(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n981), .B1(new_n978), .B2(new_n980), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n977), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(KEYINPUT127), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n986), .B(new_n977), .C1(new_n982), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n985), .A2(new_n987), .ZN(G1354gat));
  NAND3_X1  g787(.A1(new_n961), .A2(new_n499), .A3(new_n303), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n926), .A2(new_n304), .A3(new_n964), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n499), .ZN(G1355gat));
endmodule


