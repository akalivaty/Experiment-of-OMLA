

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XOR2_X1 U323 ( .A(G78GAT), .B(G204GAT), .Z(n291) );
  XNOR2_X1 U324 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n371) );
  XNOR2_X1 U325 ( .A(n372), .B(n371), .ZN(n373) );
  INV_X1 U326 ( .A(KEYINPUT31), .ZN(n352) );
  XNOR2_X1 U327 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U328 ( .A(n423), .B(n354), .ZN(n358) );
  XNOR2_X1 U329 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n378) );
  XNOR2_X1 U330 ( .A(n361), .B(n399), .ZN(n362) );
  XNOR2_X1 U331 ( .A(n379), .B(n378), .ZN(n524) );
  XNOR2_X1 U332 ( .A(n363), .B(n362), .ZN(n365) );
  OR2_X1 U333 ( .A1(n450), .A2(KEYINPUT124), .ZN(n451) );
  XOR2_X1 U334 ( .A(n555), .B(KEYINPUT28), .Z(n527) );
  XNOR2_X1 U335 ( .A(n453), .B(G218GAT), .ZN(n454) );
  XNOR2_X1 U336 ( .A(n455), .B(n454), .ZN(G1355GAT) );
  XOR2_X1 U337 ( .A(G43GAT), .B(G29GAT), .Z(n293) );
  XNOR2_X1 U338 ( .A(G50GAT), .B(KEYINPUT7), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U340 ( .A(n294), .B(KEYINPUT71), .Z(n296) );
  XNOR2_X1 U341 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n323) );
  XOR2_X1 U343 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n298) );
  XNOR2_X1 U344 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n323), .B(n299), .ZN(n310) );
  XNOR2_X1 U347 ( .A(G99GAT), .B(G85GAT), .ZN(n364) );
  XOR2_X1 U348 ( .A(KEYINPUT10), .B(G92GAT), .Z(n301) );
  XNOR2_X1 U349 ( .A(G134GAT), .B(G162GAT), .ZN(n300) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n364), .B(n302), .ZN(n304) );
  NAND2_X1 U352 ( .A1(G232GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U353 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U354 ( .A(n305), .B(KEYINPUT9), .Z(n308) );
  XNOR2_X1 U355 ( .A(G190GAT), .B(G218GAT), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n306), .B(KEYINPUT80), .ZN(n380) );
  XNOR2_X1 U357 ( .A(n380), .B(KEYINPUT65), .ZN(n307) );
  XNOR2_X1 U358 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U359 ( .A(n310), .B(n309), .Z(n571) );
  XNOR2_X1 U360 ( .A(KEYINPUT36), .B(KEYINPUT100), .ZN(n311) );
  XOR2_X1 U361 ( .A(n571), .B(n311), .Z(n484) );
  XOR2_X1 U362 ( .A(G169GAT), .B(G8GAT), .Z(n390) );
  XOR2_X1 U363 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n313) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(KEYINPUT66), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U366 ( .A(n390), .B(n314), .Z(n316) );
  NAND2_X1 U367 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n327) );
  XOR2_X1 U369 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n318) );
  XNOR2_X1 U370 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n320) );
  XNOR2_X1 U372 ( .A(G113GAT), .B(G141GAT), .ZN(n319) );
  XNOR2_X1 U373 ( .A(n319), .B(G1GAT), .ZN(n407) );
  XOR2_X1 U374 ( .A(n320), .B(n407), .Z(n325) );
  XOR2_X1 U375 ( .A(KEYINPUT72), .B(KEYINPUT73), .Z(n322) );
  XNOR2_X1 U376 ( .A(G15GAT), .B(G22GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n337) );
  XNOR2_X1 U378 ( .A(n323), .B(n337), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n543) );
  XOR2_X1 U381 ( .A(n543), .B(KEYINPUT74), .Z(n562) );
  XOR2_X1 U382 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n350) );
  XOR2_X1 U383 ( .A(G64GAT), .B(G57GAT), .Z(n329) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(G78GAT), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U386 ( .A(KEYINPUT83), .B(KEYINPUT81), .Z(n331) );
  XNOR2_X1 U387 ( .A(G1GAT), .B(KEYINPUT82), .ZN(n330) );
  XNOR2_X1 U388 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U389 ( .A(n333), .B(n332), .Z(n339) );
  XOR2_X1 U390 ( .A(G211GAT), .B(G155GAT), .Z(n335) );
  XNOR2_X1 U391 ( .A(G127GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n348) );
  XOR2_X1 U395 ( .A(KEYINPUT85), .B(KEYINPUT12), .Z(n341) );
  XNOR2_X1 U396 ( .A(KEYINPUT84), .B(KEYINPUT14), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n346) );
  XNOR2_X1 U398 ( .A(G71GAT), .B(KEYINPUT75), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n342), .B(KEYINPUT13), .ZN(n360) );
  XOR2_X1 U400 ( .A(n360), .B(KEYINPUT15), .Z(n344) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U403 ( .A(n346), .B(n345), .Z(n347) );
  XOR2_X1 U404 ( .A(n348), .B(n347), .Z(n551) );
  INV_X1 U405 ( .A(n551), .ZN(n587) );
  NAND2_X1 U406 ( .A1(n484), .A2(n587), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n366) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n291), .B(n351), .ZN(n423) );
  NAND2_X1 U410 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XOR2_X1 U411 ( .A(KEYINPUT32), .B(KEYINPUT77), .Z(n356) );
  XNOR2_X1 U412 ( .A(G148GAT), .B(KEYINPUT33), .ZN(n355) );
  XOR2_X1 U413 ( .A(n356), .B(n355), .Z(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n363) );
  XNOR2_X1 U415 ( .A(G176GAT), .B(G92GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n359), .B(G64GAT), .ZN(n381) );
  XNOR2_X1 U417 ( .A(n360), .B(n381), .ZN(n361) );
  XOR2_X1 U418 ( .A(G120GAT), .B(G57GAT), .Z(n399) );
  XOR2_X1 U419 ( .A(n365), .B(n364), .Z(n369) );
  INV_X1 U420 ( .A(n369), .ZN(n456) );
  NAND2_X1 U421 ( .A1(n366), .A2(n456), .ZN(n367) );
  NOR2_X1 U422 ( .A1(n562), .A2(n367), .ZN(n368) );
  XOR2_X1 U423 ( .A(KEYINPUT113), .B(n368), .Z(n377) );
  INV_X1 U424 ( .A(n571), .ZN(n535) );
  INV_X1 U425 ( .A(KEYINPUT41), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n499) );
  INV_X1 U427 ( .A(n543), .ZN(n582) );
  NAND2_X1 U428 ( .A1(n499), .A2(n582), .ZN(n372) );
  NAND2_X1 U429 ( .A1(n373), .A2(n551), .ZN(n374) );
  NOR2_X1 U430 ( .A1(n535), .A2(n374), .ZN(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT47), .B(n375), .Z(n376) );
  NOR2_X1 U432 ( .A1(n377), .A2(n376), .ZN(n379) );
  XOR2_X1 U433 ( .A(n381), .B(n380), .Z(n386) );
  XOR2_X1 U434 ( .A(G183GAT), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U435 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n433) );
  XNOR2_X1 U437 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n384), .B(G211GAT), .ZN(n419) );
  XNOR2_X1 U439 ( .A(n433), .B(n419), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n386), .B(n385), .ZN(n394) );
  XOR2_X1 U441 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n388) );
  XNOR2_X1 U442 ( .A(G36GAT), .B(G204GAT), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U444 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U445 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U447 ( .A(n394), .B(n393), .Z(n516) );
  NOR2_X1 U448 ( .A1(n524), .A2(n516), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n395), .B(KEYINPUT54), .ZN(n559) );
  XOR2_X1 U450 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n397) );
  XNOR2_X1 U451 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U453 ( .A(n398), .B(G85GAT), .Z(n401) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n411) );
  XOR2_X1 U456 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n403) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U459 ( .A(n404), .B(KEYINPUT4), .Z(n409) );
  XOR2_X1 U460 ( .A(G127GAT), .B(KEYINPUT86), .Z(n406) );
  XNOR2_X1 U461 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n444) );
  XNOR2_X1 U463 ( .A(n407), .B(n444), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT3), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U467 ( .A(G155GAT), .B(G148GAT), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(KEYINPUT2), .B(n414), .ZN(n428) );
  INV_X1 U470 ( .A(n428), .ZN(n415) );
  XOR2_X1 U471 ( .A(n416), .B(n415), .Z(n469) );
  XNOR2_X1 U472 ( .A(KEYINPUT93), .B(n469), .ZN(n557) );
  NAND2_X1 U473 ( .A1(n559), .A2(n557), .ZN(n449) );
  XOR2_X1 U474 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n448) );
  XOR2_X1 U475 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n422) );
  XOR2_X1 U476 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n418) );
  XNOR2_X1 U477 ( .A(G22GAT), .B(G141GAT), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U481 ( .A(G218GAT), .B(n423), .Z(n425) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U484 ( .A(n427), .B(n426), .Z(n430) );
  XOR2_X1 U485 ( .A(G50GAT), .B(n428), .Z(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n555) );
  XOR2_X1 U487 ( .A(G99GAT), .B(G43GAT), .Z(n432) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U490 ( .A(n434), .B(n433), .Z(n442) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n436) );
  XNOR2_X1 U492 ( .A(G190GAT), .B(KEYINPUT88), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U494 ( .A(G120GAT), .B(G176GAT), .Z(n438) );
  XNOR2_X1 U495 ( .A(G169GAT), .B(G15GAT), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U499 ( .A(n443), .B(G71GAT), .Z(n446) );
  XNOR2_X1 U500 ( .A(G113GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n572) );
  NAND2_X1 U502 ( .A1(n555), .A2(n572), .ZN(n447) );
  XOR2_X1 U503 ( .A(n448), .B(n447), .Z(n541) );
  INV_X1 U504 ( .A(n541), .ZN(n465) );
  NOR2_X1 U505 ( .A1(n449), .A2(n465), .ZN(n450) );
  NAND2_X1 U506 ( .A1(n450), .A2(KEYINPUT124), .ZN(n452) );
  NAND2_X1 U507 ( .A1(n452), .A2(n451), .ZN(n581) );
  NAND2_X1 U508 ( .A1(n484), .A2(n581), .ZN(n455) );
  XOR2_X1 U509 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n453) );
  NAND2_X1 U510 ( .A1(n562), .A2(n456), .ZN(n487) );
  NOR2_X1 U511 ( .A1(n535), .A2(n551), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n457), .B(KEYINPUT16), .ZN(n473) );
  INV_X1 U513 ( .A(n527), .ZN(n459) );
  XNOR2_X1 U514 ( .A(n516), .B(KEYINPUT27), .ZN(n464) );
  NOR2_X1 U515 ( .A1(n557), .A2(n464), .ZN(n525) );
  NAND2_X1 U516 ( .A1(n572), .A2(n525), .ZN(n458) );
  NOR2_X1 U517 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT96), .ZN(n471) );
  NOR2_X1 U519 ( .A1(n572), .A2(n516), .ZN(n461) );
  NOR2_X1 U520 ( .A1(n555), .A2(n461), .ZN(n462) );
  XOR2_X1 U521 ( .A(n462), .B(KEYINPUT98), .Z(n463) );
  XNOR2_X1 U522 ( .A(KEYINPUT25), .B(n463), .ZN(n467) );
  NOR2_X1 U523 ( .A1(n465), .A2(n464), .ZN(n466) );
  NOR2_X1 U524 ( .A1(n467), .A2(n466), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n482) );
  INV_X1 U527 ( .A(n482), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n500) );
  OR2_X1 U529 ( .A1(n487), .A2(n500), .ZN(n480) );
  NOR2_X1 U530 ( .A1(n557), .A2(n480), .ZN(n474) );
  XOR2_X1 U531 ( .A(n474), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NOR2_X1 U533 ( .A1(n516), .A2(n480), .ZN(n476) );
  XOR2_X1 U534 ( .A(G8GAT), .B(n476), .Z(G1325GAT) );
  NOR2_X1 U535 ( .A1(n572), .A2(n480), .ZN(n478) );
  XNOR2_X1 U536 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U538 ( .A(G15GAT), .B(n479), .Z(G1326GAT) );
  NOR2_X1 U539 ( .A1(n527), .A2(n480), .ZN(n481) );
  XOR2_X1 U540 ( .A(G22GAT), .B(n481), .Z(G1327GAT) );
  XNOR2_X1 U541 ( .A(KEYINPUT37), .B(KEYINPUT101), .ZN(n486) );
  NOR2_X1 U542 ( .A1(n482), .A2(n587), .ZN(n483) );
  NAND2_X1 U543 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n512) );
  NOR2_X1 U545 ( .A1(n512), .A2(n487), .ZN(n489) );
  XNOR2_X1 U546 ( .A(KEYINPUT103), .B(KEYINPUT38), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT102), .B(n490), .ZN(n496) );
  NOR2_X1 U549 ( .A1(n557), .A2(n496), .ZN(n492) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n516), .A2(n496), .ZN(n493) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n493), .Z(G1329GAT) );
  NOR2_X1 U554 ( .A1(n572), .A2(n496), .ZN(n494) );
  XOR2_X1 U555 ( .A(KEYINPUT40), .B(n494), .Z(n495) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U557 ( .A1(n527), .A2(n496), .ZN(n497) );
  XOR2_X1 U558 ( .A(G50GAT), .B(n497), .Z(n498) );
  XNOR2_X1 U559 ( .A(KEYINPUT104), .B(n498), .ZN(G1331GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n543), .ZN(n513) );
  NOR2_X1 U561 ( .A1(n513), .A2(n500), .ZN(n501) );
  XNOR2_X1 U562 ( .A(KEYINPUT105), .B(n501), .ZN(n507) );
  NOR2_X1 U563 ( .A1(n557), .A2(n507), .ZN(n502) );
  XOR2_X1 U564 ( .A(G57GAT), .B(n502), .Z(n503) );
  XNOR2_X1 U565 ( .A(KEYINPUT42), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n516), .A2(n507), .ZN(n504) );
  XOR2_X1 U567 ( .A(G64GAT), .B(n504), .Z(G1333GAT) );
  NOR2_X1 U568 ( .A1(n572), .A2(n507), .ZN(n505) );
  XOR2_X1 U569 ( .A(KEYINPUT106), .B(n505), .Z(n506) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  NOR2_X1 U571 ( .A1(n507), .A2(n527), .ZN(n511) );
  XOR2_X1 U572 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n509) );
  XNOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT107), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NOR2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(KEYINPUT109), .ZN(n521) );
  NOR2_X1 U578 ( .A1(n557), .A2(n521), .ZN(n515) );
  XOR2_X1 U579 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  NOR2_X1 U580 ( .A1(n516), .A2(n521), .ZN(n517) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n572), .A2(n521), .ZN(n518) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT110), .B(KEYINPUT44), .Z(n520) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(n523) );
  NOR2_X1 U587 ( .A1(n527), .A2(n521), .ZN(n522) );
  XOR2_X1 U588 ( .A(n523), .B(n522), .Z(G1339GAT) );
  INV_X1 U589 ( .A(n525), .ZN(n526) );
  NOR2_X1 U590 ( .A1(n524), .A2(n526), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n527), .A2(n542), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n572), .A2(n528), .ZN(n536) );
  NAND2_X1 U593 ( .A1(n536), .A2(n562), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U596 ( .A1(n536), .A2(n499), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n533) );
  NAND2_X1 U599 ( .A1(n536), .A2(n587), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n538) );
  NAND2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n540) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT117), .Z(n539) );
  XNOR2_X1 U606 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n543), .A2(n553), .ZN(n544) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  INV_X1 U610 ( .A(n499), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n545), .A2(n553), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U615 ( .A(KEYINPUT53), .B(n548), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U617 ( .A1(n551), .A2(n553), .ZN(n552) );
  XOR2_X1 U618 ( .A(G155GAT), .B(n552), .Z(G1346GAT) );
  NOR2_X1 U619 ( .A1(n571), .A2(n553), .ZN(n554) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  INV_X1 U621 ( .A(n555), .ZN(n556) );
  AND2_X1 U622 ( .A1(n557), .A2(n556), .ZN(n558) );
  AND2_X1 U623 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U624 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n560) );
  XNOR2_X1 U625 ( .A(n561), .B(n560), .ZN(n574) );
  NOR2_X1 U626 ( .A1(n574), .A2(n572), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n569), .A2(n562), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n565) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(n566), .Z(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n499), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n587), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n576) );
  OR2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  OR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(n577), .ZN(G1351GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT126), .Z(n579) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(n580), .Z(n584) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  NAND2_X1 U649 ( .A1(n369), .A2(n581), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n581), .A2(n587), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
endmodule

