

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n709), .A2(n594), .ZN(n620) );
  NOR2_X4 U554 ( .A1(G651), .A2(n538), .ZN(n782) );
  XNOR2_X2 U555 ( .A(n520), .B(n519), .ZN(n889) );
  NOR2_X1 U556 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U557 ( .A1(n634), .A2(n633), .ZN(n635) );
  INV_X1 U558 ( .A(KEYINPUT17), .ZN(n519) );
  XOR2_X1 U559 ( .A(n608), .B(KEYINPUT28), .Z(n518) );
  XNOR2_X1 U560 ( .A(KEYINPUT101), .B(KEYINPUT29), .ZN(n647) );
  XNOR2_X1 U561 ( .A(n648), .B(n647), .ZN(n651) );
  NOR2_X1 U562 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U563 ( .A1(G2084), .A2(n657), .ZN(n596) );
  NOR2_X1 U564 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U565 ( .A1(n719), .A2(n679), .ZN(n681) );
  NOR2_X1 U566 ( .A1(n676), .A2(n675), .ZN(n719) );
  NOR2_X1 U567 ( .A1(n685), .A2(n684), .ZN(n715) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n709) );
  XNOR2_X1 U569 ( .A(n637), .B(KEYINPUT15), .ZN(n927) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n528), .Z(n783) );
  NAND2_X1 U571 ( .A1(n751), .A2(n750), .ZN(n752) );
  AND2_X1 U572 ( .A1(n889), .A2(G138), .ZN(n527) );
  NOR2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  INV_X1 U574 ( .A(G2104), .ZN(n521) );
  NOR2_X1 U575 ( .A1(G2105), .A2(n521), .ZN(n586) );
  BUF_X1 U576 ( .A(n586), .Z(n887) );
  NAND2_X1 U577 ( .A1(G102), .A2(n887), .ZN(n525) );
  AND2_X1 U578 ( .A1(G2105), .A2(G2104), .ZN(n883) );
  NAND2_X1 U579 ( .A1(G114), .A2(n883), .ZN(n523) );
  AND2_X1 U580 ( .A1(n521), .A2(G2105), .ZN(n881) );
  NAND2_X1 U581 ( .A1(G126), .A2(n881), .ZN(n522) );
  AND2_X1 U582 ( .A1(n523), .A2(n522), .ZN(n524) );
  NAND2_X1 U583 ( .A1(n525), .A2(n524), .ZN(n526) );
  NOR2_X1 U584 ( .A1(n527), .A2(n526), .ZN(G164) );
  INV_X1 U585 ( .A(G651), .ZN(n537) );
  NOR2_X1 U586 ( .A1(G543), .A2(n537), .ZN(n528) );
  XOR2_X1 U587 ( .A(G543), .B(KEYINPUT0), .Z(n538) );
  NAND2_X1 U588 ( .A1(G49), .A2(n782), .ZN(n530) );
  NAND2_X1 U589 ( .A1(G74), .A2(G651), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n783), .A2(n531), .ZN(n532) );
  XOR2_X1 U592 ( .A(KEYINPUT81), .B(n532), .Z(n534) );
  NAND2_X1 U593 ( .A1(n538), .A2(G87), .ZN(n533) );
  NAND2_X1 U594 ( .A1(n534), .A2(n533), .ZN(G288) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n535) );
  XNOR2_X1 U596 ( .A(n535), .B(KEYINPUT64), .ZN(n788) );
  NAND2_X1 U597 ( .A1(G89), .A2(n788), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n536), .B(KEYINPUT4), .ZN(n540) );
  NOR2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n787) );
  NAND2_X1 U600 ( .A1(G76), .A2(n787), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U602 ( .A(n541), .B(KEYINPUT5), .ZN(n547) );
  NAND2_X1 U603 ( .A1(n783), .A2(G63), .ZN(n542) );
  XNOR2_X1 U604 ( .A(n542), .B(KEYINPUT74), .ZN(n544) );
  NAND2_X1 U605 ( .A1(G51), .A2(n782), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U609 ( .A(n548), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U610 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U611 ( .A1(G52), .A2(n782), .ZN(n550) );
  NAND2_X1 U612 ( .A1(G64), .A2(n783), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G77), .A2(n787), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G90), .A2(n788), .ZN(n551) );
  NAND2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U617 ( .A(KEYINPUT67), .B(n553), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT9), .B(n554), .ZN(n555) );
  NOR2_X1 U619 ( .A1(n556), .A2(n555), .ZN(G171) );
  NAND2_X1 U620 ( .A1(G78), .A2(n787), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n557), .B(KEYINPUT68), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n782), .A2(G53), .ZN(n559) );
  NAND2_X1 U623 ( .A1(G91), .A2(n788), .ZN(n558) );
  NAND2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G65), .A2(n783), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT69), .B(n560), .ZN(n561) );
  NOR2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(G299) );
  NAND2_X1 U629 ( .A1(n782), .A2(G50), .ZN(n566) );
  NAND2_X1 U630 ( .A1(G88), .A2(n788), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G75), .A2(n787), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT82), .B(n567), .Z(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n783), .A2(G62), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(G303) );
  NAND2_X1 U637 ( .A1(n782), .A2(G48), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G86), .A2(n788), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U640 ( .A1(n787), .A2(G73), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n574), .Z(n575) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n783), .A2(G61), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G72), .A2(n787), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G85), .A2(n788), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G47), .A2(n782), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G60), .A2(n783), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U652 ( .A(KEYINPUT66), .B(n585), .Z(G290) );
  INV_X1 U653 ( .A(G303), .ZN(G166) );
  NAND2_X1 U654 ( .A1(G101), .A2(n586), .ZN(n587) );
  XNOR2_X1 U655 ( .A(n587), .B(KEYINPUT65), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT23), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G137), .A2(n889), .ZN(n589) );
  AND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n754) );
  NAND2_X1 U659 ( .A1(G113), .A2(n883), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G125), .A2(n881), .ZN(n591) );
  AND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n753) );
  AND2_X1 U662 ( .A1(G40), .A2(n753), .ZN(n593) );
  NAND2_X1 U663 ( .A1(n754), .A2(n593), .ZN(n708) );
  INV_X1 U664 ( .A(n708), .ZN(n594) );
  INV_X1 U665 ( .A(n620), .ZN(n657) );
  NAND2_X1 U666 ( .A1(G8), .A2(n657), .ZN(n724) );
  NOR2_X1 U667 ( .A1(G1976), .A2(G288), .ZN(n678) );
  NAND2_X1 U668 ( .A1(n678), .A2(KEYINPUT33), .ZN(n595) );
  NOR2_X1 U669 ( .A1(n724), .A2(n595), .ZN(n685) );
  XOR2_X1 U670 ( .A(KEYINPUT106), .B(KEYINPUT32), .Z(n666) );
  NOR2_X1 U671 ( .A1(G1966), .A2(n724), .ZN(n671) );
  XNOR2_X1 U672 ( .A(KEYINPUT97), .B(n596), .ZN(n667) );
  NAND2_X1 U673 ( .A1(G8), .A2(n667), .ZN(n597) );
  NOR2_X1 U674 ( .A1(n671), .A2(n597), .ZN(n598) );
  XOR2_X1 U675 ( .A(KEYINPUT30), .B(n598), .Z(n599) );
  NOR2_X1 U676 ( .A1(G168), .A2(n599), .ZN(n603) );
  XNOR2_X1 U677 ( .A(G2078), .B(KEYINPUT25), .ZN(n999) );
  NOR2_X1 U678 ( .A1(n657), .A2(n999), .ZN(n601) );
  XOR2_X1 U679 ( .A(KEYINPUT98), .B(G1961), .Z(n976) );
  NOR2_X1 U680 ( .A1(n620), .A2(n976), .ZN(n600) );
  NOR2_X1 U681 ( .A1(n601), .A2(n600), .ZN(n649) );
  NOR2_X1 U682 ( .A1(G171), .A2(n649), .ZN(n602) );
  XNOR2_X1 U683 ( .A(KEYINPUT31), .B(n604), .ZN(n655) );
  INV_X1 U684 ( .A(KEYINPUT102), .ZN(n653) );
  NAND2_X1 U685 ( .A1(n620), .A2(G2072), .ZN(n605) );
  XNOR2_X1 U686 ( .A(n605), .B(KEYINPUT27), .ZN(n607) );
  INV_X1 U687 ( .A(G1956), .ZN(n980) );
  NOR2_X1 U688 ( .A1(n980), .A2(n620), .ZN(n606) );
  NOR2_X1 U689 ( .A1(n607), .A2(n606), .ZN(n643) );
  INV_X1 U690 ( .A(G299), .ZN(n799) );
  NOR2_X1 U691 ( .A1(n643), .A2(n799), .ZN(n608) );
  NAND2_X1 U692 ( .A1(G56), .A2(n783), .ZN(n609) );
  XOR2_X1 U693 ( .A(KEYINPUT14), .B(n609), .Z(n615) );
  NAND2_X1 U694 ( .A1(G81), .A2(n788), .ZN(n610) );
  XNOR2_X1 U695 ( .A(n610), .B(KEYINPUT12), .ZN(n612) );
  NAND2_X1 U696 ( .A1(G68), .A2(n787), .ZN(n611) );
  NAND2_X1 U697 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U698 ( .A(KEYINPUT13), .B(n613), .Z(n614) );
  NOR2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U700 ( .A1(n782), .A2(G43), .ZN(n616) );
  NAND2_X1 U701 ( .A1(n617), .A2(n616), .ZN(n920) );
  INV_X1 U702 ( .A(G1341), .ZN(n981) );
  NOR2_X1 U703 ( .A1(n620), .A2(n981), .ZN(n622) );
  AND2_X1 U704 ( .A1(n622), .A2(KEYINPUT26), .ZN(n618) );
  NOR2_X1 U705 ( .A1(KEYINPUT100), .A2(n618), .ZN(n619) );
  NOR2_X1 U706 ( .A1(n920), .A2(n619), .ZN(n627) );
  XOR2_X1 U707 ( .A(G1996), .B(KEYINPUT99), .Z(n1007) );
  NAND2_X1 U708 ( .A1(n620), .A2(n1007), .ZN(n621) );
  XNOR2_X1 U709 ( .A(n621), .B(KEYINPUT26), .ZN(n624) );
  INV_X1 U710 ( .A(n622), .ZN(n623) );
  NAND2_X1 U711 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U712 ( .A1(KEYINPUT100), .A2(n625), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n639) );
  AND2_X1 U714 ( .A1(n657), .A2(G1348), .ZN(n629) );
  INV_X1 U715 ( .A(G2067), .ZN(n1001) );
  NOR2_X1 U716 ( .A1(n657), .A2(n1001), .ZN(n628) );
  NOR2_X1 U717 ( .A1(n629), .A2(n628), .ZN(n640) );
  NAND2_X1 U718 ( .A1(G66), .A2(n783), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G79), .A2(n787), .ZN(n631) );
  NAND2_X1 U720 ( .A1(G92), .A2(n788), .ZN(n630) );
  NAND2_X1 U721 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U722 ( .A1(G54), .A2(n782), .ZN(n632) );
  XNOR2_X1 U723 ( .A(KEYINPUT73), .B(n632), .ZN(n633) );
  NAND2_X1 U724 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U725 ( .A1(n640), .A2(n927), .ZN(n638) );
  NAND2_X1 U726 ( .A1(n639), .A2(n638), .ZN(n642) );
  OR2_X1 U727 ( .A1(n640), .A2(n927), .ZN(n641) );
  NAND2_X1 U728 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n799), .A2(n643), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n518), .A2(n646), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G171), .A2(n649), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n656), .B(KEYINPUT103), .ZN(n669) );
  NAND2_X1 U736 ( .A1(G286), .A2(n669), .ZN(n663) );
  NOR2_X1 U737 ( .A1(G1971), .A2(n724), .ZN(n659) );
  NOR2_X1 U738 ( .A1(G2090), .A2(n657), .ZN(n658) );
  NOR2_X1 U739 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U740 ( .A(KEYINPUT105), .B(n660), .Z(n661) );
  NAND2_X1 U741 ( .A1(n661), .A2(G303), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(G8), .A2(n664), .ZN(n665) );
  XNOR2_X1 U744 ( .A(n666), .B(n665), .ZN(n676) );
  INV_X1 U745 ( .A(G8), .ZN(n668) );
  NOR2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n674) );
  INV_X1 U747 ( .A(n669), .ZN(n670) );
  XOR2_X1 U748 ( .A(KEYINPUT104), .B(n672), .Z(n673) );
  NOR2_X1 U749 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U750 ( .A1(G1971), .A2(G303), .ZN(n677) );
  NOR2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n931) );
  INV_X1 U752 ( .A(n931), .ZN(n679) );
  NAND2_X1 U753 ( .A1(G288), .A2(G1976), .ZN(n680) );
  XOR2_X1 U754 ( .A(KEYINPUT107), .B(n680), .Z(n922) );
  NAND2_X1 U755 ( .A1(n681), .A2(n922), .ZN(n682) );
  NOR2_X1 U756 ( .A1(n724), .A2(n682), .ZN(n683) );
  NOR2_X1 U757 ( .A1(KEYINPUT33), .A2(n683), .ZN(n684) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n934) );
  NAND2_X1 U759 ( .A1(G141), .A2(n889), .ZN(n687) );
  NAND2_X1 U760 ( .A1(G129), .A2(n881), .ZN(n686) );
  NAND2_X1 U761 ( .A1(n687), .A2(n686), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n887), .A2(G105), .ZN(n688) );
  XOR2_X1 U763 ( .A(KEYINPUT38), .B(n688), .Z(n689) );
  NOR2_X1 U764 ( .A1(n690), .A2(n689), .ZN(n692) );
  NAND2_X1 U765 ( .A1(n883), .A2(G117), .ZN(n691) );
  NAND2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n897) );
  NOR2_X1 U767 ( .A1(G1996), .A2(n897), .ZN(n950) );
  NAND2_X1 U768 ( .A1(n897), .A2(G1996), .ZN(n703) );
  NAND2_X1 U769 ( .A1(G131), .A2(n889), .ZN(n694) );
  NAND2_X1 U770 ( .A1(G95), .A2(n887), .ZN(n693) );
  NAND2_X1 U771 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U772 ( .A(n695), .B(KEYINPUT95), .ZN(n700) );
  NAND2_X1 U773 ( .A1(G107), .A2(n883), .ZN(n697) );
  NAND2_X1 U774 ( .A1(G119), .A2(n881), .ZN(n696) );
  NAND2_X1 U775 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U776 ( .A(KEYINPUT94), .B(n698), .Z(n699) );
  NAND2_X1 U777 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U778 ( .A(n701), .B(KEYINPUT96), .ZN(n904) );
  NAND2_X1 U779 ( .A1(n904), .A2(G1991), .ZN(n702) );
  NAND2_X1 U780 ( .A1(n703), .A2(n702), .ZN(n963) );
  NOR2_X1 U781 ( .A1(G1986), .A2(G290), .ZN(n704) );
  NOR2_X1 U782 ( .A1(G1991), .A2(n904), .ZN(n943) );
  NOR2_X1 U783 ( .A1(n704), .A2(n943), .ZN(n705) );
  NOR2_X1 U784 ( .A1(n963), .A2(n705), .ZN(n706) );
  NOR2_X1 U785 ( .A1(n950), .A2(n706), .ZN(n707) );
  XNOR2_X1 U786 ( .A(KEYINPUT39), .B(n707), .ZN(n710) );
  NOR2_X1 U787 ( .A1(n709), .A2(n708), .ZN(n749) );
  AND2_X1 U788 ( .A1(n710), .A2(n749), .ZN(n726) );
  INV_X1 U789 ( .A(n963), .ZN(n711) );
  XOR2_X1 U790 ( .A(G1986), .B(G290), .Z(n930) );
  NAND2_X1 U791 ( .A1(n711), .A2(n930), .ZN(n712) );
  NAND2_X1 U792 ( .A1(n712), .A2(n749), .ZN(n713) );
  OR2_X1 U793 ( .A1(n726), .A2(n713), .ZN(n716) );
  AND2_X1 U794 ( .A1(n934), .A2(n716), .ZN(n714) );
  NAND2_X1 U795 ( .A1(n715), .A2(n714), .ZN(n732) );
  INV_X1 U796 ( .A(n716), .ZN(n730) );
  NAND2_X1 U797 ( .A1(G166), .A2(G8), .ZN(n717) );
  NOR2_X1 U798 ( .A1(G2090), .A2(n717), .ZN(n718) );
  NOR2_X1 U799 ( .A1(n719), .A2(n718), .ZN(n721) );
  INV_X1 U800 ( .A(n724), .ZN(n720) );
  NOR2_X1 U801 ( .A1(n721), .A2(n720), .ZN(n728) );
  NOR2_X1 U802 ( .A1(G1981), .A2(G305), .ZN(n722) );
  XOR2_X1 U803 ( .A(n722), .B(KEYINPUT24), .Z(n723) );
  NOR2_X1 U804 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U805 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U806 ( .A1(n728), .A2(n727), .ZN(n729) );
  OR2_X1 U807 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U808 ( .A1(n732), .A2(n731), .ZN(n747) );
  XOR2_X1 U809 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n745) );
  NAND2_X1 U810 ( .A1(G140), .A2(n889), .ZN(n734) );
  NAND2_X1 U811 ( .A1(G104), .A2(n887), .ZN(n733) );
  NAND2_X1 U812 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U813 ( .A(KEYINPUT34), .B(n735), .ZN(n742) );
  NAND2_X1 U814 ( .A1(n883), .A2(G116), .ZN(n736) );
  XNOR2_X1 U815 ( .A(n736), .B(KEYINPUT90), .ZN(n738) );
  NAND2_X1 U816 ( .A1(G128), .A2(n881), .ZN(n737) );
  NAND2_X1 U817 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U818 ( .A(KEYINPUT91), .B(n739), .ZN(n740) );
  XNOR2_X1 U819 ( .A(KEYINPUT35), .B(n740), .ZN(n741) );
  NOR2_X1 U820 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U821 ( .A(n743), .B(KEYINPUT36), .ZN(n744) );
  XNOR2_X1 U822 ( .A(n745), .B(n744), .ZN(n903) );
  XNOR2_X1 U823 ( .A(KEYINPUT37), .B(G2067), .ZN(n748) );
  NOR2_X1 U824 ( .A1(n903), .A2(n748), .ZN(n944) );
  NAND2_X1 U825 ( .A1(n944), .A2(n749), .ZN(n746) );
  NAND2_X1 U826 ( .A1(n747), .A2(n746), .ZN(n751) );
  AND2_X1 U827 ( .A1(n748), .A2(n903), .ZN(n955) );
  NAND2_X1 U828 ( .A1(n955), .A2(n749), .ZN(n750) );
  XNOR2_X1 U829 ( .A(n752), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U830 ( .A1(n754), .A2(n753), .ZN(G160) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  XOR2_X1 U832 ( .A(KEYINPUT78), .B(KEYINPUT18), .Z(n756) );
  NAND2_X1 U833 ( .A1(G123), .A2(n881), .ZN(n755) );
  XNOR2_X1 U834 ( .A(n756), .B(n755), .ZN(n760) );
  NAND2_X1 U835 ( .A1(G99), .A2(n887), .ZN(n758) );
  NAND2_X1 U836 ( .A1(G111), .A2(n883), .ZN(n757) );
  NAND2_X1 U837 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U838 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U839 ( .A1(n889), .A2(G135), .ZN(n761) );
  NAND2_X1 U840 ( .A1(n762), .A2(n761), .ZN(n956) );
  XNOR2_X1 U841 ( .A(G2096), .B(n956), .ZN(n763) );
  OR2_X1 U842 ( .A1(G2100), .A2(n763), .ZN(G156) );
  INV_X1 U843 ( .A(G57), .ZN(G237) );
  INV_X1 U844 ( .A(G132), .ZN(G219) );
  INV_X1 U845 ( .A(G82), .ZN(G220) );
  NAND2_X1 U846 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U847 ( .A(n764), .B(KEYINPUT10), .ZN(n765) );
  XNOR2_X1 U848 ( .A(KEYINPUT70), .B(n765), .ZN(G223) );
  INV_X1 U849 ( .A(G223), .ZN(n825) );
  NAND2_X1 U850 ( .A1(n825), .A2(G567), .ZN(n766) );
  XOR2_X1 U851 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U852 ( .A(G860), .ZN(n774) );
  OR2_X1 U853 ( .A1(n920), .A2(n774), .ZN(n767) );
  XOR2_X1 U854 ( .A(KEYINPUT71), .B(n767), .Z(G153) );
  XOR2_X1 U855 ( .A(G171), .B(KEYINPUT72), .Z(G301) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n769) );
  OR2_X1 U857 ( .A1(n927), .A2(G868), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(G284) );
  NOR2_X1 U859 ( .A1(G868), .A2(G299), .ZN(n770) );
  XOR2_X1 U860 ( .A(KEYINPUT75), .B(n770), .Z(n773) );
  INV_X1 U861 ( .A(G868), .ZN(n771) );
  NOR2_X1 U862 ( .A1(G286), .A2(n771), .ZN(n772) );
  NOR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U864 ( .A1(n774), .A2(G559), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n775), .A2(n927), .ZN(n776) );
  XNOR2_X1 U866 ( .A(n776), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U867 ( .A1(n927), .A2(G868), .ZN(n777) );
  NOR2_X1 U868 ( .A1(G559), .A2(n777), .ZN(n778) );
  XOR2_X1 U869 ( .A(KEYINPUT77), .B(n778), .Z(n781) );
  NOR2_X1 U870 ( .A1(G868), .A2(n920), .ZN(n779) );
  XNOR2_X1 U871 ( .A(KEYINPUT76), .B(n779), .ZN(n780) );
  NOR2_X1 U872 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U873 ( .A1(G55), .A2(n782), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G67), .A2(n783), .ZN(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U876 ( .A(KEYINPUT80), .B(n786), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G80), .A2(n787), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G93), .A2(n788), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n909) );
  NAND2_X1 U881 ( .A1(G559), .A2(n927), .ZN(n793) );
  XOR2_X1 U882 ( .A(n920), .B(n793), .Z(n804) );
  XNOR2_X1 U883 ( .A(KEYINPUT79), .B(n804), .ZN(n794) );
  NOR2_X1 U884 ( .A1(G860), .A2(n794), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n909), .B(n795), .ZN(G145) );
  XOR2_X1 U886 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n797) );
  XNOR2_X1 U887 ( .A(KEYINPUT85), .B(KEYINPUT83), .ZN(n796) );
  XNOR2_X1 U888 ( .A(n797), .B(n796), .ZN(n798) );
  XNOR2_X1 U889 ( .A(G288), .B(n798), .ZN(n801) );
  XNOR2_X1 U890 ( .A(G166), .B(n799), .ZN(n800) );
  XNOR2_X1 U891 ( .A(n801), .B(n800), .ZN(n802) );
  XNOR2_X1 U892 ( .A(G290), .B(n802), .ZN(n803) );
  XNOR2_X1 U893 ( .A(n803), .B(G305), .ZN(n908) );
  XNOR2_X1 U894 ( .A(n908), .B(n804), .ZN(n805) );
  NAND2_X1 U895 ( .A1(n805), .A2(G868), .ZN(n807) );
  INV_X1 U896 ( .A(n909), .ZN(n806) );
  XNOR2_X1 U897 ( .A(n807), .B(n806), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2078), .A2(G2084), .ZN(n808) );
  XOR2_X1 U899 ( .A(KEYINPUT20), .B(n808), .Z(n809) );
  NAND2_X1 U900 ( .A1(G2090), .A2(n809), .ZN(n811) );
  XNOR2_X1 U901 ( .A(KEYINPUT21), .B(KEYINPUT86), .ZN(n810) );
  XNOR2_X1 U902 ( .A(n811), .B(n810), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n812), .A2(G2072), .ZN(n813) );
  XOR2_X1 U904 ( .A(KEYINPUT87), .B(n813), .Z(G158) );
  XNOR2_X1 U905 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U906 ( .A1(G220), .A2(G219), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT22), .B(n814), .Z(n815) );
  NOR2_X1 U908 ( .A1(G218), .A2(n815), .ZN(n816) );
  XNOR2_X1 U909 ( .A(KEYINPUT88), .B(n816), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n817), .A2(G96), .ZN(n830) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n830), .ZN(n821) );
  NAND2_X1 U912 ( .A1(G120), .A2(G69), .ZN(n818) );
  NOR2_X1 U913 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U914 ( .A1(G108), .A2(n819), .ZN(n831) );
  NAND2_X1 U915 ( .A1(G567), .A2(n831), .ZN(n820) );
  NAND2_X1 U916 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U917 ( .A(KEYINPUT89), .B(n822), .ZN(G319) );
  INV_X1 U918 ( .A(G319), .ZN(n824) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n829) );
  NAND2_X1 U921 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U922 ( .A1(n825), .A2(G2106), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n826), .B(KEYINPUT110), .ZN(G217) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U925 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U927 ( .A1(n829), .A2(n828), .ZN(G188) );
  XNOR2_X1 U928 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U934 ( .A(G2430), .B(G2435), .ZN(n840) );
  XNOR2_X1 U935 ( .A(G2454), .B(KEYINPUT108), .ZN(n838) );
  XOR2_X1 U936 ( .A(G2451), .B(G2427), .Z(n833) );
  XNOR2_X1 U937 ( .A(G2438), .B(G2446), .ZN(n832) );
  XNOR2_X1 U938 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U939 ( .A(n834), .B(G2443), .Z(n836) );
  XNOR2_X1 U940 ( .A(G1341), .B(G1348), .ZN(n835) );
  XNOR2_X1 U941 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U942 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U943 ( .A(n840), .B(n839), .ZN(n841) );
  NAND2_X1 U944 ( .A1(n841), .A2(G14), .ZN(n842) );
  XNOR2_X1 U945 ( .A(KEYINPUT109), .B(n842), .ZN(G401) );
  XOR2_X1 U946 ( .A(G2474), .B(G1976), .Z(n844) );
  XNOR2_X1 U947 ( .A(G1961), .B(G1966), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U949 ( .A(n845), .B(KEYINPUT112), .Z(n847) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U952 ( .A(G1986), .B(G1981), .Z(n849) );
  XNOR2_X1 U953 ( .A(G1971), .B(G1956), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U955 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U956 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U957 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U958 ( .A(G2100), .B(G2096), .Z(n855) );
  XNOR2_X1 U959 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U960 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U961 ( .A(KEYINPUT43), .B(G2072), .Z(n857) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2090), .ZN(n856) );
  XNOR2_X1 U963 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U964 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U966 ( .A(n861), .B(n860), .ZN(G227) );
  NAND2_X1 U967 ( .A1(G124), .A2(n881), .ZN(n862) );
  XNOR2_X1 U968 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n887), .A2(G100), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U971 ( .A1(G136), .A2(n889), .ZN(n866) );
  NAND2_X1 U972 ( .A1(G112), .A2(n883), .ZN(n865) );
  NAND2_X1 U973 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U974 ( .A1(n868), .A2(n867), .ZN(G162) );
  XOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT120), .Z(n870) );
  XNOR2_X1 U976 ( .A(KEYINPUT119), .B(KEYINPUT46), .ZN(n869) );
  XNOR2_X1 U977 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U978 ( .A(n871), .B(KEYINPUT118), .Z(n880) );
  NAND2_X1 U979 ( .A1(G139), .A2(n889), .ZN(n873) );
  NAND2_X1 U980 ( .A1(G103), .A2(n887), .ZN(n872) );
  NAND2_X1 U981 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U982 ( .A1(G115), .A2(n883), .ZN(n875) );
  NAND2_X1 U983 ( .A1(G127), .A2(n881), .ZN(n874) );
  NAND2_X1 U984 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U986 ( .A1(n878), .A2(n877), .ZN(n945) );
  XNOR2_X1 U987 ( .A(n945), .B(KEYINPUT117), .ZN(n879) );
  XNOR2_X1 U988 ( .A(n880), .B(n879), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G130), .A2(n881), .ZN(n882) );
  XNOR2_X1 U990 ( .A(n882), .B(KEYINPUT114), .ZN(n886) );
  NAND2_X1 U991 ( .A1(G118), .A2(n883), .ZN(n884) );
  XOR2_X1 U992 ( .A(KEYINPUT115), .B(n884), .Z(n885) );
  NAND2_X1 U993 ( .A1(n886), .A2(n885), .ZN(n894) );
  NAND2_X1 U994 ( .A1(n887), .A2(G106), .ZN(n888) );
  XNOR2_X1 U995 ( .A(n888), .B(KEYINPUT116), .ZN(n891) );
  NAND2_X1 U996 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U997 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U998 ( .A(n892), .B(KEYINPUT45), .Z(n893) );
  NOR2_X1 U999 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U1000 ( .A(n896), .B(n895), .Z(n900) );
  XNOR2_X1 U1001 ( .A(G162), .B(n897), .ZN(n898) );
  XNOR2_X1 U1002 ( .A(n898), .B(n956), .ZN(n899) );
  XOR2_X1 U1003 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U1004 ( .A(G164), .B(G160), .ZN(n901) );
  XNOR2_X1 U1005 ( .A(n902), .B(n901), .ZN(n906) );
  XOR2_X1 U1006 ( .A(n904), .B(n903), .Z(n905) );
  XNOR2_X1 U1007 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n907), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(G171), .B(n910), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(n920), .B(n927), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1013 ( .A(n913), .B(G286), .ZN(n914) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n916), .ZN(n917) );
  AND2_X1 U1018 ( .A1(G319), .A2(n917), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1020 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1023 ( .A(G16), .B(KEYINPUT56), .Z(n942) );
  XNOR2_X1 U1024 ( .A(n920), .B(n981), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(G1971), .A2(G303), .ZN(n921) );
  NAND2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n924) );
  XNOR2_X1 U1027 ( .A(G1956), .B(G299), .ZN(n923) );
  NOR2_X1 U1028 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(G171), .B(G1961), .ZN(n929) );
  XNOR2_X1 U1031 ( .A(n927), .B(G1348), .ZN(n928) );
  NAND2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n933) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(G168), .B(G1966), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(n936), .B(KEYINPUT57), .ZN(n937) );
  NAND2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n969) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n961) );
  XOR2_X1 U1042 ( .A(G2072), .B(n945), .Z(n947) );
  XOR2_X1 U1043 ( .A(G164), .B(G2078), .Z(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT50), .B(n948), .ZN(n953) );
  XOR2_X1 U1046 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1048 ( .A(KEYINPUT51), .B(n951), .Z(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n959) );
  XOR2_X1 U1050 ( .A(G2084), .B(G160), .Z(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1056 ( .A(KEYINPUT52), .B(n964), .Z(n965) );
  NOR2_X1 U1057 ( .A1(KEYINPUT55), .A2(n965), .ZN(n967) );
  INV_X1 U1058 ( .A(G29), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1060 ( .A1(n969), .A2(n968), .ZN(n1025) );
  XOR2_X1 U1061 ( .A(G1976), .B(KEYINPUT126), .Z(n970) );
  XNOR2_X1 U1062 ( .A(G23), .B(n970), .ZN(n974) );
  XNOR2_X1 U1063 ( .A(G1971), .B(G22), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(G24), .B(G1986), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n975), .B(KEYINPUT58), .ZN(n979) );
  XOR2_X1 U1068 ( .A(n976), .B(G5), .Z(n977) );
  XNOR2_X1 U1069 ( .A(KEYINPUT124), .B(n977), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n992) );
  XNOR2_X1 U1071 ( .A(n980), .B(G20), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(n981), .B(G19), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n983), .A2(n982), .ZN(n989) );
  XOR2_X1 U1074 ( .A(G1981), .B(G6), .Z(n987) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(G4), .ZN(n984) );
  XOR2_X1 U1076 ( .A(n984), .B(G1348), .Z(n985) );
  XNOR2_X1 U1077 ( .A(n985), .B(KEYINPUT59), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(n990), .B(KEYINPUT60), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G21), .B(G1966), .ZN(n993) );
  NOR2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1084 ( .A(KEYINPUT61), .B(n995), .ZN(n997) );
  INV_X1 U1085 ( .A(G16), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n998), .A2(G11), .ZN(n1023) );
  XOR2_X1 U1088 ( .A(G29), .B(KEYINPUT123), .Z(n1021) );
  XNOR2_X1 U1089 ( .A(G27), .B(n999), .ZN(n1011) );
  XNOR2_X1 U1090 ( .A(G25), .B(G1991), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(n1000), .B(KEYINPUT121), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G26), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(G28), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G33), .B(G2072), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(G32), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT53), .B(n1012), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(G34), .B(KEYINPUT122), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(G2084), .B(KEYINPUT54), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(n1014), .B(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(G35), .B(G2090), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT55), .B(n1019), .Z(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1111 ( .A(KEYINPUT127), .B(n1026), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1027), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

