//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT67), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT70), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  OR4_X1    g030(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n455), .A2(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(G325), .B(KEYINPUT71), .ZN(G261));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT72), .B1(new_n463), .B2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT72), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n465), .A2(new_n466), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n466), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(new_n469), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n473), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(G2104), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G101), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n472), .A2(new_n478), .A3(new_n481), .ZN(G160));
  OR2_X1    g057(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n471), .A2(KEYINPUT73), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n464), .A2(new_n467), .A3(G2105), .A4(new_n469), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT74), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  MUX2_X1   g065(.A(G100), .B(G112), .S(G2105), .Z(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2104), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  AND3_X1   g069(.A1(new_n464), .A2(new_n467), .A3(new_n469), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT75), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G126), .A4(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT75), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  MUX2_X1   g074(.A(G102), .B(G114), .S(G2105), .Z(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2104), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n497), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT76), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n497), .A2(new_n499), .A3(new_n504), .A4(new_n501), .ZN(new_n505));
  INV_X1    g080(.A(G138), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n470), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g082(.A1(new_n506), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n474), .A3(new_n469), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n503), .A2(new_n505), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT77), .B1(new_n517), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n513), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n516), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n524), .A2(G62), .ZN(new_n529));
  NAND2_X1  g104(.A1(G75), .A2(G543), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT78), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n528), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(G166));
  AND2_X1   g108(.A1(new_n524), .A2(new_n513), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n515), .A2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n536), .A2(KEYINPUT79), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT79), .B1(new_n536), .B2(new_n537), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(G168));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT80), .B(G52), .Z(new_n545));
  OAI22_X1  g120(.A1(new_n525), .A2(new_n544), .B1(new_n514), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT81), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n528), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  AOI22_X1  g126(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n528), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n515), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n525), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n522), .A2(new_n523), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT82), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(KEYINPUT82), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(G651), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(G53), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n514), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n514), .B2(new_n571), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n534), .A2(G91), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  OAI21_X1  g152(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT83), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n534), .A2(G87), .B1(G49), .B2(new_n515), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n528), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n515), .A2(G48), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n525), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n584), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n534), .A2(G85), .B1(G47), .B2(new_n515), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n528), .B2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(new_n534), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT84), .B(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n565), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(G54), .B2(new_n515), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  MUX2_X1   g174(.A(new_n599), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g175(.A(new_n599), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g176(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g177(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g178(.A(new_n599), .ZN(new_n604));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n557), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(KEYINPUT85), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(KEYINPUT85), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n489), .A2(G123), .ZN(new_n613));
  NOR3_X1   g188(.A1(new_n468), .A2(KEYINPUT87), .A3(G111), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT87), .B1(new_n468), .B2(G111), .ZN(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(G2104), .A3(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n613), .B1(new_n614), .B2(new_n617), .C1(new_n485), .C2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(G2096), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(G2096), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n468), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT86), .B(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n620), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT88), .ZN(G156));
  INV_X1    g203(.A(KEYINPUT14), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2427), .ZN(new_n632));
  INV_X1    g207(.A(G2430), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT89), .B(KEYINPUT16), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n635), .A2(new_n642), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT90), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT17), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2084), .B(G2090), .ZN(new_n650));
  NOR3_X1   g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n650), .B1(new_n647), .B2(new_n649), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n648), .B2(new_n649), .ZN(new_n653));
  INV_X1    g228(.A(new_n649), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n654), .A2(new_n650), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT18), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n651), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2100), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(KEYINPUT92), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n667), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n664), .B2(new_n668), .ZN(new_n673));
  OR2_X1    g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1991), .B(G1996), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT93), .ZN(new_n680));
  XOR2_X1   g255(.A(G1981), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n678), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  NOR2_X1   g259(.A1(G16), .A2(G23), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n581), .B2(G16), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT98), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  NOR2_X1   g264(.A1(G6), .A2(G16), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n584), .A2(new_n587), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n690), .B1(new_n691), .B2(G16), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT97), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT32), .B(G1981), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(KEYINPUT96), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G22), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1971), .ZN(new_n703));
  NOR4_X1   g278(.A1(new_n689), .A2(new_n695), .A3(new_n696), .A4(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G25), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT94), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n486), .A2(G131), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT95), .ZN(new_n711));
  MUX2_X1   g286(.A(G95), .B(G107), .S(G2105), .Z(new_n712));
  AOI22_X1  g287(.A1(new_n489), .A2(G119), .B1(G2104), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n709), .B1(new_n714), .B2(G29), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT35), .B(G1991), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G24), .B(G290), .S(new_n700), .Z(new_n719));
  INV_X1    g294(.A(G1986), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n706), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n704), .A2(new_n705), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT36), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n707), .A2(G33), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n486), .A2(G139), .ZN(new_n727));
  NAND2_X1  g302(.A1(G115), .A2(G2104), .ZN(new_n728));
  INV_X1    g303(.A(G127), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n475), .B2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT25), .ZN(new_n731));
  INV_X1    g306(.A(G103), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n479), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n480), .A2(KEYINPUT25), .A3(G103), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n730), .A2(G2105), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n727), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n726), .B1(new_n737), .B2(new_n707), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(G2072), .Z(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  AND2_X1   g315(.A1(KEYINPUT24), .A2(G34), .ZN(new_n741));
  NOR2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n707), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G160), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n707), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n707), .A2(G32), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n486), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n489), .A2(G129), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT26), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(G105), .B2(new_n480), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n747), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n746), .B1(new_n755), .B2(new_n707), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT27), .B(G1996), .Z(new_n757));
  OAI221_X1 g332(.A(new_n739), .B1(new_n740), .B2(new_n745), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT100), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT29), .Z(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NOR2_X1   g340(.A1(G27), .A2(G29), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G164), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2078), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n764), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n697), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n697), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n772), .A2(G1966), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n700), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n557), .B2(new_n700), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1341), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n604), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G4), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n773), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n698), .A2(G20), .A3(new_n699), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n772), .A2(G1966), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT101), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n780), .A2(new_n784), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n778), .A2(new_n779), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n619), .A2(new_n707), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n745), .A2(new_n740), .ZN(new_n790));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G11), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT30), .B(G28), .Z(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G29), .ZN(new_n793));
  NOR4_X1   g368(.A1(new_n788), .A2(new_n789), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n707), .A2(G26), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT28), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n489), .A2(G128), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  MUX2_X1   g373(.A(G104), .B(G116), .S(G2105), .Z(new_n799));
  AOI22_X1  g374(.A1(new_n486), .A2(G140), .B1(G2104), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n796), .B1(new_n801), .B2(G29), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n697), .A2(G5), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G171), .B2(new_n697), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(G1961), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n805), .A2(G1961), .B1(new_n756), .B2(new_n757), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n794), .A2(new_n803), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n759), .A2(new_n770), .A3(new_n787), .A4(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n725), .A2(new_n810), .ZN(G311));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n724), .B(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(new_n809), .ZN(G150));
  AOI22_X1  g389(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT102), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(G651), .A3(new_n817), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n534), .A2(G93), .B1(G55), .B2(new_n515), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G860), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  INV_X1    g397(.A(new_n557), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n818), .A2(new_n557), .A3(new_n819), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT38), .Z(new_n827));
  NOR2_X1   g402(.A1(new_n599), .A2(new_n605), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(G860), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(new_n830), .B2(KEYINPUT39), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n822), .B1(new_n831), .B2(new_n833), .ZN(G145));
  INV_X1    g409(.A(KEYINPUT105), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n489), .A2(G130), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT103), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n468), .A2(G106), .ZN(new_n839));
  NAND2_X1  g414(.A1(G118), .A2(G2105), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n463), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n486), .B2(G142), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n623), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n714), .A2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n714), .A2(new_n845), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n844), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n711), .A2(new_n713), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(new_n623), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n851), .A2(new_n843), .A3(new_n846), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n801), .B(new_n736), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n510), .A2(new_n499), .A3(new_n497), .A4(new_n501), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n754), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n835), .B1(new_n853), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n493), .B(new_n744), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n619), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n853), .B2(new_n860), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n849), .A2(new_n859), .A3(KEYINPUT105), .A4(new_n852), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT106), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT106), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n861), .A2(new_n864), .A3(new_n868), .A4(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT104), .B1(new_n853), .B2(new_n860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n853), .A2(new_n860), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n849), .A2(new_n859), .A3(new_n873), .A4(new_n852), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G37), .B1(new_n875), .B2(new_n863), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g453(.A1(new_n820), .A2(G868), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G299), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n599), .A2(new_n881), .A3(KEYINPUT107), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT107), .B1(new_n599), .B2(new_n881), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n882), .A2(new_n883), .B1(new_n881), .B2(new_n599), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n607), .B(new_n826), .Z(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n581), .B(G290), .Z(new_n891));
  XNOR2_X1  g466(.A(new_n691), .B(G166), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n891), .B(new_n892), .Z(new_n893));
  NAND2_X1  g468(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(new_n887), .B2(new_n884), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n882), .A2(new_n883), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n599), .A2(new_n881), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n888), .A2(new_n900), .A3(KEYINPUT108), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n890), .A2(new_n895), .A3(new_n897), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n897), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n893), .B(new_n894), .C1(new_n903), .C2(new_n889), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n904), .B(new_n902), .C1(KEYINPUT109), .C2(KEYINPUT42), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G868), .ZN(new_n910));
  OAI211_X1 g485(.A(KEYINPUT110), .B(new_n880), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(new_n879), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n911), .A2(new_n914), .ZN(G295));
  NOR2_X1   g490(.A1(new_n913), .A2(new_n879), .ZN(G331));
  XNOR2_X1  g491(.A(G301), .B(G286), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n917), .A2(new_n826), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n826), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n884), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n886), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n923), .B2(new_n893), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n900), .A2(KEYINPUT41), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n884), .A2(new_n885), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n922), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n920), .ZN(new_n928));
  INV_X1    g503(.A(new_n893), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT111), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n931));
  AOI211_X1 g506(.A(new_n931), .B(new_n893), .C1(new_n927), .C2(new_n920), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n924), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n924), .B(new_n935), .C1(new_n930), .C2(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n937), .B(KEYINPUT44), .Z(G397));
  NOR2_X1   g513(.A1(new_n850), .A2(new_n716), .ZN(new_n939));
  INV_X1    g514(.A(G2067), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n801), .B(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1996), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n754), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n714), .A2(new_n717), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n939), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(G290), .B(new_n720), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n855), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G160), .A2(G40), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n948), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT125), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT116), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n502), .A2(KEYINPUT76), .B1(new_n507), .B2(new_n509), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n960), .B2(new_n505), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT50), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n511), .A2(new_n949), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n964), .A2(KEYINPUT116), .A3(KEYINPUT50), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n509), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n464), .A2(new_n469), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(G138), .A3(new_n468), .A4(new_n467), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n969), .B2(KEYINPUT4), .ZN(new_n970));
  OAI211_X1 g545(.A(KEYINPUT115), .B(new_n949), .C1(new_n502), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT115), .B1(new_n855), .B2(new_n949), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n955), .B1(new_n974), .B2(new_n962), .ZN(new_n975));
  XOR2_X1   g550(.A(KEYINPUT121), .B(G2084), .Z(new_n976));
  NAND3_X1  g551(.A1(new_n966), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT123), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n972), .B2(new_n973), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n961), .A2(new_n953), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n956), .ZN(new_n982));
  INV_X1    g557(.A(G1966), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n977), .A2(new_n978), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n978), .B1(new_n977), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  NOR2_X1   g563(.A1(G168), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT124), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n992), .B(G8), .C1(new_n985), .C2(new_n986), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n977), .A2(new_n984), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT123), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n977), .A2(new_n978), .A3(new_n984), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n992), .B1(new_n998), .B2(G8), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT51), .B1(new_n994), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n990), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n991), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G305), .A2(G1981), .ZN(new_n1005));
  OR3_X1    g580(.A1(new_n584), .A2(new_n587), .A3(G1981), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT49), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n974), .A2(new_n956), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1005), .A2(KEYINPUT49), .A3(new_n1006), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(G8), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT119), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1010), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G288), .A2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1014), .A2(new_n1016), .A3(new_n988), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1017), .B(new_n1018), .C1(G1976), .C2(new_n581), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1013), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(G303), .A2(G8), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n1022), .B(KEYINPUT55), .Z(new_n1023));
  XOR2_X1   g598(.A(KEYINPUT113), .B(G1971), .Z(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n961), .A2(new_n953), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n956), .B1(new_n950), .B2(new_n979), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(KEYINPUT50), .B2(new_n961), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n956), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT117), .B(G2090), .Z(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1028), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1023), .B1(new_n1034), .B2(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1021), .A2(new_n1035), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n966), .A2(new_n975), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1028), .A2(KEYINPUT114), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1039), .B(new_n1025), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1037), .A2(new_n1032), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n988), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n966), .A2(new_n975), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1045), .B2(new_n1033), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(KEYINPUT118), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1043), .A2(new_n1047), .A3(new_n1023), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT53), .B1(new_n1049), .B2(new_n768), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1045), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n982), .A2(new_n1053), .A3(G2078), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(G301), .B(KEYINPUT54), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1027), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n954), .A2(new_n1053), .A3(G2078), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1055), .A2(new_n1056), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1036), .A2(new_n1048), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n958), .B1(new_n1004), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1003), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT124), .B1(new_n987), .B2(new_n988), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(new_n993), .A3(new_n990), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1064), .B1(new_n1066), .B2(KEYINPUT51), .ZN(new_n1067));
  OAI211_X1 g642(.A(KEYINPUT125), .B(new_n1063), .C1(new_n1067), .C2(new_n991), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT56), .B(G2072), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1031), .A2(new_n1069), .B1(new_n1049), .B2(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(G299), .B(KEYINPUT57), .Z(new_n1072));
  NOR2_X1   g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1045), .A2(new_n779), .B1(new_n940), .B2(new_n1014), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(new_n599), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1073), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1076), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1073), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  AOI22_X1  g656(.A1(new_n1049), .A2(new_n942), .B1(new_n1010), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n823), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1083), .B(KEYINPUT59), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1084), .B1(new_n1074), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1079), .B1(new_n1078), .B2(new_n1073), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1080), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1075), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1074), .A2(new_n599), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1077), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1062), .A2(new_n1068), .A3(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1013), .A2(new_n1015), .A3(new_n581), .ZN(new_n1095));
  XOR2_X1   g670(.A(new_n1006), .B(KEYINPUT120), .Z(new_n1096));
  OAI211_X1 g671(.A(G8), .B(new_n1010), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1048), .B2(new_n1021), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1023), .ZN(new_n1099));
  OAI21_X1  g674(.A(G8), .B1(new_n1046), .B2(KEYINPUT118), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1021), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(KEYINPUT122), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1023), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1021), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT63), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1001), .A2(new_n1108), .A3(G286), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1048), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1104), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1001), .A2(G286), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1036), .A2(new_n1048), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1108), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1098), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n1116));
  INV_X1    g691(.A(new_n991), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n988), .B1(new_n996), .B2(new_n997), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n989), .B1(new_n1118), .B2(new_n992), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1002), .B1(new_n1119), .B2(new_n1065), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1116), .B(new_n1117), .C1(new_n1120), .C2(new_n1064), .ZN(new_n1121));
  AND4_X1   g696(.A1(G171), .A2(new_n1036), .A3(new_n1048), .A4(new_n1055), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1004), .A2(new_n1116), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1115), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n957), .B1(new_n1094), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n954), .A2(new_n956), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n941), .B2(new_n755), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT46), .B1(new_n1127), .B2(G1996), .ZN(new_n1129));
  OR3_X1    g704(.A1(new_n1127), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT47), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n946), .A2(new_n1127), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1127), .A2(G1986), .A3(G290), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1134), .B(KEYINPUT48), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n945), .A2(new_n941), .A3(new_n943), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n798), .A2(new_n940), .A3(new_n800), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1127), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1133), .A2(new_n1135), .B1(new_n1138), .B2(KEYINPUT126), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1132), .B(new_n1139), .C1(KEYINPUT126), .C2(new_n1138), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1126), .A2(new_n1140), .ZN(G329));
  assign    G231 = 1'b0;
  OR4_X1    g716(.A1(new_n461), .A2(G227), .A3(G229), .A4(G401), .ZN(new_n1143));
  AOI21_X1  g717(.A(new_n1143), .B1(new_n870), .B2(new_n876), .ZN(new_n1144));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n1145));
  AND3_X1   g719(.A1(new_n937), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n937), .B2(new_n1144), .ZN(new_n1147));
  NOR2_X1   g721(.A1(new_n1146), .A2(new_n1147), .ZN(G308));
  NAND2_X1  g722(.A1(new_n937), .A2(new_n1144), .ZN(G225));
endmodule


