

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  XNOR2_X1 U321 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U322 ( .A(n377), .B(n290), .ZN(n378) );
  NOR2_X1 U323 ( .A1(n466), .A2(n508), .ZN(n565) );
  XNOR2_X1 U324 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n417) );
  XNOR2_X1 U325 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U326 ( .A(n467), .B(KEYINPUT28), .Z(n521) );
  XOR2_X1 U327 ( .A(n369), .B(n368), .Z(n508) );
  AND2_X1 U328 ( .A1(G228GAT), .A2(G233GAT), .ZN(n289) );
  XOR2_X1 U329 ( .A(n376), .B(n375), .Z(n290) );
  XOR2_X1 U330 ( .A(G99GAT), .B(G85GAT), .Z(n438) );
  XNOR2_X1 U331 ( .A(n370), .B(n289), .ZN(n371) );
  XNOR2_X1 U332 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U333 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U334 ( .A(n334), .B(KEYINPUT10), .ZN(n335) );
  XNOR2_X1 U335 ( .A(n336), .B(n335), .ZN(n339) );
  XNOR2_X1 U336 ( .A(n418), .B(n417), .ZN(n505) );
  XNOR2_X1 U337 ( .A(n405), .B(KEYINPUT26), .ZN(n564) );
  INV_X1 U338 ( .A(n564), .ZN(n537) );
  XOR2_X1 U339 ( .A(n446), .B(n445), .Z(n571) );
  XNOR2_X1 U340 ( .A(n345), .B(n344), .ZN(n546) );
  XNOR2_X1 U341 ( .A(n448), .B(n447), .ZN(n493) );
  XNOR2_X1 U342 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n449) );
  XNOR2_X1 U344 ( .A(n474), .B(n473), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n450), .B(n449), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n292) );
  XNOR2_X1 U347 ( .A(KEYINPUT81), .B(G183GAT), .ZN(n291) );
  XNOR2_X1 U348 ( .A(n292), .B(n291), .ZN(n311) );
  XOR2_X1 U349 ( .A(G99GAT), .B(G134GAT), .Z(n294) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U352 ( .A(KEYINPUT65), .B(G176GAT), .Z(n296) );
  XNOR2_X1 U353 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U355 ( .A(n298), .B(n297), .Z(n309) );
  XNOR2_X1 U356 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n299), .B(KEYINPUT17), .ZN(n300) );
  XOR2_X1 U358 ( .A(n300), .B(KEYINPUT82), .Z(n302) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n400) );
  XOR2_X1 U361 ( .A(G120GAT), .B(G127GAT), .Z(n304) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n361) );
  XOR2_X1 U364 ( .A(n361), .B(G71GAT), .Z(n306) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n400), .B(n307), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U369 ( .A(n311), .B(n310), .Z(n412) );
  INV_X1 U370 ( .A(n412), .ZN(n549) );
  XOR2_X1 U371 ( .A(G8GAT), .B(G183GAT), .Z(n388) );
  XOR2_X1 U372 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n313) );
  XNOR2_X1 U373 ( .A(KEYINPUT78), .B(KEYINPUT14), .ZN(n312) );
  XNOR2_X1 U374 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U375 ( .A(n388), .B(n314), .Z(n317) );
  XNOR2_X1 U376 ( .A(G15GAT), .B(G1GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n315), .B(KEYINPUT69), .ZN(n419) );
  XOR2_X1 U378 ( .A(G22GAT), .B(G155GAT), .Z(n370) );
  XNOR2_X1 U379 ( .A(n419), .B(n370), .ZN(n316) );
  XNOR2_X1 U380 ( .A(n317), .B(n316), .ZN(n327) );
  XOR2_X1 U381 ( .A(KEYINPUT76), .B(G64GAT), .Z(n319) );
  XNOR2_X1 U382 ( .A(G127GAT), .B(G211GAT), .ZN(n318) );
  XNOR2_X1 U383 ( .A(n319), .B(n318), .ZN(n325) );
  XOR2_X1 U384 ( .A(KEYINPUT13), .B(G57GAT), .Z(n321) );
  XNOR2_X1 U385 ( .A(G71GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n321), .B(n320), .ZN(n442) );
  XOR2_X1 U387 ( .A(n442), .B(KEYINPUT12), .Z(n323) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U389 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U390 ( .A(n325), .B(n324), .Z(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n574) );
  XOR2_X1 U392 ( .A(KEYINPUT73), .B(KEYINPUT66), .Z(n329) );
  XNOR2_X1 U393 ( .A(KEYINPUT9), .B(G92GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U395 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n331) );
  XOR2_X1 U396 ( .A(G134GAT), .B(KEYINPUT74), .Z(n360) );
  XNOR2_X1 U397 ( .A(n360), .B(n438), .ZN(n330) );
  XNOR2_X1 U398 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n336) );
  AND2_X1 U400 ( .A1(G232GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U401 ( .A(G36GAT), .B(G190GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n337), .B(G218GAT), .ZN(n392) );
  XOR2_X1 U403 ( .A(n392), .B(KEYINPUT67), .Z(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n345) );
  XOR2_X1 U405 ( .A(G29GAT), .B(G43GAT), .Z(n341) );
  XNOR2_X1 U406 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n340) );
  XNOR2_X1 U407 ( .A(n341), .B(n340), .ZN(n432) );
  XOR2_X1 U408 ( .A(G106GAT), .B(G162GAT), .Z(n343) );
  XNOR2_X1 U409 ( .A(G50GAT), .B(KEYINPUT72), .ZN(n342) );
  XNOR2_X1 U410 ( .A(n343), .B(n342), .ZN(n374) );
  XOR2_X1 U411 ( .A(n432), .B(n374), .Z(n344) );
  INV_X1 U412 ( .A(KEYINPUT102), .ZN(n346) );
  XNOR2_X1 U413 ( .A(n546), .B(n346), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n347), .B(KEYINPUT36), .ZN(n578) );
  XOR2_X1 U415 ( .A(G57GAT), .B(KEYINPUT5), .Z(n349) );
  XNOR2_X1 U416 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n348) );
  XNOR2_X1 U417 ( .A(n349), .B(n348), .ZN(n369) );
  XOR2_X1 U418 ( .A(KEYINPUT90), .B(KEYINPUT4), .Z(n351) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(G155GAT), .ZN(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U421 ( .A(KEYINPUT1), .B(KEYINPUT92), .Z(n353) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n352) );
  XNOR2_X1 U423 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U424 ( .A(n355), .B(n354), .Z(n367) );
  XOR2_X1 U425 ( .A(G148GAT), .B(KEYINPUT3), .Z(n357) );
  XNOR2_X1 U426 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n356) );
  XNOR2_X1 U427 ( .A(n357), .B(n356), .ZN(n372) );
  XOR2_X1 U428 ( .A(n372), .B(KEYINPUT94), .Z(n359) );
  NAND2_X1 U429 ( .A1(G225GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U430 ( .A(n359), .B(n358), .ZN(n365) );
  XOR2_X1 U431 ( .A(G85GAT), .B(n360), .Z(n363) );
  XNOR2_X1 U432 ( .A(n361), .B(G162GAT), .ZN(n362) );
  XNOR2_X1 U433 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U434 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U435 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U436 ( .A(n373), .B(KEYINPUT24), .Z(n379) );
  XNOR2_X1 U437 ( .A(n374), .B(KEYINPUT87), .ZN(n377) );
  XOR2_X1 U438 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n376) );
  XNOR2_X1 U439 ( .A(G218GAT), .B(KEYINPUT84), .ZN(n375) );
  XOR2_X1 U440 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n381) );
  XNOR2_X1 U441 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U443 ( .A(G197GAT), .B(n382), .Z(n389) );
  XOR2_X1 U444 ( .A(KEYINPUT89), .B(G78GAT), .Z(n384) );
  XNOR2_X1 U445 ( .A(KEYINPUT88), .B(G204GAT), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n389), .B(n385), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n467) );
  XOR2_X1 U449 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n391) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n396) );
  XOR2_X1 U452 ( .A(n392), .B(KEYINPUT97), .Z(n394) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U454 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U455 ( .A(n396), .B(n395), .Z(n402) );
  XOR2_X1 U456 ( .A(KEYINPUT71), .B(G64GAT), .Z(n398) );
  XNOR2_X1 U457 ( .A(G204GAT), .B(G92GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U459 ( .A(G176GAT), .B(n399), .Z(n445) );
  XNOR2_X1 U460 ( .A(n400), .B(n445), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n510) );
  NAND2_X1 U462 ( .A1(n510), .A2(n549), .ZN(n403) );
  NAND2_X1 U463 ( .A1(n467), .A2(n403), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n404), .B(KEYINPUT25), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n510), .B(KEYINPUT27), .ZN(n410) );
  NOR2_X1 U466 ( .A1(n467), .A2(n549), .ZN(n405) );
  AND2_X1 U467 ( .A1(n410), .A2(n564), .ZN(n406) );
  NOR2_X1 U468 ( .A1(n407), .A2(n406), .ZN(n408) );
  NOR2_X1 U469 ( .A1(n508), .A2(n408), .ZN(n409) );
  XOR2_X1 U470 ( .A(KEYINPUT99), .B(n409), .Z(n415) );
  NAND2_X1 U471 ( .A1(n410), .A2(n508), .ZN(n411) );
  XOR2_X1 U472 ( .A(KEYINPUT98), .B(n411), .Z(n518) );
  NAND2_X1 U473 ( .A1(n412), .A2(n518), .ZN(n413) );
  NOR2_X1 U474 ( .A1(n521), .A2(n413), .ZN(n414) );
  NOR2_X1 U475 ( .A1(n415), .A2(n414), .ZN(n476) );
  NOR2_X1 U476 ( .A1(n578), .A2(n476), .ZN(n416) );
  NAND2_X1 U477 ( .A1(n574), .A2(n416), .ZN(n418) );
  XOR2_X1 U478 ( .A(G50GAT), .B(n419), .Z(n421) );
  NAND2_X1 U479 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U481 ( .A(n422), .B(G36GAT), .Z(n430) );
  XOR2_X1 U482 ( .A(G141GAT), .B(G197GAT), .Z(n424) );
  XNOR2_X1 U483 ( .A(G169GAT), .B(G22GAT), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U485 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n426) );
  XNOR2_X1 U486 ( .A(G113GAT), .B(G8GAT), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n431), .B(KEYINPUT68), .Z(n434) );
  XNOR2_X1 U491 ( .A(n432), .B(KEYINPUT70), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n548) );
  XOR2_X1 U493 ( .A(KEYINPUT31), .B(G148GAT), .Z(n436) );
  XNOR2_X1 U494 ( .A(G120GAT), .B(G106GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n440) );
  AND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n437) );
  XOR2_X1 U497 ( .A(KEYINPUT32), .B(n441), .Z(n444) );
  XNOR2_X1 U498 ( .A(n442), .B(KEYINPUT33), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n446) );
  NAND2_X1 U500 ( .A1(n548), .A2(n571), .ZN(n479) );
  OR2_X1 U501 ( .A1(n505), .A2(n479), .ZN(n448) );
  XOR2_X1 U502 ( .A(KEYINPUT104), .B(KEYINPUT38), .Z(n447) );
  NAND2_X1 U503 ( .A1(n549), .A2(n493), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n571), .B(KEYINPUT64), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n451), .B(KEYINPUT41), .ZN(n558) );
  NAND2_X1 U506 ( .A1(n548), .A2(n558), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n452), .B(KEYINPUT46), .ZN(n453) );
  XNOR2_X1 U508 ( .A(KEYINPUT110), .B(n574), .ZN(n562) );
  NAND2_X1 U509 ( .A1(n453), .A2(n562), .ZN(n454) );
  NOR2_X1 U510 ( .A1(n454), .A2(n546), .ZN(n456) );
  XNOR2_X1 U511 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n455) );
  XNOR2_X1 U512 ( .A(n456), .B(n455), .ZN(n461) );
  NOR2_X1 U513 ( .A1(n578), .A2(n574), .ZN(n457) );
  XNOR2_X1 U514 ( .A(KEYINPUT45), .B(n457), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n458), .A2(n571), .ZN(n459) );
  NOR2_X1 U516 ( .A1(n548), .A2(n459), .ZN(n460) );
  NOR2_X1 U517 ( .A1(n461), .A2(n460), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT48), .ZN(n517) );
  XOR2_X1 U519 ( .A(KEYINPUT118), .B(n510), .Z(n463) );
  NOR2_X1 U520 ( .A1(n517), .A2(n463), .ZN(n465) );
  INV_X1 U521 ( .A(KEYINPUT54), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n565), .A2(n467), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n468) );
  XNOR2_X1 U525 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT55), .ZN(n551) );
  NAND2_X1 U527 ( .A1(n551), .A2(n549), .ZN(n561) );
  INV_X1 U528 ( .A(n561), .ZN(n557) );
  NAND2_X1 U529 ( .A1(n557), .A2(n546), .ZN(n474) );
  XOR2_X1 U530 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n472) );
  XNOR2_X1 U531 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n471) );
  XNOR2_X1 U532 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n481) );
  NOR2_X1 U533 ( .A1(n546), .A2(n574), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT16), .ZN(n478) );
  INV_X1 U535 ( .A(n476), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n495) );
  NOR2_X1 U537 ( .A1(n479), .A2(n495), .ZN(n487) );
  NAND2_X1 U538 ( .A1(n508), .A2(n487), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U540 ( .A1(n487), .A2(n510), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n484) );
  NAND2_X1 U543 ( .A1(n487), .A2(n549), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(n486) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT100), .Z(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U547 ( .A1(n487), .A2(n521), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U549 ( .A1(n493), .A2(n508), .ZN(n491) );
  XNOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n493), .A2(n510), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U555 ( .A1(n493), .A2(n521), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n494), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n498) );
  INV_X1 U558 ( .A(n548), .ZN(n566) );
  NAND2_X1 U559 ( .A1(n558), .A2(n566), .ZN(n506) );
  NOR2_X1 U560 ( .A1(n506), .A2(n495), .ZN(n496) );
  XNOR2_X1 U561 ( .A(KEYINPUT106), .B(n496), .ZN(n502) );
  NAND2_X1 U562 ( .A1(n508), .A2(n502), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U565 ( .A1(n502), .A2(n510), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U567 ( .A1(n502), .A2(n549), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n501), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(G78GAT), .B(KEYINPUT43), .Z(n504) );
  NAND2_X1 U570 ( .A1(n521), .A2(n502), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n504), .B(n503), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n506), .A2(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(KEYINPUT108), .ZN(n513) );
  NAND2_X1 U574 ( .A1(n513), .A2(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n510), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n513), .A2(n549), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n515) );
  NAND2_X1 U581 ( .A1(n521), .A2(n513), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n516), .ZN(G1339GAT) );
  INV_X1 U584 ( .A(n517), .ZN(n519) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U586 ( .A(KEYINPUT112), .B(n520), .ZN(n536) );
  NOR2_X1 U587 ( .A1(n521), .A2(n536), .ZN(n522) );
  NAND2_X1 U588 ( .A1(n522), .A2(n549), .ZN(n523) );
  XNOR2_X1 U589 ( .A(KEYINPUT113), .B(n523), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n548), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT114), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n527) );
  NAND2_X1 U594 ( .A1(n533), .A2(n558), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U596 ( .A(G120GAT), .B(n528), .Z(G1341GAT) );
  INV_X1 U597 ( .A(n533), .ZN(n529) );
  NOR2_X1 U598 ( .A1(n562), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n532), .Z(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n535) );
  NAND2_X1 U603 ( .A1(n533), .A2(n546), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n548), .A2(n545), .ZN(n538) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n538), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n540) );
  NAND2_X1 U609 ( .A1(n545), .A2(n558), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(n541), .ZN(G1345GAT) );
  XOR2_X1 U612 ( .A(G155GAT), .B(KEYINPUT117), .Z(n544) );
  INV_X1 U613 ( .A(n574), .ZN(n542) );
  NAND2_X1 U614 ( .A1(n545), .A2(n542), .ZN(n543) );
  XNOR2_X1 U615 ( .A(n544), .B(n543), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n547), .B(G162GAT), .ZN(G1347GAT) );
  AND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U620 ( .A(n552), .B(KEYINPUT121), .Z(n553) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n555) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U624 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(n556), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n563), .Z(G1350GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n566), .A2(n577), .ZN(n570) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n577), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n577), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U643 ( .A(KEYINPUT62), .B(n579), .Z(n580) );
  XNOR2_X1 U644 ( .A(G218GAT), .B(n580), .ZN(G1355GAT) );
endmodule

