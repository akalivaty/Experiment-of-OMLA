//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n194), .B2(new_n188), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n195), .B(G146), .ZN(new_n196));
  INV_X1    g010(.A(G237), .ZN(new_n197));
  INV_X1    g011(.A(G953), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G214), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n197), .A2(new_n198), .A3(G143), .A4(G214), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT17), .A3(G131), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT90), .B1(new_n203), .B2(G131), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT90), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n201), .A2(new_n207), .A3(new_n208), .A4(new_n202), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n196), .B(new_n204), .C1(new_n210), .C2(KEYINPUT17), .ZN(new_n211));
  XNOR2_X1  g025(.A(G113), .B(G122), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n212), .B(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT18), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n201), .B(new_n202), .C1(new_n215), .C2(new_n208), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n216), .B(KEYINPUT89), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n191), .A2(new_n193), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT88), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n194), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(G146), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n215), .A2(new_n208), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n222), .A2(new_n224), .B1(new_n203), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n211), .A2(new_n214), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n195), .A2(new_n223), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(KEYINPUT19), .A3(new_n221), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(KEYINPUT19), .B2(new_n194), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n210), .B(new_n230), .C1(new_n232), .C2(G146), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n214), .B1(new_n233), .B2(new_n227), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n187), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n236), .A2(KEYINPUT20), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(KEYINPUT20), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n233), .A2(new_n227), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n228), .B1(new_n240), .B2(new_n214), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n241), .A2(new_n236), .A3(KEYINPUT20), .A4(new_n187), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n214), .B1(new_n211), .B2(new_n227), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n229), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G475), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n239), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n200), .A2(G128), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G128), .B2(new_n200), .ZN(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n252), .A2(KEYINPUT93), .A3(G143), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n249), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT95), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(KEYINPUT95), .B(new_n249), .C1(new_n251), .C2(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  INV_X1    g073(.A(G107), .ZN(new_n260));
  INV_X1    g074(.A(G122), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G116), .ZN(new_n262));
  INV_X1    g076(.A(G116), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G122), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT92), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G116), .B(G122), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(KEYINPUT92), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n260), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n265), .A2(new_n266), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(KEYINPUT92), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G107), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n258), .A2(new_n259), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT13), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n251), .B2(new_n253), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT94), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(new_n249), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT93), .B1(new_n252), .B2(G143), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n250), .A2(new_n200), .A3(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT13), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT94), .B1(new_n281), .B2(new_n248), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT13), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n278), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G134), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n274), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n264), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n260), .B1(new_n287), .B2(KEYINPUT14), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n288), .B1(KEYINPUT14), .B2(new_n265), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n256), .A2(G134), .A3(new_n257), .ZN(new_n290));
  AOI21_X1  g104(.A(G134), .B1(new_n256), .B2(new_n257), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n270), .B(new_n289), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT9), .B(G234), .ZN(new_n293));
  INV_X1    g107(.A(G217), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(new_n294), .A3(G953), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n286), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n286), .B2(new_n292), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n243), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT96), .ZN(new_n299));
  INV_X1    g113(.A(G478), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT15), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT96), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n302), .B(new_n243), .C1(new_n296), .C2(new_n297), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n298), .A2(new_n301), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT97), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT97), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n304), .A2(new_n308), .A3(new_n305), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n247), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G140), .ZN(new_n311));
  INV_X1    g125(.A(G227), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n312), .A2(G953), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n311), .B(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G101), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n260), .A2(G104), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n213), .A2(G107), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT80), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT1), .B1(new_n200), .B2(G146), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n200), .A2(G146), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n223), .A2(G143), .ZN(new_n323));
  OAI211_X1 g137(.A(G128), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n223), .A2(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n200), .A2(G146), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n325), .B(new_n326), .C1(KEYINPUT1), .C2(new_n252), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT3), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n260), .A3(G104), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n330), .A2(new_n332), .A3(new_n316), .A4(new_n318), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n320), .A2(new_n329), .A3(KEYINPUT10), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT0), .A2(G128), .ZN(new_n335));
  OR2_X1    g149(.A1(KEYINPUT0), .A2(G128), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n335), .B(new_n336), .C1(new_n322), .C2(new_n323), .ZN(new_n337));
  AND2_X1   g151(.A1(KEYINPUT0), .A2(G128), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n325), .A2(new_n326), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n330), .A2(new_n332), .A3(new_n318), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G101), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n342), .A2(G101), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n333), .A2(KEYINPUT4), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n341), .B(new_n344), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n334), .A2(new_n347), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n317), .A2(new_n318), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT80), .B1(new_n349), .B2(new_n316), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n319), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n333), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT81), .B1(new_n353), .B2(new_n328), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n320), .A2(new_n329), .A3(new_n355), .A4(new_n333), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G137), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G134), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT11), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(G134), .B2(new_n359), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n259), .A2(KEYINPUT11), .A3(G137), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n208), .B(new_n361), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT65), .ZN(new_n366));
  OAI21_X1  g180(.A(KEYINPUT11), .B1(new_n259), .B2(G137), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n362), .A2(new_n359), .A3(G134), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n360), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT65), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n208), .ZN(new_n371));
  INV_X1    g185(.A(new_n369), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n366), .A2(new_n371), .B1(G131), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n348), .A2(new_n358), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n353), .A2(new_n328), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n354), .A2(new_n356), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n372), .A2(G131), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n367), .A2(new_n368), .ZN(new_n378));
  AND4_X1   g192(.A1(new_n370), .A2(new_n378), .A3(new_n208), .A4(new_n361), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n370), .B1(new_n369), .B2(new_n208), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n376), .A2(KEYINPUT12), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT12), .B1(new_n376), .B2(new_n381), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n315), .B(new_n374), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n374), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n373), .B1(new_n348), .B2(new_n358), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n314), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G469), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(new_n243), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n374), .A2(new_n315), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n392), .A2(new_n387), .ZN(new_n393));
  INV_X1    g207(.A(new_n384), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n386), .B1(new_n382), .B2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n393), .B(G469), .C1(new_n395), .C2(new_n315), .ZN(new_n396));
  NAND2_X1  g210(.A1(G469), .A2(G902), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(G221), .B1(new_n293), .B2(G902), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n340), .A2(G125), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n328), .A2(new_n192), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT83), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n340), .A2(new_n404), .A3(G125), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n198), .A2(G224), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n407), .B(KEYINPUT84), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n406), .B(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G119), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G116), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n263), .A2(G119), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT2), .B(G113), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT5), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n417), .B(G113), .C1(KEYINPUT5), .C2(new_n412), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n320), .A2(new_n333), .A3(new_n416), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n415), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(new_n344), .C1(new_n345), .C2(new_n346), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G122), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n419), .A2(new_n422), .A3(new_n424), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n429), .A3(new_n425), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n410), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n418), .A2(new_n416), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n353), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n419), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n424), .B(KEYINPUT8), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n405), .A2(new_n403), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n437), .A2(KEYINPUT7), .A3(new_n408), .A4(new_n402), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n403), .A2(new_n401), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT85), .B(KEYINPUT7), .Z(new_n440));
  NAND2_X1  g254(.A1(new_n408), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n436), .A2(new_n438), .A3(KEYINPUT86), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n427), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n434), .A2(new_n435), .B1(new_n439), .B2(new_n441), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT86), .B1(new_n445), .B2(new_n438), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n431), .B(new_n243), .C1(new_n444), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n448), .B(KEYINPUT87), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G214), .B1(G237), .B2(G902), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n452), .B(KEYINPUT82), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n436), .A2(new_n438), .A3(new_n442), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n427), .A3(new_n443), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n458), .A2(new_n243), .A3(new_n449), .A4(new_n431), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(new_n454), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G952), .ZN(new_n462));
  AOI211_X1 g276(.A(G953), .B(new_n462), .C1(G234), .C2(G237), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n243), .B(new_n198), .C1(G234), .C2(G237), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  XOR2_X1   g280(.A(KEYINPUT21), .B(G898), .Z(new_n467));
  OAI21_X1  g281(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND4_X1   g282(.A1(new_n310), .A2(new_n400), .A3(new_n461), .A4(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT70), .ZN(new_n470));
  NOR2_X1   g284(.A1(G472), .A2(G902), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n421), .B1(new_n381), .B2(new_n341), .ZN(new_n473));
  AOI21_X1  g287(.A(KEYINPUT66), .B1(new_n259), .B2(G137), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n259), .A2(G137), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n360), .A2(KEYINPUT66), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n208), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n366), .B2(new_n371), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n329), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n477), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G131), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n379), .B2(new_n380), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n473), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n197), .A2(new_n198), .A3(G210), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT27), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G101), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n488), .B(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT64), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n336), .A2(new_n335), .ZN(new_n493));
  XNOR2_X1  g307(.A(G143), .B(G146), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n339), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n492), .B1(new_n337), .B2(new_n339), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n381), .A2(new_n498), .B1(new_n479), .B2(new_n329), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT67), .B1(new_n499), .B2(KEYINPUT30), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n329), .B(new_n483), .C1(new_n379), .C2(new_n380), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n340), .A2(KEYINPUT64), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n495), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n501), .B1(new_n373), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n500), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n421), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n479), .A2(new_n480), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n329), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n506), .B1(new_n381), .B2(new_n341), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n491), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT31), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n486), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n512), .A2(new_n473), .B1(new_n421), .B2(new_n504), .ZN(new_n519));
  XNOR2_X1  g333(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n490), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n515), .A2(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n512), .B2(new_n473), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n381), .A2(new_n498), .ZN(new_n525));
  AOI211_X1 g339(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n525), .C2(new_n501), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n512), .A2(new_n513), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n421), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n524), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT31), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n472), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n470), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n516), .B(new_n524), .C1(new_n528), .C2(new_n530), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n504), .A2(new_n421), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n520), .B1(new_n486), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT28), .B1(new_n512), .B2(new_n473), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n522), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n515), .A2(new_n516), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n471), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT32), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(KEYINPUT70), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n508), .A2(new_n514), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n490), .B1(new_n546), .B2(new_n486), .ZN(new_n547));
  NOR3_X1   g361(.A1(new_n537), .A2(new_n522), .A3(new_n538), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n547), .A2(KEYINPUT29), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n381), .A2(new_n341), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n509), .B1(new_n512), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n486), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT28), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n518), .A2(KEYINPUT71), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT71), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n538), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(new_n490), .A2(KEYINPUT29), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n553), .A2(new_n554), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n243), .ZN(new_n559));
  OAI21_X1  g373(.A(G472), .B1(new_n549), .B2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n534), .A2(new_n544), .A3(new_n545), .A4(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT22), .B(G137), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n198), .A2(G221), .A3(G234), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n195), .B(new_n223), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n252), .A2(G119), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n411), .A2(G128), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT24), .B(G110), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  OR2_X1    g386(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n573));
  NAND2_X1  g387(.A1(KEYINPUT72), .A2(KEYINPUT23), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n567), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(new_n574), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n576), .A2(KEYINPUT73), .A3(new_n568), .A4(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n568), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n575), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n581), .A3(G110), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT74), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n572), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n569), .A2(new_n570), .ZN(new_n587));
  OR2_X1    g401(.A1(new_n580), .A2(new_n575), .ZN(new_n588));
  XOR2_X1   g402(.A(KEYINPUT75), .B(G110), .Z(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n590), .A2(new_n224), .A3(new_n230), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n565), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n582), .A2(new_n583), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n582), .A2(new_n583), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n566), .B(new_n571), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n591), .A3(new_n564), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n294), .B1(G234), .B2(new_n243), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(G902), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT77), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n593), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT78), .Z(new_n603));
  NAND3_X1  g417(.A1(new_n593), .A2(new_n597), .A3(new_n243), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT76), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(KEYINPUT25), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n606), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n593), .A2(new_n597), .A3(new_n243), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n603), .B1(new_n598), .B2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n561), .A2(KEYINPUT79), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(KEYINPUT79), .B1(new_n561), .B2(new_n611), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n469), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT98), .B(G101), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G3));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n400), .ZN(new_n617));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n523), .A2(new_n532), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(new_n243), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n542), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n617), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n299), .A2(new_n300), .A3(new_n303), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  INV_X1    g439(.A(new_n297), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n286), .A2(new_n292), .A3(new_n295), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n296), .A2(new_n297), .A3(KEYINPUT33), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n243), .A2(G478), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n624), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n247), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n451), .A2(new_n459), .A3(new_n454), .A4(new_n468), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n623), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT34), .B(G104), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  AND3_X1   g452(.A1(new_n304), .A2(new_n308), .A3(new_n305), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n308), .B1(new_n304), .B2(new_n305), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n211), .A2(new_n227), .ZN(new_n642));
  INV_X1    g456(.A(new_n214), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n644), .B2(new_n228), .ZN(new_n645));
  INV_X1    g459(.A(G475), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n245), .A2(KEYINPUT99), .A3(G475), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n239), .A3(new_n648), .A4(new_n242), .ZN(new_n649));
  NOR4_X1   g463(.A1(new_n634), .A2(new_n639), .A3(new_n640), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n623), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NAND2_X1  g467(.A1(new_n610), .A2(new_n598), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n586), .A2(KEYINPUT100), .A3(new_n592), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n596), .B2(new_n591), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n565), .A2(KEYINPUT36), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI22_X1  g474(.A1(new_n655), .A2(new_n657), .B1(KEYINPUT36), .B2(new_n565), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n601), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n622), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n469), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT101), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G12));
  NOR3_X1   g483(.A1(new_n639), .A2(new_n640), .A3(new_n649), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT102), .B(G900), .Z(new_n671));
  AOI21_X1  g485(.A(new_n463), .B1(new_n465), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n670), .A2(KEYINPUT103), .A3(new_n461), .A4(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  INV_X1    g489(.A(new_n649), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n307), .A2(new_n309), .A3(new_n676), .A4(new_n673), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n675), .B1(new_n677), .B2(new_n460), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n561), .A2(new_n400), .A3(new_n663), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n252), .ZN(G30));
  OAI21_X1  g496(.A(new_n486), .B1(new_n528), .B2(new_n530), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n490), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n551), .A2(new_n552), .ZN(new_n685));
  AOI21_X1  g499(.A(G902), .B1(new_n685), .B2(new_n522), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n618), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n533), .B2(KEYINPUT32), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n534), .A2(new_n688), .A3(new_n544), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(KEYINPUT104), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n534), .A2(new_n688), .A3(new_n691), .A4(new_n544), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n451), .A2(new_n459), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT38), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n696), .A2(new_n453), .A3(new_n663), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n672), .B(KEYINPUT39), .Z(new_n698));
  NAND2_X1  g512(.A1(new_n400), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  INV_X1    g514(.A(new_n247), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n639), .A2(new_n640), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n697), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n694), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n200), .ZN(G45));
  NAND2_X1  g520(.A1(new_n398), .A2(new_n399), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n632), .A2(new_n247), .A3(new_n673), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n708), .A3(new_n460), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n709), .A2(new_n561), .A3(new_n663), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n223), .ZN(G48));
  INV_X1    g525(.A(new_n389), .ZN(new_n712));
  OAI21_X1  g526(.A(G469), .B1(new_n712), .B2(G902), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n399), .A3(new_n391), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n561), .A2(new_n611), .A3(new_n635), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NAND4_X1  g532(.A1(new_n561), .A2(new_n650), .A3(new_n611), .A4(new_n715), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NOR2_X1   g534(.A1(new_n714), .A2(new_n634), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n561), .A2(new_n310), .A3(new_n663), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  AND2_X1   g537(.A1(new_n554), .A2(new_n556), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n490), .B1(new_n724), .B2(new_n553), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT105), .B1(new_n725), .B2(new_n541), .ZN(new_n726));
  INV_X1    g540(.A(new_n553), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n554), .A2(new_n556), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n522), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n729), .A2(new_n730), .A3(new_n532), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n726), .A2(new_n535), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n620), .B1(new_n732), .B2(new_n471), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(new_n611), .A3(new_n702), .A4(new_n721), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  NOR3_X1   g549(.A1(new_n714), .A2(new_n708), .A3(new_n460), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n733), .A2(new_n736), .A3(new_n663), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  AOI21_X1  g552(.A(KEYINPUT106), .B1(new_n695), .B2(new_n454), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n740), .B(new_n453), .C1(new_n451), .C2(new_n459), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n707), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n708), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n561), .A3(new_n611), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n542), .B2(new_n543), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n533), .A2(KEYINPUT107), .A3(KEYINPUT32), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n542), .A2(new_n543), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n560), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n750), .A2(new_n611), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n632), .A2(KEYINPUT42), .A3(new_n247), .A4(new_n673), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n707), .A2(new_n752), .A3(new_n739), .A4(new_n741), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n744), .A2(new_n745), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n208), .ZN(G33));
  INV_X1    g569(.A(new_n677), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n742), .A2(new_n561), .A3(new_n611), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  OAI21_X1  g572(.A(new_n393), .B1(new_n395), .B2(new_n315), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n390), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n760), .B2(new_n759), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n397), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n397), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n391), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n399), .ZN(new_n768));
  INV_X1    g582(.A(new_n698), .ZN(new_n769));
  OR3_X1    g583(.A1(new_n768), .A2(KEYINPUT108), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(KEYINPUT108), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  INV_X1    g585(.A(new_n622), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n632), .A2(new_n701), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n247), .B2(KEYINPUT109), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n773), .B(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n772), .A2(new_n776), .A3(new_n664), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT44), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n739), .A2(new_n741), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n777), .B2(KEYINPUT44), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n770), .A2(new_n771), .A3(new_n778), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  INV_X1    g597(.A(new_n768), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n785), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n768), .A2(new_n787), .ZN(new_n788));
  NOR4_X1   g602(.A1(new_n780), .A2(new_n561), .A3(new_n611), .A4(new_n708), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND2_X1  g605(.A1(new_n779), .A2(new_n715), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n776), .A2(new_n464), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n751), .A3(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT117), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(KEYINPUT48), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT48), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n796), .A2(KEYINPUT117), .A3(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n733), .A2(new_n611), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n795), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n461), .A3(new_n715), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(G952), .A3(new_n198), .ZN(new_n806));
  INV_X1    g620(.A(new_n633), .ZN(new_n807));
  AND4_X1   g621(.A1(new_n463), .A2(new_n794), .A3(new_n611), .A4(new_n694), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n808), .A2(new_n807), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT116), .B1(new_n812), .B2(new_n806), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n802), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n786), .A2(new_n788), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n713), .A2(new_n391), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n399), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n779), .B(new_n804), .C1(new_n815), .C2(new_n817), .ZN(new_n818));
  AND4_X1   g632(.A1(new_n663), .A2(new_n794), .A3(new_n733), .A4(new_n795), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n632), .A2(new_n247), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n819), .B1(new_n808), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n696), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n454), .A3(new_n714), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n804), .A2(KEYINPUT50), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n803), .A2(new_n823), .A3(new_n795), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n818), .A2(new_n821), .A3(KEYINPUT51), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n824), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n831), .A2(new_n818), .A3(new_n821), .A4(new_n832), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n814), .B(new_n829), .C1(KEYINPUT51), .C2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n737), .B1(new_n679), .B2(new_n680), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n663), .A2(new_n672), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n702), .A3(new_n461), .A4(new_n400), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n690), .B2(new_n692), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n710), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT52), .B1(new_n836), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n835), .A2(new_n839), .A3(new_n842), .A4(new_n710), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n734), .A2(new_n716), .A3(new_n719), .A4(new_n722), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n754), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n306), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n633), .B1(new_n247), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n634), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n623), .A2(new_n850), .B1(new_n665), .B2(new_n469), .ZN(new_n851));
  INV_X1    g665(.A(new_n757), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n733), .A2(new_n743), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n306), .A2(new_n649), .A3(new_n672), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n561), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n742), .A2(new_n663), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n852), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n846), .A2(new_n614), .A3(new_n851), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n844), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n860), .B1(new_n844), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT54), .ZN(new_n864));
  INV_X1    g678(.A(new_n838), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n542), .A2(KEYINPUT70), .A3(new_n543), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT70), .B1(new_n542), .B2(new_n543), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n691), .B1(new_n868), .B2(new_n688), .ZN(new_n869));
  INV_X1    g683(.A(new_n692), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n865), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n710), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n842), .B1(new_n873), .B2(new_n835), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n836), .A2(new_n840), .A3(KEYINPUT52), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n754), .A2(new_n845), .A3(new_n860), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n614), .A2(new_n851), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n856), .A2(new_n857), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n757), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n878), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n858), .A2(KEYINPUT113), .A3(new_n614), .A4(new_n851), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n876), .A2(new_n877), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n862), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n864), .B1(KEYINPUT54), .B2(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n834), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n816), .B(KEYINPUT49), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n611), .A2(new_n454), .A3(new_n399), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT111), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n890), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n891), .A2(new_n701), .A3(new_n632), .A4(new_n892), .ZN(new_n893));
  AOI211_X1 g707(.A(new_n822), .B(new_n888), .C1(new_n893), .C2(KEYINPUT112), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n894), .B(new_n694), .C1(KEYINPUT112), .C2(new_n893), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n887), .A2(new_n895), .ZN(G75));
  AOI21_X1  g710(.A(new_n243), .B1(new_n862), .B2(new_n884), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n449), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n428), .A2(new_n430), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n410), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n198), .A2(G952), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G51));
  XOR2_X1   g720(.A(new_n397), .B(KEYINPUT57), .Z(new_n907));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n862), .A2(new_n908), .A3(new_n884), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n862), .B2(new_n884), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(KEYINPUT118), .B(new_n907), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n389), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n897), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n916), .A2(new_n762), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n905), .B1(new_n915), .B2(new_n917), .ZN(G54));
  AND4_X1   g732(.A1(KEYINPUT58), .A2(new_n897), .A3(G475), .A4(new_n241), .ZN(new_n919));
  NAND2_X1  g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n241), .B1(new_n897), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n919), .A2(new_n905), .A3(new_n922), .ZN(G60));
  XOR2_X1   g737(.A(new_n630), .B(KEYINPUT119), .Z(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n300), .A2(new_n243), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n886), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n924), .B(new_n927), .C1(new_n909), .C2(new_n910), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(G952), .B2(new_n198), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n928), .A2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT121), .Z(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n885), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n593), .A2(new_n597), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n905), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n934), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n862), .B2(new_n884), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n660), .A2(new_n661), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n940), .B1(new_n939), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n937), .B(KEYINPUT61), .C1(new_n943), .C2(new_n944), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(G66));
  AOI21_X1  g763(.A(new_n198), .B1(new_n467), .B2(G224), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n879), .A2(new_n845), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT123), .Z(new_n952));
  AOI21_X1  g766(.A(new_n950), .B1(new_n952), .B2(new_n198), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n900), .B1(G898), .B2(new_n198), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT124), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  NAND2_X1  g770(.A1(new_n508), .A2(new_n529), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(new_n232), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n780), .A2(new_n699), .A3(new_n849), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n612), .A2(new_n613), .ZN(new_n961));
  AOI22_X1  g775(.A1(new_n815), .A2(new_n789), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n836), .A2(new_n872), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n963), .A2(new_n705), .A3(KEYINPUT62), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT62), .B1(new_n963), .B2(new_n705), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n962), .A2(new_n782), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(G953), .ZN(new_n967));
  NAND3_X1  g781(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n959), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n963), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n782), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n754), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n790), .A2(new_n972), .A3(new_n757), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n702), .A2(new_n461), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n770), .A2(new_n751), .A3(new_n771), .A4(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n971), .A2(new_n974), .A3(KEYINPUT126), .A4(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n782), .A2(new_n977), .A3(new_n970), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n980), .B2(new_n973), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n198), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n312), .A2(G900), .A3(G953), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n969), .B1(new_n985), .B2(new_n959), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  OAI21_X1  g802(.A(new_n988), .B1(new_n982), .B2(new_n952), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n989), .A2(new_n546), .A3(new_n486), .A4(new_n522), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n966), .B2(new_n952), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n993), .B(new_n988), .C1(new_n966), .C2(new_n952), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n992), .A2(new_n490), .A3(new_n683), .A4(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(new_n988), .ZN(new_n996));
  INV_X1    g810(.A(new_n547), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n531), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n905), .B1(new_n863), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n990), .A2(new_n995), .A3(new_n999), .ZN(G57));
endmodule


