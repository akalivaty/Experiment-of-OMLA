

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n683), .B(KEYINPUT91), .ZN(n684) );
  AND2_X1 U551 ( .A1(n684), .A2(n583), .ZN(n686) );
  INV_X1 U552 ( .A(n680), .ZN(n708) );
  NAND2_X1 U553 ( .A1(n678), .A2(n791), .ZN(n680) );
  BUF_X1 U554 ( .A(n680), .Z(n723) );
  NOR2_X1 U555 ( .A1(G651), .A2(n628), .ZN(n642) );
  XNOR2_X1 U556 ( .A(G543), .B(KEYINPUT0), .ZN(n517) );
  XNOR2_X1 U557 ( .A(n517), .B(KEYINPUT67), .ZN(n628) );
  INV_X1 U558 ( .A(G651), .ZN(n523) );
  NOR2_X1 U559 ( .A1(n628), .A2(n523), .ZN(n637) );
  NAND2_X1 U560 ( .A1(n637), .A2(G77), .ZN(n518) );
  XNOR2_X1 U561 ( .A(KEYINPUT70), .B(n518), .ZN(n521) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U563 ( .A1(n636), .A2(G90), .ZN(n519) );
  XOR2_X1 U564 ( .A(KEYINPUT69), .B(n519), .Z(n520) );
  NAND2_X1 U565 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U566 ( .A(KEYINPUT9), .B(n522), .ZN(n529) );
  NOR2_X1 U567 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n524), .Z(n635) );
  NAND2_X1 U569 ( .A1(G64), .A2(n635), .ZN(n526) );
  NAND2_X1 U570 ( .A1(G52), .A2(n642), .ZN(n525) );
  NAND2_X1 U571 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U572 ( .A(KEYINPUT68), .B(n527), .Z(n528) );
  NAND2_X1 U573 ( .A1(n529), .A2(n528), .ZN(G301) );
  INV_X1 U574 ( .A(G301), .ZN(G171) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n530), .Z(n888) );
  NAND2_X1 U577 ( .A1(G137), .A2(n888), .ZN(n531) );
  XNOR2_X1 U578 ( .A(n531), .B(KEYINPUT66), .ZN(n541) );
  XOR2_X1 U579 ( .A(KEYINPUT65), .B(KEYINPUT23), .Z(n533) );
  INV_X1 U580 ( .A(G2104), .ZN(n534) );
  NOR2_X2 U581 ( .A1(G2105), .A2(n534), .ZN(n889) );
  NAND2_X1 U582 ( .A1(G101), .A2(n889), .ZN(n532) );
  XNOR2_X1 U583 ( .A(n533), .B(n532), .ZN(n539) );
  INV_X1 U584 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U585 ( .A1(n534), .A2(n535), .ZN(n896) );
  NAND2_X1 U586 ( .A1(G113), .A2(n896), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G2104), .A2(n535), .ZN(n893) );
  NAND2_X1 U588 ( .A1(G125), .A2(n893), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n543) );
  INV_X1 U592 ( .A(KEYINPUT64), .ZN(n542) );
  XNOR2_X1 U593 ( .A(n543), .B(n542), .ZN(n677) );
  BUF_X1 U594 ( .A(n677), .Z(G160) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U596 ( .A1(G135), .A2(n888), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G111), .A2(n896), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n893), .A2(G123), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT18), .B(n546), .Z(n547) );
  NOR2_X1 U601 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n889), .A2(G99), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n550), .A2(n549), .ZN(n1009) );
  XNOR2_X1 U604 ( .A(G2096), .B(n1009), .ZN(n551) );
  OR2_X1 U605 ( .A1(G2100), .A2(n551), .ZN(G156) );
  NAND2_X1 U606 ( .A1(G65), .A2(n635), .ZN(n553) );
  NAND2_X1 U607 ( .A1(G53), .A2(n642), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G91), .A2(n636), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G78), .A2(n637), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n701) );
  INV_X1 U613 ( .A(n701), .ZN(G299) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U617 ( .A(KEYINPUT76), .B(KEYINPUT7), .ZN(n569) );
  NAND2_X1 U618 ( .A1(n636), .A2(G89), .ZN(n558) );
  XNOR2_X1 U619 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U620 ( .A1(G76), .A2(n637), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U622 ( .A(KEYINPUT5), .B(n561), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n635), .A2(G63), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT75), .B(n562), .Z(n564) );
  NAND2_X1 U625 ( .A1(n642), .A2(G51), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U629 ( .A(n569), .B(n568), .ZN(G168) );
  XOR2_X1 U630 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U632 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n824) );
  NAND2_X1 U634 ( .A1(n824), .A2(G567), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n636), .A2(G81), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G68), .A2(n637), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n635), .A2(G56), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n577), .Z(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(KEYINPUT72), .ZN(n582) );
  NAND2_X1 U646 ( .A1(G43), .A2(n642), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n959) );
  INV_X1 U648 ( .A(n959), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n583), .A2(G860), .ZN(G153) );
  NAND2_X1 U650 ( .A1(G171), .A2(G868), .ZN(n593) );
  NAND2_X1 U651 ( .A1(G54), .A2(n642), .ZN(n590) );
  NAND2_X1 U652 ( .A1(G92), .A2(n636), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G66), .A2(n635), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G79), .A2(n637), .ZN(n586) );
  XNOR2_X1 U656 ( .A(KEYINPUT73), .B(n586), .ZN(n587) );
  NOR2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U659 ( .A(n591), .B(KEYINPUT15), .ZN(n954) );
  INV_X1 U660 ( .A(G868), .ZN(n656) );
  NAND2_X1 U661 ( .A1(n954), .A2(n656), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U663 ( .A(KEYINPUT74), .B(n594), .Z(G284) );
  NAND2_X1 U664 ( .A1(G868), .A2(G286), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G299), .A2(n656), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(G297) );
  INV_X1 U667 ( .A(G559), .ZN(n597) );
  NOR2_X1 U668 ( .A1(G860), .A2(n597), .ZN(n598) );
  XNOR2_X1 U669 ( .A(KEYINPUT77), .B(n598), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n954), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n959), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G868), .A2(n954), .ZN(n601) );
  NOR2_X1 U674 ( .A1(G559), .A2(n601), .ZN(n602) );
  NOR2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G559), .A2(n954), .ZN(n604) );
  XNOR2_X1 U677 ( .A(n604), .B(n959), .ZN(n652) );
  NOR2_X1 U678 ( .A1(n652), .A2(G860), .ZN(n612) );
  NAND2_X1 U679 ( .A1(G55), .A2(n642), .ZN(n605) );
  XNOR2_X1 U680 ( .A(n605), .B(KEYINPUT78), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n636), .A2(G93), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G80), .A2(n637), .ZN(n609) );
  NAND2_X1 U684 ( .A1(G67), .A2(n635), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n655) );
  XOR2_X1 U687 ( .A(n612), .B(n655), .Z(G145) );
  NAND2_X1 U688 ( .A1(G88), .A2(n636), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G75), .A2(n637), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G62), .A2(n635), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G50), .A2(n642), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n618), .A2(n617), .ZN(G166) );
  NAND2_X1 U695 ( .A1(G86), .A2(n636), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G61), .A2(n635), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n625) );
  XOR2_X1 U698 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n622) );
  NAND2_X1 U699 ( .A1(G73), .A2(n637), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n622), .B(n621), .ZN(n623) );
  XOR2_X1 U701 ( .A(KEYINPUT80), .B(n623), .Z(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n642), .A2(G48), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(G305) );
  NAND2_X1 U705 ( .A1(G87), .A2(n628), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U708 ( .A1(n635), .A2(n631), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G49), .A2(n642), .ZN(n632) );
  XOR2_X1 U710 ( .A(KEYINPUT79), .B(n632), .Z(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(G288) );
  AND2_X1 U712 ( .A1(n635), .A2(G60), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G85), .A2(n636), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G72), .A2(n637), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n642), .A2(G47), .ZN(n643) );
  NAND2_X1 U718 ( .A1(n644), .A2(n643), .ZN(G290) );
  XOR2_X1 U719 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n646) );
  XNOR2_X1 U720 ( .A(G166), .B(KEYINPUT19), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n649) );
  XOR2_X1 U722 ( .A(n655), .B(G305), .Z(n647) );
  XNOR2_X1 U723 ( .A(n647), .B(G288), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n649), .B(n648), .ZN(n651) );
  XNOR2_X1 U725 ( .A(G290), .B(n701), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(n910) );
  XNOR2_X1 U727 ( .A(n910), .B(n652), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n653), .A2(G868), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(KEYINPUT84), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(G295) );
  NAND2_X1 U732 ( .A1(G2084), .A2(G2078), .ZN(n659) );
  XOR2_X1 U733 ( .A(KEYINPUT20), .B(n659), .Z(n660) );
  NAND2_X1 U734 ( .A1(G2090), .A2(n660), .ZN(n661) );
  XNOR2_X1 U735 ( .A(KEYINPUT21), .B(n661), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n662), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U738 ( .A1(G220), .A2(G219), .ZN(n663) );
  XOR2_X1 U739 ( .A(KEYINPUT22), .B(n663), .Z(n664) );
  NOR2_X1 U740 ( .A1(G218), .A2(n664), .ZN(n665) );
  NAND2_X1 U741 ( .A1(G96), .A2(n665), .ZN(n828) );
  NAND2_X1 U742 ( .A1(n828), .A2(G2106), .ZN(n669) );
  NAND2_X1 U743 ( .A1(G69), .A2(G120), .ZN(n666) );
  NOR2_X1 U744 ( .A1(G237), .A2(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(G108), .A2(n667), .ZN(n829) );
  NAND2_X1 U746 ( .A1(n829), .A2(G567), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n669), .A2(n668), .ZN(n844) );
  NAND2_X1 U748 ( .A1(G483), .A2(G661), .ZN(n670) );
  NOR2_X1 U749 ( .A1(n844), .A2(n670), .ZN(n827) );
  NAND2_X1 U750 ( .A1(n827), .A2(G36), .ZN(G176) );
  NAND2_X1 U751 ( .A1(G138), .A2(n888), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G102), .A2(n889), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n676) );
  NAND2_X1 U754 ( .A1(G114), .A2(n896), .ZN(n674) );
  NAND2_X1 U755 ( .A1(G126), .A2(n893), .ZN(n673) );
  NAND2_X1 U756 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U757 ( .A1(n676), .A2(n675), .ZN(G164) );
  INV_X1 U758 ( .A(G166), .ZN(G303) );
  NAND2_X1 U759 ( .A1(G40), .A2(n677), .ZN(n790) );
  INV_X1 U760 ( .A(n790), .ZN(n678) );
  NOR2_X1 U761 ( .A1(G164), .A2(G1384), .ZN(n791) );
  NAND2_X1 U762 ( .A1(G1996), .A2(n708), .ZN(n679) );
  XNOR2_X1 U763 ( .A(n679), .B(KEYINPUT26), .ZN(n682) );
  NAND2_X1 U764 ( .A1(G1341), .A2(n723), .ZN(n681) );
  NAND2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U766 ( .A1(n686), .A2(n954), .ZN(n685) );
  XNOR2_X1 U767 ( .A(n685), .B(KEYINPUT93), .ZN(n698) );
  NAND2_X1 U768 ( .A1(n686), .A2(n954), .ZN(n691) );
  NAND2_X1 U769 ( .A1(G1348), .A2(n723), .ZN(n688) );
  NAND2_X1 U770 ( .A1(G2067), .A2(n708), .ZN(n687) );
  NAND2_X1 U771 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U772 ( .A(KEYINPUT92), .B(n689), .ZN(n690) );
  NAND2_X1 U773 ( .A1(n691), .A2(n690), .ZN(n696) );
  NAND2_X1 U774 ( .A1(n708), .A2(G2072), .ZN(n692) );
  XNOR2_X1 U775 ( .A(n692), .B(KEYINPUT27), .ZN(n694) );
  INV_X1 U776 ( .A(G1956), .ZN(n972) );
  NOR2_X1 U777 ( .A1(n972), .A2(n708), .ZN(n693) );
  NOR2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n700) );
  NOR2_X1 U779 ( .A1(n701), .A2(n700), .ZN(n695) );
  XOR2_X1 U780 ( .A(n695), .B(KEYINPUT28), .Z(n699) );
  AND2_X1 U781 ( .A1(n696), .A2(n699), .ZN(n697) );
  NAND2_X1 U782 ( .A1(n698), .A2(n697), .ZN(n705) );
  INV_X1 U783 ( .A(n699), .ZN(n703) );
  NAND2_X1 U784 ( .A1(n701), .A2(n700), .ZN(n702) );
  OR2_X1 U785 ( .A1(n703), .A2(n702), .ZN(n704) );
  AND2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n707) );
  XOR2_X1 U787 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n706) );
  XNOR2_X1 U788 ( .A(n707), .B(n706), .ZN(n713) );
  INV_X1 U789 ( .A(G1961), .ZN(n983) );
  NAND2_X1 U790 ( .A1(n723), .A2(n983), .ZN(n710) );
  XNOR2_X1 U791 ( .A(G2078), .B(KEYINPUT25), .ZN(n928) );
  NAND2_X1 U792 ( .A1(n708), .A2(n928), .ZN(n709) );
  NAND2_X1 U793 ( .A1(n710), .A2(n709), .ZN(n714) );
  AND2_X1 U794 ( .A1(n714), .A2(G171), .ZN(n711) );
  XOR2_X1 U795 ( .A(KEYINPUT90), .B(n711), .Z(n712) );
  NAND2_X1 U796 ( .A1(n713), .A2(n712), .ZN(n736) );
  NOR2_X1 U797 ( .A1(G171), .A2(n714), .ZN(n719) );
  NAND2_X1 U798 ( .A1(G8), .A2(n723), .ZN(n765) );
  NOR2_X1 U799 ( .A1(G1966), .A2(n765), .ZN(n738) );
  NOR2_X1 U800 ( .A1(G2084), .A2(n723), .ZN(n737) );
  NOR2_X1 U801 ( .A1(n738), .A2(n737), .ZN(n715) );
  NAND2_X1 U802 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U803 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U804 ( .A1(n717), .A2(G168), .ZN(n718) );
  NOR2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n722) );
  XNOR2_X1 U806 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n720) );
  XNOR2_X1 U807 ( .A(n720), .B(KEYINPUT31), .ZN(n721) );
  XNOR2_X1 U808 ( .A(n722), .B(n721), .ZN(n735) );
  NOR2_X1 U809 ( .A1(G1971), .A2(n765), .ZN(n725) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n723), .ZN(n724) );
  NOR2_X1 U811 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U812 ( .A(KEYINPUT97), .B(n726), .Z(n727) );
  NAND2_X1 U813 ( .A1(n727), .A2(G303), .ZN(n729) );
  AND2_X1 U814 ( .A1(n735), .A2(n729), .ZN(n728) );
  NAND2_X1 U815 ( .A1(n736), .A2(n728), .ZN(n733) );
  INV_X1 U816 ( .A(n729), .ZN(n730) );
  OR2_X1 U817 ( .A1(n730), .A2(G286), .ZN(n731) );
  AND2_X1 U818 ( .A1(G8), .A2(n731), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U820 ( .A(n734), .B(KEYINPUT32), .ZN(n759) );
  NAND2_X1 U821 ( .A1(n736), .A2(n735), .ZN(n741) );
  AND2_X1 U822 ( .A1(G8), .A2(n737), .ZN(n739) );
  NOR2_X1 U823 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U824 ( .A1(n741), .A2(n740), .ZN(n757) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n952) );
  INV_X1 U826 ( .A(n952), .ZN(n742) );
  OR2_X1 U827 ( .A1(n742), .A2(n765), .ZN(n746) );
  INV_X1 U828 ( .A(n746), .ZN(n743) );
  AND2_X1 U829 ( .A1(n757), .A2(n743), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n759), .A2(n744), .ZN(n750) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n751) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n745) );
  NOR2_X1 U833 ( .A1(n751), .A2(n745), .ZN(n948) );
  OR2_X1 U834 ( .A1(n746), .A2(n948), .ZN(n748) );
  INV_X1 U835 ( .A(KEYINPUT33), .ZN(n747) );
  AND2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n756) );
  NAND2_X1 U838 ( .A1(n751), .A2(KEYINPUT33), .ZN(n752) );
  NOR2_X1 U839 ( .A1(n765), .A2(n752), .ZN(n754) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n942) );
  INV_X1 U841 ( .A(n942), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n755) );
  AND2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n771) );
  AND2_X1 U844 ( .A1(n757), .A2(n765), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n759), .A2(n758), .ZN(n769) );
  INV_X1 U846 ( .A(n765), .ZN(n762) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G8), .A2(n760), .ZN(n761) );
  NOR2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n767) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U851 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U856 ( .A(n772), .B(KEYINPUT98), .ZN(n793) );
  NAND2_X1 U857 ( .A1(G105), .A2(n889), .ZN(n773) );
  XNOR2_X1 U858 ( .A(n773), .B(KEYINPUT38), .ZN(n780) );
  NAND2_X1 U859 ( .A1(G141), .A2(n888), .ZN(n775) );
  NAND2_X1 U860 ( .A1(G117), .A2(n896), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U862 ( .A1(n893), .A2(G129), .ZN(n776) );
  XOR2_X1 U863 ( .A(KEYINPUT88), .B(n776), .Z(n777) );
  NOR2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n876) );
  NAND2_X1 U866 ( .A1(G1996), .A2(n876), .ZN(n789) );
  NAND2_X1 U867 ( .A1(G95), .A2(n889), .ZN(n782) );
  NAND2_X1 U868 ( .A1(G119), .A2(n893), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U870 ( .A1(G131), .A2(n888), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G107), .A2(n896), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U874 ( .A(n787), .B(KEYINPUT87), .ZN(n903) );
  NAND2_X1 U875 ( .A1(G1991), .A2(n903), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n789), .A2(n788), .ZN(n1007) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n819) );
  NAND2_X1 U878 ( .A1(n1007), .A2(n819), .ZN(n792) );
  XNOR2_X1 U879 ( .A(n792), .B(KEYINPUT89), .ZN(n811) );
  NOR2_X1 U880 ( .A1(n793), .A2(n811), .ZN(n805) );
  XNOR2_X1 U881 ( .A(KEYINPUT37), .B(G2067), .ZN(n817) );
  NAND2_X1 U882 ( .A1(n896), .A2(G116), .ZN(n794) );
  XOR2_X1 U883 ( .A(KEYINPUT85), .B(n794), .Z(n796) );
  NAND2_X1 U884 ( .A1(n893), .A2(G128), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U886 ( .A(n797), .B(KEYINPUT35), .ZN(n802) );
  NAND2_X1 U887 ( .A1(G140), .A2(n888), .ZN(n799) );
  NAND2_X1 U888 ( .A1(G104), .A2(n889), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U890 ( .A(KEYINPUT34), .B(n800), .Z(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XOR2_X1 U892 ( .A(n803), .B(KEYINPUT36), .Z(n906) );
  OR2_X1 U893 ( .A1(n817), .A2(n906), .ZN(n804) );
  XOR2_X1 U894 ( .A(KEYINPUT86), .B(n804), .Z(n1016) );
  NAND2_X1 U895 ( .A1(n819), .A2(n1016), .ZN(n815) );
  NAND2_X1 U896 ( .A1(n805), .A2(n815), .ZN(n806) );
  XNOR2_X1 U897 ( .A(n806), .B(KEYINPUT99), .ZN(n808) );
  XNOR2_X1 U898 ( .A(G1986), .B(G290), .ZN(n950) );
  NAND2_X1 U899 ( .A1(n950), .A2(n819), .ZN(n807) );
  NAND2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n822) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n903), .ZN(n1008) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n1008), .A2(n809), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U905 ( .A1(G1996), .A2(n876), .ZN(n1004) );
  NOR2_X1 U906 ( .A1(n812), .A2(n1004), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n813), .B(KEYINPUT39), .ZN(n814) );
  XNOR2_X1 U908 ( .A(n814), .B(KEYINPUT100), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n816), .A2(n815), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n817), .A2(n906), .ZN(n1021) );
  NAND2_X1 U911 ( .A1(n818), .A2(n1021), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U914 ( .A(KEYINPUT40), .B(n823), .ZN(G329) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n824), .ZN(G217) );
  AND2_X1 U916 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U917 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U918 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U921 ( .A(G120), .ZN(G236) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  INV_X1 U923 ( .A(G69), .ZN(G235) );
  NOR2_X1 U924 ( .A1(n829), .A2(n828), .ZN(G325) );
  INV_X1 U925 ( .A(G325), .ZN(G261) );
  XOR2_X1 U926 ( .A(KEYINPUT101), .B(G2435), .Z(n831) );
  XNOR2_X1 U927 ( .A(G1341), .B(G1348), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n831), .B(n830), .ZN(n841) );
  XOR2_X1 U929 ( .A(G2446), .B(KEYINPUT104), .Z(n833) );
  XNOR2_X1 U930 ( .A(G2430), .B(G2438), .ZN(n832) );
  XNOR2_X1 U931 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U932 ( .A(KEYINPUT103), .B(KEYINPUT102), .Z(n835) );
  XNOR2_X1 U933 ( .A(G2427), .B(G2454), .ZN(n834) );
  XNOR2_X1 U934 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U935 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2443), .B(G2451), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(n842) );
  NAND2_X1 U939 ( .A1(n842), .A2(G14), .ZN(n843) );
  XNOR2_X1 U940 ( .A(n843), .B(KEYINPUT105), .ZN(n918) );
  XNOR2_X1 U941 ( .A(n918), .B(KEYINPUT106), .ZN(G401) );
  INV_X1 U942 ( .A(n844), .ZN(G319) );
  XOR2_X1 U943 ( .A(G1976), .B(G1971), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n856) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G2474), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1966), .B(KEYINPUT108), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(G1981), .B(G1956), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1961), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U956 ( .A(G2678), .B(G2072), .Z(n858) );
  XNOR2_X1 U957 ( .A(G2084), .B(G2078), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U959 ( .A(n859), .B(G2100), .Z(n861) );
  XNOR2_X1 U960 ( .A(G2067), .B(G2090), .ZN(n860) );
  XNOR2_X1 U961 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U962 ( .A(G2096), .B(KEYINPUT107), .Z(n863) );
  XNOR2_X1 U963 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U965 ( .A(n865), .B(n864), .Z(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n893), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n896), .A2(G112), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G136), .A2(n888), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G100), .A2(n889), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(G162) );
  XOR2_X1 U974 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U977 ( .A(G164), .B(G162), .Z(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n902) );
  NAND2_X1 U980 ( .A1(n896), .A2(G115), .ZN(n879) );
  XOR2_X1 U981 ( .A(KEYINPUT113), .B(n879), .Z(n881) );
  NAND2_X1 U982 ( .A1(n893), .A2(G127), .ZN(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U984 ( .A(KEYINPUT47), .B(n882), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G139), .A2(n888), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G103), .A2(n889), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U988 ( .A(KEYINPUT112), .B(n885), .Z(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n997) );
  NAND2_X1 U990 ( .A1(G142), .A2(n888), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G106), .A2(n889), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n892), .B(KEYINPUT45), .ZN(n895) );
  NAND2_X1 U994 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G118), .A2(n896), .ZN(n897) );
  XNOR2_X1 U997 ( .A(KEYINPUT111), .B(n897), .ZN(n898) );
  NOR2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n997), .B(n900), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n908) );
  XOR2_X1 U1001 ( .A(G160), .B(n903), .Z(n904) );
  XNOR2_X1 U1002 ( .A(n1009), .B(n904), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(G286), .B(n910), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(G171), .B(n954), .ZN(n911) );
  XNOR2_X1 U1008 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1009 ( .A(n913), .B(n959), .Z(n914) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G229), .A2(G227), .ZN(n915) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n916), .ZN(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1019 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n1024) );
  XNOR2_X1 U1020 ( .A(G1996), .B(G32), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(G33), .B(G2072), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n927) );
  XOR2_X1 U1023 ( .A(G2067), .B(G26), .Z(n923) );
  NAND2_X1 U1024 ( .A1(n923), .A2(G28), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(G25), .B(G1991), .ZN(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1028 ( .A(G27), .B(n928), .Z(n929) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1030 ( .A(KEYINPUT53), .B(n931), .Z(n935) );
  XNOR2_X1 U1031 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(n932), .B(G34), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G2084), .B(n933), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(G35), .B(G2090), .ZN(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(n1024), .B(n938), .ZN(n939) );
  NOR2_X1 U1038 ( .A1(G29), .A2(n939), .ZN(n940) );
  XOR2_X1 U1039 ( .A(KEYINPUT124), .B(n940), .Z(n941) );
  NAND2_X1 U1040 ( .A1(G11), .A2(n941), .ZN(n995) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .ZN(n965) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G168), .ZN(n943) );
  NAND2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1044 ( .A(KEYINPUT57), .B(n944), .ZN(n963) );
  XNOR2_X1 U1045 ( .A(G299), .B(G1956), .ZN(n946) );
  AND2_X1 U1046 ( .A1(G1971), .A2(G303), .ZN(n945) );
  NOR2_X1 U1047 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(n953), .B(KEYINPUT125), .ZN(n958) );
  XOR2_X1 U1052 ( .A(n954), .B(G1348), .Z(n956) );
  XOR2_X1 U1053 ( .A(G171), .B(G1961), .Z(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G1341), .B(n959), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n993) );
  INV_X1 U1060 ( .A(G16), .ZN(n991) );
  XOR2_X1 U1061 ( .A(G1986), .B(G24), .Z(n969) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G22), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(G23), .B(G1976), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n971) );
  XNOR2_X1 U1066 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(n971), .B(n970), .ZN(n988) );
  XOR2_X1 U1068 ( .A(G1966), .B(G21), .Z(n982) );
  XNOR2_X1 U1069 ( .A(G20), .B(n972), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G1341), .B(G19), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G6), .ZN(n973) );
  NOR2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n979) );
  XOR2_X1 U1074 ( .A(KEYINPUT59), .B(G1348), .Z(n977) );
  XNOR2_X1 U1075 ( .A(G4), .B(n977), .ZN(n978) );
  NOR2_X1 U1076 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(KEYINPUT60), .B(n980), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n986) );
  XOR2_X1 U1079 ( .A(KEYINPUT126), .B(n983), .Z(n984) );
  XNOR2_X1 U1080 ( .A(G5), .B(n984), .ZN(n985) );
  NOR2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1083 ( .A(KEYINPUT61), .B(n989), .Z(n990) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n1028) );
  XOR2_X1 U1087 ( .A(G2072), .B(KEYINPUT118), .Z(n996) );
  XNOR2_X1 U1088 ( .A(n997), .B(n996), .ZN(n1000) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n998) );
  XNOR2_X1 U1090 ( .A(KEYINPUT119), .B(n998), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(KEYINPUT50), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT120), .B(n1002), .ZN(n1019) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT51), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(KEYINPUT116), .B(n1006), .ZN(n1014) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(G2084), .B(G160), .Z(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(KEYINPUT117), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT121), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(n1023), .B(KEYINPUT52), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(G29), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

