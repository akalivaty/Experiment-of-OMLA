//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:59 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT65), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(KEYINPUT65), .B1(G567), .B2(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G125), .ZN(new_n463));
  OR2_X1    g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G2105), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n465), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n470), .A2(new_n472), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT66), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n470), .A2(new_n482), .A3(new_n471), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n480), .A2(new_n471), .ZN(new_n486));
  NOR2_X1   g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT67), .ZN(new_n488));
  INV_X1    g063(.A(G112), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n473), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(G124), .A2(new_n486), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n485), .A2(new_n491), .ZN(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n478), .B2(new_n479), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n470), .A2(new_n497), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  OAI211_X1 g076(.A(new_n501), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n502));
  NAND2_X1  g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n502), .B(KEYINPUT68), .C1(new_n480), .C2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n464), .B2(new_n465), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n471), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n499), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT69), .B1(new_n514), .B2(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT6), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(new_n518), .B1(new_n514), .B2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n522), .B2(KEYINPUT70), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(KEYINPUT5), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n513), .A2(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n526), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n517), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n529), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(KEYINPUT7), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n526), .A2(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G89), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n538), .B1(new_n527), .B2(new_n539), .C1(new_n540), .C2(new_n520), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G168));
  NAND2_X1  g120(.A1(G77), .A2(G543), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n523), .A2(new_n525), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G651), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G52), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n552), .A2(new_n520), .B1(new_n527), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  AND2_X1   g130(.A1(new_n526), .A2(G56), .ZN(new_n556));
  AND2_X1   g131(.A1(G68), .A2(G543), .ZN(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  INV_X1    g136(.A(new_n527), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n515), .A2(new_n518), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n514), .A2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n522), .ZN(new_n566));
  AOI22_X1  g141(.A1(G81), .A2(new_n562), .B1(new_n566), .B2(G43), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n560), .A2(G860), .A3(new_n561), .A4(new_n567), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT73), .Z(G188));
  NAND3_X1  g148(.A1(new_n519), .A2(G91), .A3(new_n526), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT74), .ZN(new_n575));
  NAND2_X1  g150(.A1(G53), .A2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT9), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n519), .A2(new_n578), .A3(G53), .A4(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n547), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n577), .A2(new_n579), .B1(new_n582), .B2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n575), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND2_X1  g161(.A1(new_n562), .A2(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n566), .A2(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n523), .B2(new_n525), .ZN(new_n592));
  AND2_X1   g167(.A1(G73), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n519), .A2(G86), .A3(new_n526), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n519), .A2(KEYINPUT76), .A3(G86), .A4(new_n526), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n519), .A2(G48), .A3(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n594), .B2(KEYINPUT75), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(G72), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G60), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n547), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT77), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(KEYINPUT77), .B(new_n605), .C1(new_n547), .C2(new_n606), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(G651), .A3(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  AOI22_X1  g189(.A1(G85), .A2(new_n562), .B1(new_n566), .B2(G47), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(G290));
  NAND2_X1  g191(.A1(G301), .A2(G868), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n526), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(new_n517), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n566), .A2(G54), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n621));
  INV_X1    g196(.A(G92), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n527), .B2(new_n622), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n619), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n527), .A2(new_n622), .A3(new_n621), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n617), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n617), .B1(new_n626), .B2(G868), .ZN(G321));
  NOR2_X1   g203(.A1(G299), .A2(G868), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(G168), .B2(G868), .ZN(G297));
  AOI21_X1  g205(.A(new_n629), .B1(G168), .B2(G868), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND3_X1  g208(.A1(new_n560), .A2(new_n561), .A3(new_n567), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n624), .A2(new_n625), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n636), .A2(G559), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT80), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n635), .B1(new_n638), .B2(G868), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n486), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n471), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(G135), .B2(new_n484), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT81), .Z(new_n646));
  INV_X1    g221(.A(G2096), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n470), .A2(new_n474), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT12), .Z(new_n650));
  XOR2_X1   g225(.A(KEYINPUT13), .B(G2100), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT82), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT83), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT85), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT17), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT86), .B(G2100), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2072), .B(G2078), .Z(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n677), .B2(KEYINPUT18), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(new_n647), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n687), .A2(new_n688), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n689), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(KEYINPUT87), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n692), .A2(new_n693), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT20), .Z(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G1981), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT88), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n705), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n703), .B(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n707), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n708), .A2(new_n712), .ZN(G229));
  XNOR2_X1  g288(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G34), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(new_n716), .B2(new_n476), .ZN(new_n718));
  INV_X1    g293(.A(G2084), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(G33), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT25), .Z(new_n724));
  AOI22_X1  g299(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n471), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G139), .B2(new_n484), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n722), .B1(new_n727), .B2(new_n716), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(G2072), .Z(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G35), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G162), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT29), .B(G2090), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G16), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G5), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G171), .B2(new_n735), .ZN(new_n737));
  AOI211_X1 g312(.A(new_n721), .B(new_n734), .C1(G1961), .C2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  NOR2_X1   g314(.A1(G164), .A2(new_n716), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G27), .B2(new_n716), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n716), .A2(G26), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n484), .A2(G140), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n745));
  INV_X1    g320(.A(G116), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G2105), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n486), .B2(G128), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n743), .B1(new_n750), .B2(new_n716), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n739), .A2(new_n741), .B1(new_n751), .B2(G2067), .ZN(new_n752));
  OAI221_X1 g327(.A(new_n752), .B1(G2067), .B2(new_n751), .C1(new_n716), .C2(new_n646), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT94), .B(G28), .Z(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(KEYINPUT30), .B2(new_n754), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n718), .B2(new_n719), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n759), .B1(new_n737), .B2(G1961), .C1(new_n741), .C2(new_n739), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n753), .A2(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G19), .B(new_n634), .S(G16), .Z(new_n762));
  INV_X1    g337(.A(G1341), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n474), .A2(G105), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT26), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n765), .B(new_n767), .C1(G129), .C2(new_n486), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n484), .A2(G141), .ZN(new_n769));
  AND3_X1   g344(.A1(new_n768), .A2(new_n769), .A3(KEYINPUT92), .ZN(new_n770));
  AOI21_X1  g345(.A(KEYINPUT92), .B1(new_n768), .B2(new_n769), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(KEYINPUT93), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G29), .B2(G32), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n774), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT27), .B(G1996), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n738), .A2(new_n761), .A3(new_n764), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n735), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n735), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n626), .B2(new_n735), .ZN(new_n786));
  INV_X1    g361(.A(G1348), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n784), .B(new_n788), .C1(new_n777), .C2(new_n778), .ZN(new_n789));
  NOR2_X1   g364(.A1(G16), .A2(G21), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G168), .B2(G16), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1966), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n780), .A2(new_n789), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n735), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G166), .B2(new_n735), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G6), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n603), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT32), .B(G1981), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n799), .A2(new_n800), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n735), .A2(G23), .ZN(new_n803));
  INV_X1    g378(.A(G288), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n735), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n797), .A2(new_n801), .A3(new_n802), .A4(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  MUX2_X1   g385(.A(G24), .B(G290), .S(G16), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G1986), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(G1986), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n716), .A2(G25), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n484), .A2(G131), .ZN(new_n815));
  OAI21_X1  g390(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n816));
  INV_X1    g391(.A(G107), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(G2105), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(new_n486), .B2(G119), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n814), .B1(new_n821), .B2(new_n716), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  NOR3_X1   g399(.A1(new_n813), .A2(KEYINPUT89), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n809), .A2(new_n810), .A3(new_n812), .A4(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n793), .A2(new_n828), .A3(new_n829), .ZN(G150));
  INV_X1    g405(.A(G150), .ZN(G311));
  NOR2_X1   g406(.A1(new_n636), .A2(new_n632), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT38), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n547), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n517), .B1(new_n836), .B2(KEYINPUT95), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(KEYINPUT95), .B2(new_n836), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT97), .B(G93), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT96), .B(G55), .ZN(new_n840));
  AOI22_X1  g415(.A1(new_n562), .A2(new_n839), .B1(new_n566), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n634), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n634), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n833), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT98), .B(G860), .Z(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n849), .B1(new_n838), .B2(new_n841), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  XNOR2_X1  g428(.A(new_n646), .B(G160), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n820), .B(KEYINPUT99), .ZN(new_n856));
  INV_X1    g431(.A(new_n650), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  INV_X1    g434(.A(G118), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n860), .B2(G2105), .ZN(new_n861));
  AND2_X1   g436(.A1(new_n484), .A2(G142), .ZN(new_n862));
  AOI211_X1 g437(.A(new_n861), .B(new_n862), .C1(G130), .C2(new_n486), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n858), .B(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n727), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n506), .A2(new_n509), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n499), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n772), .A2(new_n750), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n772), .A2(new_n750), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n870), .A2(new_n871), .A3(new_n868), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n865), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n727), .A3(new_n872), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n864), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n864), .B1(new_n875), .B2(new_n877), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n855), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(KEYINPUT100), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(new_n855), .C1(new_n879), .C2(new_n880), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n875), .A2(new_n877), .ZN(new_n886));
  INV_X1    g461(.A(new_n864), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n855), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT101), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n864), .A2(new_n875), .A3(new_n877), .A4(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n878), .A2(KEYINPUT101), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n885), .A2(KEYINPUT40), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT40), .B1(new_n885), .B2(new_n894), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(G395));
  INV_X1    g472(.A(G868), .ZN(new_n898));
  XNOR2_X1  g473(.A(G290), .B(G305), .ZN(new_n899));
  XNOR2_X1  g474(.A(G303), .B(G288), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n899), .B(new_n900), .Z(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT42), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n899), .B(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n626), .A2(G299), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n636), .A2(new_n575), .A3(new_n583), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n912));
  MUX2_X1   g487(.A(new_n911), .B(new_n909), .S(KEYINPUT102), .Z(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n913), .B2(KEYINPUT41), .ZN(new_n914));
  INV_X1    g489(.A(new_n845), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n638), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n638), .B(new_n845), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n918), .A2(new_n913), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n908), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n903), .B(new_n907), .C1(new_n917), .C2(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n898), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n842), .A2(new_n898), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  OR3_X1    g500(.A1(new_n923), .A2(KEYINPUT104), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT104), .B1(new_n923), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(G295));
  OR2_X1    g503(.A1(new_n923), .A2(new_n925), .ZN(G331));
  XNOR2_X1  g504(.A(G168), .B(G301), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(new_n845), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT41), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n911), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n934), .B(new_n901), .C1(new_n913), .C2(new_n933), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n930), .B(new_n915), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n914), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n931), .A2(new_n913), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n904), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n935), .A2(KEYINPUT43), .A3(new_n936), .A4(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n936), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n904), .B1(new_n938), .B2(new_n939), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT44), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n935), .A2(new_n942), .A3(new_n936), .A4(new_n940), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n943), .B2(new_n944), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(new_n952), .ZN(G397));
  OAI21_X1  g528(.A(new_n472), .B1(new_n479), .B2(new_n478), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n474), .A2(G101), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n954), .A2(G40), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(G125), .B1(new_n478), .B2(new_n479), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n471), .B1(new_n957), .B2(new_n467), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT105), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n469), .A2(new_n960), .A3(G40), .A4(new_n475), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1384), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n867), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR4_X1   g541(.A1(G290), .A2(G1986), .A3(new_n962), .A4(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT127), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(KEYINPUT48), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(KEYINPUT48), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n772), .B(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n749), .B(G2067), .Z(new_n974));
  NAND2_X1  g549(.A1(new_n821), .A2(new_n823), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n821), .A2(new_n823), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n966), .A2(new_n962), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n969), .A2(new_n970), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT46), .B1(new_n978), .B2(new_n971), .ZN(new_n981));
  XOR2_X1   g556(.A(new_n981), .B(KEYINPUT125), .Z(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(KEYINPUT46), .A3(new_n971), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT126), .Z(new_n984));
  INV_X1    g559(.A(new_n974), .ZN(new_n985));
  INV_X1    g560(.A(new_n772), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n982), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n972), .A2(new_n985), .A3(new_n975), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n749), .A2(G2067), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n978), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n980), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT123), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  NOR2_X1   g571(.A1(G168), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1966), .ZN(new_n999));
  AOI21_X1  g574(.A(G1384), .B1(new_n499), .B2(new_n866), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n959), .B(new_n961), .C1(new_n1000), .C2(KEYINPUT45), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n1002));
  OAI211_X1 g577(.A(KEYINPUT110), .B(new_n999), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n511), .A2(new_n963), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1005));
  AOI211_X1 g580(.A(KEYINPUT50), .B(G1384), .C1(new_n499), .C2(new_n866), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n959), .A2(new_n961), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n719), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n511), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n966), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(KEYINPUT110), .B1(new_n1012), .B2(new_n999), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT119), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n1009), .A4(new_n1003), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n998), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(G168), .A3(new_n1019), .ZN(new_n1021));
  AND2_X1   g596(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n997), .A2(KEYINPUT51), .ZN(new_n1024));
  OAI21_X1  g599(.A(G8), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1020), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT62), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n995), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n739), .A2(KEYINPUT53), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n966), .A2(new_n1008), .A3(new_n1011), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n511), .B2(new_n963), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1033), .A2(new_n1006), .A3(new_n962), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT120), .B(G1961), .Z(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n511), .B2(new_n963), .ZN(new_n1037));
  AOI211_X1 g612(.A(new_n965), .B(G1384), .C1(new_n499), .C2(new_n866), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n962), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n1039), .B2(new_n739), .ZN(new_n1040));
  OAI21_X1  g615(.A(G171), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT121), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1035), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n867), .A2(KEYINPUT45), .A3(new_n963), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1046), .A2(new_n959), .A3(new_n961), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1047), .A2(G2078), .A3(new_n1037), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1045), .B(new_n1031), .C1(new_n1048), .C2(KEYINPUT53), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1050), .A3(G171), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n529), .B2(new_n531), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n796), .B1(new_n1047), .B2(new_n1037), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n964), .A2(KEYINPUT50), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(new_n1008), .C1(KEYINPUT50), .C2(new_n1004), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1058), .B2(G2090), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1059), .B2(G8), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT106), .ZN(new_n1061));
  INV_X1    g636(.A(G2090), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1056), .A2(new_n1061), .B1(new_n1062), .B2(new_n1034), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT106), .B(new_n796), .C1(new_n1047), .C2(new_n1037), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n996), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1060), .B1(new_n1065), .B2(new_n1055), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G288), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT108), .B(G1976), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT52), .B1(G288), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1000), .A2(new_n959), .A3(new_n961), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1072), .A2(KEYINPUT107), .A3(G8), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT107), .B1(new_n1072), .B2(G8), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1069), .B(new_n1071), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(G8), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT107), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1072), .A2(KEYINPUT107), .A3(G8), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1068), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n594), .A2(new_n601), .A3(new_n596), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(G1981), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT109), .B1(new_n603), .B2(new_n701), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT109), .ZN(new_n1087));
  NOR4_X1   g662(.A1(new_n600), .A2(new_n1087), .A3(new_n602), .A4(G1981), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT49), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1083), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT49), .B(new_n1085), .C1(new_n1086), .C2(new_n1088), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1082), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1052), .A2(new_n1066), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1021), .A2(new_n1022), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT123), .B(KEYINPUT62), .C1(new_n1096), .C2(new_n1020), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1029), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1065), .A2(new_n1055), .ZN(new_n1099));
  OAI211_X1 g674(.A(G8), .B(G168), .C1(new_n1010), .C2(new_n1013), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1034), .A2(new_n1062), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1064), .A3(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1104), .A2(G8), .A3(new_n1055), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1101), .A2(new_n1093), .A3(KEYINPUT63), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT111), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1083), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1092), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1060), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1082), .ZN(new_n1112));
  AND4_X1   g687(.A1(new_n1110), .A2(new_n1111), .A3(new_n1105), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1100), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1107), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1066), .A2(new_n1093), .A3(new_n1107), .A4(new_n1114), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1106), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT112), .B(G1956), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n959), .B(new_n961), .C1(new_n1000), .C2(new_n1032), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1038), .A2(new_n962), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1037), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1129));
  OR2_X1    g704(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1128), .A2(KEYINPUT113), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1130), .A2(new_n1123), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT113), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1130), .A2(new_n1129), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1072), .A2(G2067), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1043), .B2(new_n787), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n636), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT61), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1143), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n636), .A2(KEYINPUT60), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1144), .A2(new_n1132), .B1(new_n1140), .B2(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1140), .A2(new_n636), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1140), .A2(new_n636), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT60), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n634), .A2(KEYINPUT117), .ZN(new_n1150));
  XOR2_X1   g725(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n1151));
  INV_X1    g726(.A(KEYINPUT114), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1124), .A2(new_n1125), .A3(new_n1152), .A4(new_n971), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n1154));
  XNOR2_X1  g729(.A(KEYINPUT115), .B(KEYINPUT58), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(new_n763), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1072), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1072), .A2(new_n1156), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT116), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1039), .B2(new_n971), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1150), .B(new_n1151), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1150), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1151), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1146), .A2(new_n1149), .A3(new_n1162), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT61), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1142), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1027), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1040), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n956), .A2(new_n958), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n966), .A2(new_n1172), .A3(new_n1046), .A4(new_n1030), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT122), .ZN(new_n1174));
  AOI21_X1  g749(.A(G301), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT54), .B1(new_n1049), .B2(G171), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1171), .A2(new_n1174), .A3(G301), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1042), .A2(new_n1178), .A3(new_n1051), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1168), .A2(new_n1169), .A3(new_n1113), .A4(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1110), .A2(new_n1067), .A3(new_n804), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1183), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1105), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1184), .A2(new_n1109), .B1(new_n1093), .B2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1098), .A2(new_n1119), .A3(new_n1182), .A4(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(G290), .B(G1986), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n978), .B1(new_n977), .B2(new_n1188), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1187), .A2(KEYINPUT124), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT124), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n994), .B1(new_n1190), .B2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g767(.A1(new_n461), .A2(G227), .ZN(new_n1194));
  AND4_X1   g768(.A1(new_n672), .A2(new_n708), .A3(new_n712), .A4(new_n1194), .ZN(new_n1195));
  NAND2_X1  g769(.A1(new_n885), .A2(new_n894), .ZN(new_n1196));
  AND3_X1   g770(.A1(new_n1195), .A2(new_n1196), .A3(new_n950), .ZN(G308));
  NAND3_X1  g771(.A1(new_n1195), .A2(new_n1196), .A3(new_n950), .ZN(G225));
endmodule


