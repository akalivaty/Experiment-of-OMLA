//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT84), .ZN(new_n203));
  XOR2_X1   g002(.A(G57gat), .B(G85gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  INV_X1    g009(.A(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G162gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n216), .A2(new_n218), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(KEYINPUT79), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(G148gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n220), .B1(new_n224), .B2(new_n210), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT80), .B(G155gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n226), .B2(new_n215), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n219), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G113gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n229), .A2(KEYINPUT72), .A3(G120gat), .ZN(new_n230));
  INV_X1    g029(.A(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G127gat), .ZN(new_n232));
  INV_X1    g031(.A(G127gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G134gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n236));
  NOR2_X1   g035(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G120gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n229), .A2(G120gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT72), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n241), .A2(new_n242), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT1), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n234), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n239), .A2(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n228), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT82), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n248), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT73), .B(KEYINPUT1), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n244), .A2(new_n254), .A3(new_n255), .A4(new_n230), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT81), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n225), .A2(new_n227), .ZN(new_n259));
  INV_X1    g058(.A(new_n219), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT81), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n253), .A2(new_n262), .A3(new_n256), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n228), .A2(new_n249), .A3(KEYINPUT82), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n252), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G225gat), .A2(G233gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n208), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n252), .A2(new_n270), .A3(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n228), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n272), .A2(new_n258), .A3(new_n263), .A4(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n228), .A2(new_n249), .A3(KEYINPUT4), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n271), .A2(new_n275), .A3(new_n267), .A4(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n274), .A2(new_n258), .A3(new_n263), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n268), .B1(new_n279), .B2(new_n272), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n228), .A2(new_n249), .A3(KEYINPUT82), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT82), .B1(new_n228), .B2(new_n249), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT4), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n250), .A2(new_n270), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n280), .A2(new_n208), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n207), .B1(new_n278), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT6), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n278), .A2(new_n285), .A3(new_n207), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(new_n290), .B2(new_n286), .ZN(new_n291));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292));
  INV_X1    g091(.A(G211gat), .ZN(new_n293));
  INV_X1    g092(.A(G218gat), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295));
  OAI22_X1  g094(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(KEYINPUT22), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(KEYINPUT22), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G211gat), .B(G218gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n299), .B(new_n292), .C1(new_n296), .C2(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT65), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT65), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n310), .A2(new_n311), .A3(new_n315), .A4(new_n312), .ZN(new_n316));
  INV_X1    g115(.A(G169gat), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT23), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT23), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(G169gat), .B2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n314), .A2(new_n316), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n308), .A2(KEYINPUT66), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(G183gat), .A3(G190gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n329), .A3(new_n309), .ZN(new_n330));
  INV_X1    g129(.A(G183gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(KEYINPUT67), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT67), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G183gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g134(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(KEYINPUT68), .A2(G190gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n330), .B(new_n312), .C1(new_n335), .C2(new_n338), .ZN(new_n339));
  AND4_X1   g138(.A1(KEYINPUT25), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT70), .B(KEYINPUT28), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT69), .B1(new_n331), .B2(KEYINPUT27), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT69), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT27), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(G183gat), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n344), .A2(new_n347), .A3(new_n336), .A4(new_n337), .ZN(new_n348));
  AND3_X1   g147(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT27), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n351), .A2(KEYINPUT28), .A3(new_n336), .A4(new_n337), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NOR3_X1   g152(.A1(KEYINPUT71), .A2(G169gat), .A3(G176gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n322), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NOR4_X1   g155(.A1(KEYINPUT71), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n308), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n307), .B1(new_n342), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n324), .A2(new_n325), .B1(new_n339), .B2(new_n340), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n350), .B2(new_n352), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n362), .A2(new_n363), .A3(new_n306), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n304), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n360), .A3(new_n305), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n362), .A2(new_n363), .B1(KEYINPUT29), .B2(new_n306), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n366), .A2(new_n367), .A3(new_n303), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  NAND3_X1  g170(.A1(new_n365), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(KEYINPUT78), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT78), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n365), .A2(new_n368), .A3(new_n374), .A4(new_n371), .ZN(new_n375));
  INV_X1    g174(.A(new_n371), .ZN(new_n376));
  INV_X1    g175(.A(new_n368), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n303), .B1(new_n366), .B2(new_n367), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n376), .A2(KEYINPUT37), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n368), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n379), .A2(new_n380), .B1(new_n381), .B2(KEYINPUT37), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT38), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n373), .B(new_n375), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n291), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT38), .B1(new_n379), .B2(new_n380), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n377), .A2(KEYINPUT92), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(KEYINPUT37), .C1(new_n381), .C2(KEYINPUT92), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n386), .A2(KEYINPUT93), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT93), .B1(new_n386), .B2(new_n388), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT88), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT29), .B1(new_n301), .B2(new_n302), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n261), .B1(new_n393), .B2(KEYINPUT3), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT29), .B1(new_n228), .B2(new_n273), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n303), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT86), .B1(new_n395), .B2(new_n303), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n396), .A2(new_n397), .A3(G228gat), .A4(G233gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399));
  OAI221_X1 g198(.A(new_n394), .B1(KEYINPUT86), .B2(new_n399), .C1(new_n303), .C2(new_n395), .ZN(new_n400));
  AOI21_X1  g199(.A(G22gat), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(G22gat), .A3(new_n400), .ZN(new_n405));
  XNOR2_X1  g204(.A(G78gat), .B(G106gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT31), .B(G50gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n405), .B(new_n409), .C1(new_n401), .C2(new_n402), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n392), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n398), .A2(new_n400), .ZN(new_n412));
  INV_X1    g211(.A(G22gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT87), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n405), .A2(new_n409), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT88), .A4(new_n403), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n409), .B1(new_n414), .B2(new_n405), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n385), .A2(new_n391), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n373), .A2(new_n422), .A3(new_n375), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n365), .A2(new_n368), .A3(KEYINPUT30), .A4(new_n371), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n379), .A2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT90), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT90), .B1(new_n423), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT40), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n283), .A2(new_n275), .A3(new_n284), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n268), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n207), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n252), .A2(new_n264), .A3(new_n265), .A4(new_n267), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT39), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n268), .B2(new_n430), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n429), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n286), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n430), .A2(new_n268), .ZN(new_n439));
  INV_X1    g238(.A(new_n435), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(KEYINPUT40), .A3(new_n207), .A4(new_n432), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n437), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT91), .B1(new_n428), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n425), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT90), .ZN(new_n448));
  AND4_X1   g247(.A1(KEYINPUT91), .A2(new_n443), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n421), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT94), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT94), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n421), .B(new_n452), .C1(new_n444), .C2(new_n449), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n342), .A2(new_n360), .A3(new_n257), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n249), .B1(new_n362), .B2(new_n363), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G227gat), .A2(G233gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT64), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT75), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT34), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n457), .A2(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT74), .B(G71gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(G99gat), .ZN(new_n466));
  XOR2_X1   g265(.A(G15gat), .B(G43gat), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n455), .A2(new_n456), .A3(new_n459), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(KEYINPUT32), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n461), .A2(new_n462), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n469), .B(KEYINPUT32), .C1(new_n470), .C2(new_n468), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n475), .B1(new_n473), .B2(new_n476), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n464), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n479), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n463), .A3(new_n477), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n480), .A2(new_n482), .B1(KEYINPUT76), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n480), .A2(new_n482), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n419), .B1(new_n411), .B2(new_n417), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n286), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n283), .A2(new_n284), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n275), .A2(new_n208), .A3(new_n267), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n493), .A2(new_n495), .B1(new_n269), .B2(new_n277), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT85), .B1(new_n496), .B2(new_n207), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT6), .B1(new_n496), .B2(new_n207), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n492), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n287), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n490), .B1(new_n501), .B2(new_n445), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT89), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n489), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n488), .ZN(new_n505));
  INV_X1    g304(.A(new_n490), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n445), .B1(new_n499), .B2(new_n287), .ZN(new_n507));
  OAI22_X1  g306(.A1(new_n505), .A2(new_n484), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT89), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n454), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n480), .A2(new_n482), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n490), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n507), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n512), .A2(new_n490), .A3(new_n428), .ZN(new_n515));
  INV_X1    g314(.A(new_n291), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n514), .A2(KEYINPUT35), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT97), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT97), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT15), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n526), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n524), .B1(KEYINPUT95), .B2(new_n522), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT96), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT96), .ZN(new_n542));
  AOI211_X1 g341(.A(new_n542), .B(new_n539), .C1(new_n536), .C2(new_n537), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n533), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(G1gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G1gat), .B2(new_n545), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G8gat), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n549), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n544), .A2(new_n551), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n521), .B(new_n550), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n544), .B(new_n549), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n521), .B(KEYINPUT13), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n544), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT17), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n553), .A3(new_n552), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(KEYINPUT18), .A3(new_n521), .A4(new_n550), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT11), .B(G169gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n571), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n558), .A2(new_n565), .A3(new_n573), .A4(new_n561), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G190gat), .B(G218gat), .Z(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n578));
  NAND2_X1  g377(.A1(G85gat), .A2(G92gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT7), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT100), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n579), .B2(KEYINPUT7), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(KEYINPUT101), .A3(G85gat), .A4(G92gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT100), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n579), .A2(new_n586), .A3(KEYINPUT7), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n581), .A2(new_n583), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G99gat), .B(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n594), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n552), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n578), .B1(new_n599), .B2(new_n555), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n563), .A2(KEYINPUT102), .A3(new_n552), .A4(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n598), .ZN(new_n603));
  AND2_X1   g402(.A1(G232gat), .A2(G233gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n544), .A2(new_n603), .B1(KEYINPUT41), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n577), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G134gat), .B(G162gat), .Z(new_n608));
  NOR2_X1   g407(.A1(new_n604), .A2(KEYINPUT41), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n602), .A2(new_n605), .A3(new_n577), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n607), .A2(KEYINPUT103), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n610), .B(KEYINPUT103), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n602), .A2(new_n605), .A3(new_n577), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(new_n606), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G71gat), .A2(G78gat), .ZN(new_n618));
  OR2_X1    g417(.A1(G71gat), .A2(G78gat), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT9), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(G57gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(G64gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(G64gat), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n624), .B2(KEYINPUT98), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n626), .A2(new_n622), .A3(G64gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n621), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G64gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(G57gat), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT9), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n631), .A2(new_n618), .A3(new_n619), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n549), .B1(KEYINPUT21), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT99), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G231gat), .A2(G233gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n233), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n636), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G155gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(G183gat), .B(G211gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n642), .B(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT104), .B1(new_n617), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n613), .A2(new_n616), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n598), .A2(new_n633), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n634), .A2(new_n596), .A3(new_n597), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n634), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G230gat), .A2(G233gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(KEYINPUT105), .A3(new_n660), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n654), .A2(new_n655), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(G230gat), .A3(G233gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n661), .A2(new_n667), .A3(new_n671), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n520), .A2(new_n575), .A3(new_n653), .A4(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(new_n500), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT106), .B(G1gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1324gat));
  INV_X1    g479(.A(new_n428), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT16), .B(G8gat), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT107), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT42), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT107), .B(new_n686), .C1(new_n682), .C2(new_n683), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(G8gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n677), .B2(new_n489), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n512), .A2(G15gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n677), .B2(new_n691), .ZN(G1326gat));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n506), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  NOR2_X1   g494(.A1(new_n649), .A2(new_n675), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n520), .A2(new_n575), .A3(new_n617), .A4(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(G29gat), .A3(new_n500), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n508), .B1(new_n451), .B2(new_n453), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n518), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n703), .B2(new_n650), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n650), .A2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n509), .A2(new_n504), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n451), .B2(new_n453), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n707), .B2(new_n518), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n572), .A2(KEYINPUT109), .A3(new_n574), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT109), .B1(new_n572), .B2(new_n574), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n696), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n704), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G29gat), .B1(new_n713), .B2(new_n500), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n700), .A2(new_n714), .ZN(G1328gat));
  NOR3_X1   g514(.A1(new_n697), .A2(G36gat), .A3(new_n681), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  OAI21_X1  g516(.A(G36gat), .B1(new_n713), .B2(new_n681), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1329gat));
  NOR2_X1   g518(.A1(new_n697), .A2(new_n512), .ZN(new_n720));
  INV_X1    g519(.A(new_n489), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n720), .A2(G43gat), .B1(new_n713), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g523(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n725));
  INV_X1    g524(.A(new_n575), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n510), .B2(new_n519), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n727), .A2(new_n728), .A3(new_n617), .A4(new_n696), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n506), .A2(G50gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n725), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT111), .B1(new_n713), .B2(new_n506), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G50gat), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n713), .A2(KEYINPUT111), .A3(new_n506), .ZN(new_n734));
  OAI211_X1 g533(.A(KEYINPUT48), .B(new_n731), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(G50gat), .B1(new_n713), .B2(new_n506), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT48), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n735), .A2(new_n739), .ZN(G1331gat));
  INV_X1    g539(.A(new_n703), .ZN(new_n741));
  INV_X1    g540(.A(new_n711), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n653), .A2(new_n675), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n500), .B(KEYINPUT112), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g547(.A1(new_n744), .A2(new_n681), .ZN(new_n749));
  NOR2_X1   g548(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n750));
  AND2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n749), .B2(new_n750), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n744), .B2(new_n489), .ZN(new_n754));
  INV_X1    g553(.A(G71gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n511), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n744), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g557(.A1(new_n745), .A2(new_n490), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n711), .A2(new_n649), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT113), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(new_n675), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n704), .A2(new_n708), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n500), .ZN(new_n765));
  OAI211_X1 g564(.A(new_n617), .B(new_n762), .C1(new_n702), .C2(new_n518), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n676), .A2(new_n500), .A3(G85gat), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT114), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n765), .B1(new_n770), .B2(new_n772), .ZN(G1336gat));
  INV_X1    g572(.A(new_n770), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n681), .A2(new_n676), .A3(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n704), .A2(new_n708), .A3(new_n428), .A4(new_n763), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G92gat), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n777), .A2(KEYINPUT115), .A3(G92gat), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT115), .B1(new_n777), .B2(G92gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n767), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n783), .A3(KEYINPUT51), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n785), .A2(new_n786), .A3(new_n775), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n781), .A2(new_n782), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n780), .B1(new_n788), .B2(new_n779), .ZN(G1337gat));
  OAI21_X1  g588(.A(G99gat), .B1(new_n764), .B2(new_n489), .ZN(new_n790));
  OR3_X1    g589(.A1(new_n512), .A2(new_n676), .A3(G99gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n770), .B2(new_n791), .ZN(G1338gat));
  NOR3_X1   g591(.A1(new_n506), .A2(new_n676), .A3(G106gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n785), .A2(new_n786), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT117), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n785), .A2(new_n796), .A3(new_n786), .A4(new_n793), .ZN(new_n797));
  OAI21_X1  g596(.A(G106gat), .B1(new_n764), .B2(new_n506), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n774), .B2(new_n793), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n663), .A2(new_n805), .A3(new_n664), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n661), .A2(KEYINPUT54), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n659), .A2(new_n660), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n672), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n804), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n808), .A2(new_n809), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n672), .A4(new_n806), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n811), .A2(new_n674), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT118), .A4(new_n674), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n711), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n521), .B1(new_n564), .B2(new_n550), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n559), .A2(new_n560), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n570), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n574), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n675), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n617), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n816), .A2(new_n817), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n613), .A2(new_n616), .A3(new_n822), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n647), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n653), .A2(new_n676), .A3(new_n742), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n746), .ZN(new_n831));
  INV_X1    g630(.A(new_n513), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n831), .A2(new_n832), .A3(new_n428), .ZN(new_n833));
  AOI21_X1  g632(.A(G113gat), .B1(new_n833), .B2(new_n711), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n490), .B1(new_n828), .B2(new_n829), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n835), .A2(new_n501), .A3(new_n511), .A4(new_n681), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n836), .A2(new_n229), .A3(new_n726), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n834), .A2(new_n837), .ZN(G1340gat));
  AOI21_X1  g637(.A(G120gat), .B1(new_n833), .B2(new_n675), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n836), .A2(new_n240), .A3(new_n676), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(G1341gat));
  NAND3_X1  g640(.A1(new_n833), .A2(new_n233), .A3(new_n649), .ZN(new_n842));
  OAI21_X1  g641(.A(G127gat), .B1(new_n836), .B2(new_n647), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(G1342gat));
  NAND3_X1  g643(.A1(new_n833), .A2(new_n231), .A3(new_n617), .ZN(new_n845));
  OR2_X1    g644(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n846));
  OAI21_X1  g645(.A(G134gat), .B1(new_n836), .B2(new_n650), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(KEYINPUT56), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(G1343gat));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n721), .A2(new_n506), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n681), .A3(new_n746), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n726), .A2(G141gat), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n721), .A2(new_n500), .A3(new_n428), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n830), .B2(new_n490), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n506), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n575), .A2(new_n811), .A3(new_n674), .A4(new_n813), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n617), .B1(new_n861), .B2(new_n823), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n647), .B1(new_n827), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n860), .B1(new_n829), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n575), .B(new_n856), .C1(new_n857), .C2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n221), .A2(new_n223), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n855), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI211_X1 g668(.A(KEYINPUT119), .B(new_n855), .C1(new_n865), .C2(new_n866), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n711), .B(new_n856), .C1(new_n857), .C2(new_n864), .ZN(new_n871));
  INV_X1    g670(.A(new_n852), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n871), .A2(new_n866), .B1(new_n872), .B2(new_n853), .ZN(new_n873));
  OAI22_X1  g672(.A1(new_n869), .A2(new_n870), .B1(new_n873), .B2(new_n850), .ZN(G1344gat));
  AOI21_X1  g673(.A(new_n860), .B1(new_n828), .B2(new_n829), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n826), .A2(new_n814), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n647), .B1(new_n862), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n648), .A2(new_n726), .A3(new_n652), .A4(new_n676), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n879), .B2(new_n490), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n856), .A2(new_n675), .ZN(new_n882));
  OAI21_X1  g681(.A(G148gat), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT59), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n675), .B(new_n856), .C1(new_n857), .C2(new_n864), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n209), .A2(KEYINPUT59), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n885), .B2(new_n887), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n872), .A2(new_n209), .A3(new_n675), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1345gat));
  NAND3_X1  g691(.A1(new_n872), .A2(new_n226), .A3(new_n649), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n856), .B1(new_n857), .B2(new_n864), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n647), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n895), .B2(new_n226), .ZN(G1346gat));
  NOR3_X1   g695(.A1(new_n894), .A2(new_n215), .A3(new_n650), .ZN(new_n897));
  AOI21_X1  g696(.A(G162gat), .B1(new_n872), .B2(new_n617), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(G1347gat));
  OR2_X1    g698(.A1(new_n746), .A2(new_n681), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n512), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n835), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n902), .A2(new_n317), .A3(new_n726), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n501), .B1(new_n828), .B2(new_n829), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n428), .B1(new_n904), .B2(KEYINPUT121), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  AOI211_X1 g705(.A(new_n906), .B(new_n501), .C1(new_n828), .C2(new_n829), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n832), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n711), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n903), .B1(new_n909), .B2(new_n317), .ZN(G1348gat));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n318), .A3(new_n675), .ZN(new_n911));
  OAI21_X1  g710(.A(G176gat), .B1(new_n902), .B2(new_n676), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  NAND2_X1  g712(.A1(new_n830), .A2(new_n500), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n681), .B1(new_n914), .B2(new_n906), .ZN(new_n915));
  INV_X1    g714(.A(new_n907), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n649), .A2(new_n351), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n915), .A2(new_n513), .A3(new_n916), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n335), .B1(new_n902), .B2(new_n647), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g720(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n922));
  NAND2_X1  g721(.A1(KEYINPUT122), .A2(KEYINPUT60), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n919), .A2(KEYINPUT122), .A3(KEYINPUT60), .A4(new_n920), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n902), .B2(new_n650), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n928), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(KEYINPUT61), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n927), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n650), .A2(new_n338), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT123), .B1(new_n908), .B2(new_n934), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n908), .A2(KEYINPUT123), .A3(new_n934), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n931), .B(new_n933), .C1(new_n935), .C2(new_n936), .ZN(G1351gat));
  NAND2_X1  g736(.A1(new_n830), .A2(new_n859), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n879), .A2(new_n490), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(new_n858), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n900), .A2(new_n721), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n941), .A2(KEYINPUT125), .A3(new_n575), .A4(new_n942), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n575), .B(new_n942), .C1(new_n875), .C2(new_n880), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(G197gat), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n742), .A2(G197gat), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n915), .A2(new_n851), .A3(new_n916), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT126), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n952), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1352gat));
  NOR2_X1   g753(.A1(new_n676), .A2(G204gat), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n915), .A2(new_n851), .A3(new_n916), .A4(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(G204gat), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n881), .A2(new_n721), .A3(new_n900), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n675), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n956), .B1(new_n959), .B2(KEYINPUT62), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n956), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n961));
  OAI21_X1  g760(.A(KEYINPUT127), .B1(new_n956), .B2(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G1353gat));
  NOR4_X1   g762(.A1(new_n905), .A2(new_n907), .A3(new_n506), .A4(new_n721), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n293), .A3(new_n649), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n958), .A2(new_n649), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n966), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n966), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(G1354gat));
  NAND3_X1  g768(.A1(new_n964), .A2(new_n294), .A3(new_n617), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n958), .A2(new_n617), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n970), .B1(new_n972), .B2(new_n294), .ZN(G1355gat));
endmodule


