//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G113), .ZN(new_n191));
  AND2_X1   g005(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n191), .A2(KEYINPUT2), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n188), .B(new_n190), .C1(new_n192), .C2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(new_n190), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT2), .B(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(new_n199), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n203), .B2(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n200), .A2(KEYINPUT66), .A3(G137), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n200), .A2(G137), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(KEYINPUT11), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n207), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(G131), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  AND2_X1   g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  INV_X1    g034(.A(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n219), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n226));
  XNOR2_X1  g040(.A(G143), .B(G146), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n218), .B(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(G143), .B2(new_n221), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n223), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n221), .A2(G143), .ZN(new_n233));
  OAI22_X1  g047(.A1(new_n231), .A2(new_n219), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n218), .B1(new_n234), .B2(new_n225), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n198), .B1(new_n217), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n205), .B1(new_n204), .B2(new_n199), .ZN(new_n238));
  AOI211_X1 g052(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n203), .C2(G134), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n210), .A2(new_n211), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n212), .A2(KEYINPUT11), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n214), .ZN(new_n246));
  OAI211_X1 g060(.A(KEYINPUT67), .B(G131), .C1(new_n240), .C2(new_n243), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT64), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n227), .B2(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n227), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n222), .A2(new_n224), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n255), .A3(KEYINPUT64), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n250), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n246), .A2(new_n247), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n237), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XOR2_X1   g077(.A(new_n263), .B(KEYINPUT27), .Z(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n237), .A2(new_n258), .A3(KEYINPUT69), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT69), .B1(new_n237), .B2(new_n258), .ZN(new_n269));
  INV_X1    g083(.A(new_n198), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n234), .A2(new_n225), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n217), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n258), .B2(new_n272), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n261), .B(new_n267), .C1(new_n274), .C2(new_n260), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n258), .A2(new_n272), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n217), .A2(new_n236), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n258), .A2(KEYINPUT30), .A3(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n278), .A2(new_n198), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n259), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n237), .A2(new_n258), .A3(KEYINPUT69), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n266), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n275), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n266), .A2(new_n287), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n261), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n258), .A2(new_n279), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n198), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n283), .A2(new_n292), .A3(new_n284), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n290), .B1(new_n293), .B2(KEYINPUT28), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT71), .B1(new_n294), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n268), .A2(new_n269), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n260), .B1(new_n298), .B2(new_n292), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n296), .B(new_n297), .C1(new_n299), .C2(new_n290), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n288), .A2(new_n295), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G472), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n278), .A2(new_n198), .A3(new_n280), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n298), .A3(new_n267), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n304), .A2(new_n298), .A3(KEYINPUT31), .A4(new_n267), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n261), .B1(new_n274), .B2(new_n260), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n266), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT70), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n307), .A2(new_n308), .B1(new_n310), .B2(new_n266), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT32), .B1(new_n318), .B2(new_n315), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n301), .A2(new_n321), .A3(G472), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n303), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G469), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G140), .ZN(new_n325));
  INV_X1    g139(.A(G953), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(G227), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n325), .B(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n329));
  INV_X1    g143(.A(G104), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT3), .B1(new_n330), .B2(G107), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT3), .ZN(new_n332));
  INV_X1    g146(.A(G107), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(G104), .ZN(new_n334));
  INV_X1    g148(.A(G101), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(G107), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n331), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n330), .A2(G107), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n333), .A2(G104), .ZN(new_n339));
  OAI21_X1  g153(.A(G101), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n342), .A4(new_n228), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n334), .A3(new_n336), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G101), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n347), .A3(G101), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n257), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n350));
  INV_X1    g164(.A(new_n225), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT1), .B1(new_n223), .B2(G146), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT79), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT79), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n222), .A2(new_n354), .A3(KEYINPUT1), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(G128), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n351), .B1(new_n356), .B2(new_n253), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n350), .B1(new_n357), .B2(new_n341), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n343), .A2(new_n349), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n246), .B2(new_n247), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n246), .A2(new_n360), .A3(new_n247), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n328), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n246), .A2(new_n247), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n341), .A2(new_n234), .A3(new_n225), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n357), .B2(new_n341), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n365), .A2(new_n366), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n246), .A3(new_n247), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT12), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n368), .A2(new_n246), .A3(new_n247), .A4(new_n369), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT83), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n328), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n359), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n343), .A2(new_n349), .A3(new_n358), .A4(KEYINPUT84), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n365), .A3(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n343), .A2(new_n349), .A3(new_n358), .ZN(new_n383));
  INV_X1    g197(.A(new_n361), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n363), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n378), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n324), .B(new_n297), .C1(new_n377), .C2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n376), .A2(new_n385), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n328), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n364), .A2(new_n382), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(G469), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n324), .A2(new_n297), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n387), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT9), .B(G234), .ZN(new_n395));
  OAI21_X1  g209(.A(G221), .B1(new_n395), .B2(G902), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n400));
  OAI21_X1  g214(.A(G131), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n400), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(new_n208), .A3(new_n398), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT17), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G125), .ZN(new_n406));
  NOR3_X1   g220(.A1(new_n406), .A2(KEYINPUT16), .A3(G140), .ZN(new_n407));
  XNOR2_X1  g221(.A(G125), .B(G140), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G146), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n409), .A2(G146), .ZN(new_n411));
  OAI211_X1 g225(.A(KEYINPUT17), .B(G131), .C1(new_n399), .C2(new_n400), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n405), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G113), .B(G122), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(new_n330), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n408), .B(new_n221), .ZN(new_n416));
  OAI211_X1 g230(.A(KEYINPUT18), .B(G131), .C1(new_n399), .C2(new_n400), .ZN(new_n417));
  NAND2_X1  g231(.A1(KEYINPUT18), .A2(G131), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n402), .A2(new_n398), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n413), .A2(new_n415), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n415), .B1(new_n413), .B2(new_n420), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n297), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G475), .ZN(new_n425));
  INV_X1    g239(.A(new_n420), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n408), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT19), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n428), .B(KEYINPUT88), .C1(new_n429), .C2(new_n408), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n408), .A2(new_n427), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n221), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n221), .B(new_n407), .C1(KEYINPUT16), .C2(new_n408), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n401), .B2(new_n403), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n426), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n421), .B1(new_n437), .B2(new_n415), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n439));
  NOR2_X1   g253(.A1(G475), .A2(G902), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n425), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n189), .A2(G122), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT89), .B(G122), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n444), .B1(new_n445), .B2(new_n189), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(new_n445), .B2(new_n189), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n447), .A3(G107), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n333), .A2(KEYINPUT14), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n223), .A2(G128), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n219), .A2(G143), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT91), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n453), .A2(G134), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(G134), .B1(new_n453), .B2(new_n455), .ZN(new_n457));
  OAI221_X1 g271(.A(new_n448), .B1(new_n446), .B2(new_n449), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n457), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n223), .A2(KEYINPUT13), .A3(G128), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT90), .A3(new_n451), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT13), .B1(new_n223), .B2(G128), .ZN(new_n462));
  OAI221_X1 g276(.A(G134), .B1(KEYINPUT90), .B2(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n446), .A2(G107), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n446), .A2(G107), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n459), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G217), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n395), .A2(new_n467), .A3(G953), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n458), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n458), .B2(new_n466), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n297), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G478), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(KEYINPUT15), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI221_X1 g289(.A(new_n297), .B1(KEYINPUT15), .B2(new_n473), .C1(new_n470), .C2(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(G234), .A2(G237), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n478), .A2(G952), .A3(new_n326), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n478), .A2(G902), .A3(G953), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(G898), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n443), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  OAI21_X1  g298(.A(G210), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G110), .B(G122), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT8), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT5), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(G113), .C1(KEYINPUT5), .C2(new_n188), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n342), .B1(new_n194), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n490), .A2(new_n194), .A3(new_n340), .A4(new_n337), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n337), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n198), .A2(new_n348), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n492), .B(new_n487), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n271), .A2(new_n406), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n250), .A2(new_n256), .A3(G125), .A4(new_n252), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n500));
  INV_X1    g314(.A(G224), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(G953), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n494), .A2(new_n497), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n498), .B2(new_n499), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n502), .A2(KEYINPUT7), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n297), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n511));
  INV_X1    g325(.A(new_n487), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT6), .A3(new_n497), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n506), .A2(new_n507), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n511), .A2(new_n516), .A3(new_n512), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT85), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT85), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n514), .A2(new_n515), .A3(new_n520), .A4(new_n517), .ZN(new_n521));
  AOI211_X1 g335(.A(new_n486), .B(new_n510), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n510), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n485), .B(KEYINPUT86), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n483), .B(new_n484), .C1(new_n522), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n397), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n219), .A2(G119), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n187), .A2(G128), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n530), .A2(new_n531), .A3(new_n529), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT24), .B(G110), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT23), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n531), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT23), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT74), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n530), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(G110), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n409), .A2(G146), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n537), .B(new_n545), .C1(new_n546), .C2(new_n435), .ZN(new_n547));
  XNOR2_X1  g361(.A(KEYINPUT22), .B(G137), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(G221), .A2(G234), .ZN(new_n550));
  OAI21_X1  g364(.A(KEYINPUT76), .B1(new_n550), .B2(G953), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT76), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n552), .A2(new_n326), .A3(G221), .A4(G234), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT77), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n551), .B2(new_n553), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n557), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n548), .A3(new_n555), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n539), .A2(new_n543), .ZN(new_n562));
  INV_X1    g376(.A(new_n530), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G110), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n564), .A2(new_n565), .A3(new_n531), .A4(new_n540), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n530), .A2(new_n531), .A3(new_n529), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n535), .B1(new_n567), .B2(new_n532), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n408), .A2(new_n221), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n409), .B2(G146), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n569), .A2(KEYINPUT75), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT75), .B1(new_n569), .B2(new_n571), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n547), .B(new_n561), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n547), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n569), .A2(new_n571), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(KEYINPUT75), .A3(new_n571), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n558), .A2(new_n560), .A3(KEYINPUT78), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT78), .B1(new_n558), .B2(new_n560), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n574), .B(new_n297), .C1(new_n580), .C2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n547), .B1(new_n572), .B2(new_n573), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n582), .B2(new_n583), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n589), .A2(KEYINPUT25), .A3(new_n297), .A4(new_n574), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n467), .B1(G234), .B2(new_n297), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n574), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n592), .A2(G902), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n591), .A2(new_n592), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n323), .A2(new_n528), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  NAND2_X1  g412(.A1(new_n519), .A2(new_n521), .ZN(new_n599));
  INV_X1    g413(.A(new_n510), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n599), .A2(KEYINPUT92), .A3(new_n485), .A4(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(new_n485), .B2(new_n523), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n522), .A2(KEYINPUT92), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n484), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n472), .A2(new_n473), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT93), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n470), .B2(new_n471), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n458), .A2(new_n466), .ZN(new_n610));
  INV_X1    g424(.A(new_n468), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n469), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n297), .A2(G478), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n605), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n443), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(new_n443), .A3(KEYINPUT94), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n604), .A2(new_n623), .A3(new_n482), .ZN(new_n624));
  OAI21_X1  g438(.A(G472), .B1(new_n318), .B2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n312), .A2(new_n316), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n394), .A2(new_n596), .A3(new_n396), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n624), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT95), .ZN(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT34), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n523), .A2(new_n485), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT92), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n523), .A2(new_n485), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n638), .A3(new_n601), .ZN(new_n639));
  INV_X1    g453(.A(new_n482), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n413), .A2(new_n420), .ZN(new_n642));
  INV_X1    g456(.A(new_n415), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n644), .B2(new_n421), .ZN(new_n645));
  INV_X1    g459(.A(G475), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n424), .A2(KEYINPUT96), .A3(G475), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n438), .A2(new_n440), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT20), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n649), .A2(new_n653), .A3(new_n477), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n639), .A2(new_n484), .A3(new_n640), .A4(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(new_n627), .A3(new_n628), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT98), .B(G107), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NAND2_X1  g474(.A1(new_n588), .A2(KEYINPUT99), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT36), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(new_n547), .C1(new_n572), .C2(new_n573), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n662), .B1(new_n661), .B2(new_n664), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n595), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT100), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n591), .A2(new_n592), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n670), .B(new_n595), .C1(new_n665), .C2(new_n666), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n397), .A2(new_n527), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n627), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  NAND3_X1  g491(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n678));
  INV_X1    g492(.A(new_n479), .ZN(new_n679));
  INV_X1    g493(.A(new_n480), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n679), .B1(new_n680), .B2(G900), .ZN(new_n681));
  AND4_X1   g495(.A1(new_n653), .A2(new_n649), .A3(new_n477), .A4(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n604), .A2(new_n397), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n323), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  NOR2_X1   g500(.A1(new_n526), .A2(new_n522), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  INV_X1    g502(.A(new_n484), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n443), .A2(new_n477), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n688), .A2(new_n689), .A3(new_n678), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n681), .B(KEYINPUT39), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n394), .A2(new_n396), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n691), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n281), .A2(new_n285), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n266), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n297), .B1(new_n293), .B2(new_n267), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n320), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT101), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n696), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n223), .ZN(G45));
  NAND3_X1  g518(.A1(new_n618), .A2(new_n443), .A3(new_n681), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n678), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n604), .A2(new_n397), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n313), .B1(new_n312), .B2(new_n316), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n318), .A2(KEYINPUT32), .A3(new_n315), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n322), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n321), .B1(new_n301), .B2(G472), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n708), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  NAND2_X1  g528(.A1(new_n382), .A2(new_n385), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n715), .A2(new_n328), .B1(new_n364), .B2(new_n376), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n716), .B2(G902), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n387), .A3(new_n396), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(KEYINPUT102), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n387), .A3(new_n720), .A4(new_n396), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n719), .A2(new_n596), .A3(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n323), .A2(new_n624), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT41), .B(G113), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT103), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n723), .B(new_n725), .ZN(G15));
  NAND3_X1  g540(.A1(new_n719), .A2(new_n596), .A3(new_n721), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n655), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n323), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT104), .B1(new_n728), .B2(new_n323), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n189), .ZN(G18));
  INV_X1    g548(.A(new_n604), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n678), .A2(new_n483), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n721), .A3(new_n736), .A4(new_n719), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n323), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  NOR2_X1   g554(.A1(new_n604), .A2(new_n690), .ZN(new_n741));
  INV_X1    g555(.A(new_n261), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n266), .B1(new_n299), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n309), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n316), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n625), .A2(new_n745), .A3(new_n640), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n722), .A2(new_n741), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  AND2_X1   g562(.A1(new_n719), .A2(new_n721), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n667), .A2(KEYINPUT100), .B1(new_n591), .B2(new_n592), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n705), .B1(new_n750), .B2(new_n671), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n625), .A2(new_n751), .A3(new_n745), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n752), .A3(new_n735), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT105), .B(G125), .Z(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G27));
  AOI22_X1  g569(.A1(KEYINPUT83), .A2(new_n374), .B1(new_n371), .B2(new_n372), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n756), .A2(new_n370), .B1(new_n362), .B2(new_n363), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT106), .B1(new_n757), .B2(new_n378), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n388), .A2(new_n759), .A3(new_n328), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n758), .A2(new_n760), .A3(G469), .A4(new_n390), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n387), .A3(new_n393), .ZN(new_n762));
  INV_X1    g576(.A(new_n396), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n689), .ZN(new_n764));
  AND4_X1   g578(.A1(new_n596), .A2(new_n762), .A3(new_n687), .A4(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n323), .A2(new_n706), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n323), .A2(KEYINPUT42), .A3(new_n706), .A4(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  OAI211_X1 g585(.A(new_n682), .B(new_n765), .C1(new_n711), .C2(new_n712), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  AOI21_X1  g587(.A(KEYINPUT111), .B1(new_n627), .B2(new_n678), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n627), .A2(new_n678), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n651), .A2(new_n652), .B1(G475), .B2(new_n424), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n618), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT43), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT110), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n774), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(KEYINPUT44), .ZN(new_n784));
  INV_X1    g598(.A(new_n687), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n689), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n783), .B1(new_n782), .B2(KEYINPUT44), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT113), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n788), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n790), .A2(new_n791), .A3(new_n786), .A4(new_n784), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n389), .B2(new_n390), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n324), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n758), .A2(new_n760), .A3(KEYINPUT45), .A4(new_n390), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n392), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT46), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT107), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n387), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n799), .A2(KEYINPUT108), .A3(new_n387), .A4(new_n800), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n796), .A2(KEYINPUT46), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT109), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n807), .A2(new_n396), .A3(new_n692), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n782), .A2(KEYINPUT44), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n789), .A2(new_n792), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G137), .ZN(G39));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n396), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(KEYINPUT47), .A3(new_n396), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n323), .ZN(new_n817));
  INV_X1    g631(.A(new_n786), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n596), .A3(new_n705), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  NAND2_X1  g635(.A1(new_n596), .A2(new_n479), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n780), .A2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n625), .A2(new_n745), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n689), .A3(new_n688), .A4(new_n749), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT50), .Z(new_n828));
  NAND2_X1  g642(.A1(new_n749), .A2(new_n786), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n822), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n702), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n618), .A2(new_n443), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n829), .A2(new_n679), .A3(new_n780), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n678), .A3(new_n824), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n828), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n717), .A2(new_n387), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n814), .B(new_n815), .C1(new_n396), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n825), .A2(new_n818), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT51), .ZN(new_n842));
  MUX2_X1   g656(.A(new_n477), .B(new_n618), .S(new_n443), .Z(new_n843));
  AND4_X1   g657(.A1(new_n484), .A2(new_n843), .A3(new_n785), .A4(new_n640), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n844), .A2(new_n629), .B1(new_n673), .B2(new_n674), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n723), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n747), .B1(new_n817), .B2(new_n737), .ZN(new_n847));
  INV_X1    g661(.A(new_n597), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n752), .A2(new_n687), .A3(new_n762), .A4(new_n764), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n475), .A2(new_n476), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n653), .A2(new_n851), .A3(new_n649), .A4(new_n681), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n687), .A2(new_n852), .A3(new_n678), .A4(new_n484), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n853), .A2(new_n397), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n854), .B1(new_n711), .B2(new_n712), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n772), .A2(new_n850), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n768), .B2(new_n769), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n729), .B(new_n730), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n849), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n762), .A2(new_n672), .A3(new_n396), .A4(new_n681), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n701), .A2(new_n861), .A3(new_n741), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n685), .A2(new_n713), .A3(new_n862), .A4(new_n753), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT52), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n735), .A2(new_n721), .A3(new_n719), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n865), .A2(new_n752), .B1(new_n323), .B2(new_n684), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n860), .B1(new_n320), .B2(new_n700), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n867), .A2(new_n741), .B1(new_n323), .B2(new_n708), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT52), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g685(.A1(new_n859), .A2(new_n871), .A3(KEYINPUT53), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n864), .A2(new_n870), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n873), .B1(new_n864), .B2(new_n870), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n859), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n878));
  OAI211_X1 g692(.A(KEYINPUT54), .B(new_n872), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n878), .B1(new_n876), .B2(new_n859), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n864), .A2(new_n870), .A3(KEYINPUT53), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT116), .B1(new_n859), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n864), .A2(new_n870), .A3(KEYINPUT53), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n625), .A2(new_n745), .A3(new_n640), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n727), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n738), .A2(new_n323), .B1(new_n885), .B2(new_n741), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n597), .A3(new_n723), .A4(new_n845), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n733), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n883), .A2(new_n888), .A3(new_n889), .A4(new_n857), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n880), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n835), .A2(new_n323), .A3(new_n596), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n896));
  XOR2_X1   g710(.A(KEYINPUT118), .B(KEYINPUT48), .Z(new_n897));
  NAND3_X1  g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(G952), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n899), .B(G953), .C1(new_n826), .C2(new_n865), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n898), .B(new_n900), .C1(new_n623), .C2(new_n832), .ZN(new_n901));
  AOI211_X1 g715(.A(KEYINPUT118), .B(KEYINPUT48), .C1(new_n895), .C2(new_n896), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n879), .A2(new_n893), .A3(new_n903), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n842), .A2(new_n904), .B1(G952), .B2(G953), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n779), .A2(new_n763), .A3(new_n689), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n596), .C1(KEYINPUT49), .C2(new_n838), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(KEYINPUT49), .B2(new_n838), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n702), .A2(new_n688), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT114), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n910), .ZN(G75));
  NOR2_X1   g725(.A1(new_n326), .A2(G952), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT120), .Z(new_n913));
  AOI21_X1  g727(.A(new_n297), .B1(new_n880), .B2(new_n891), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(new_n524), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n514), .A2(new_n517), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n515), .ZN(new_n917));
  XNOR2_X1  g731(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT56), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n913), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n914), .A2(G210), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n923), .B2(new_n920), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(G51));
  AND3_X1   g739(.A1(new_n880), .A2(new_n891), .A3(new_n892), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n892), .B1(new_n880), .B2(new_n891), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n392), .B(KEYINPUT57), .Z(new_n929));
  OAI22_X1  g743(.A1(new_n928), .A2(new_n929), .B1(new_n377), .B2(new_n386), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n914), .A2(new_n795), .A3(new_n794), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n912), .B1(new_n930), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  INV_X1    g747(.A(new_n438), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n933), .A2(KEYINPUT121), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n912), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n933), .B2(new_n934), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT121), .B1(new_n933), .B2(new_n934), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(G60));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT59), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n609), .A2(new_n615), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n880), .A2(new_n891), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT54), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n943), .B1(new_n945), .B2(new_n893), .ZN(new_n946));
  INV_X1    g760(.A(new_n913), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(KEYINPUT122), .B(new_n913), .C1(new_n928), .C2(new_n943), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n879), .A2(new_n893), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n942), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n616), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(G63));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n954));
  NAND2_X1  g768(.A1(G217), .A2(G902), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n880), .B2(new_n891), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n954), .B(new_n913), .C1(new_n957), .C2(new_n594), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n956), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n882), .A2(new_n890), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n871), .A2(KEYINPUT115), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n864), .A2(new_n870), .A3(new_n873), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n859), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT53), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n961), .B1(new_n962), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n947), .B1(new_n968), .B2(new_n593), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n665), .A2(new_n666), .ZN(new_n971));
  AND4_X1   g785(.A1(new_n970), .A2(new_n944), .A3(new_n971), .A4(new_n961), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n970), .B1(new_n957), .B2(new_n971), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n960), .A2(new_n974), .ZN(new_n975));
  OAI221_X1 g789(.A(new_n969), .B1(new_n954), .B2(KEYINPUT61), .C1(new_n972), .C2(new_n973), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n481), .B2(new_n501), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n888), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n916), .B1(G898), .B2(new_n326), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  NAND2_X1  g795(.A1(new_n278), .A2(new_n280), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(new_n433), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n323), .A2(new_n596), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n786), .A2(new_n843), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n693), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n866), .A2(new_n713), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n703), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n991), .A2(new_n810), .A3(new_n820), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n983), .B1(new_n992), .B2(G953), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n983), .B1(G900), .B2(G953), .ZN(new_n994));
  INV_X1    g808(.A(new_n770), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n866), .A2(new_n713), .A3(new_n772), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n984), .A2(new_n604), .A3(new_n690), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n995), .B(new_n996), .C1(new_n808), .C2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n810), .A2(new_n820), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n994), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n993), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n326), .B1(G227), .B2(G900), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1002), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n993), .A2(new_n1004), .A3(new_n1000), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(G72));
  INV_X1    g820(.A(new_n698), .ZN(new_n1007));
  XOR2_X1   g821(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n697), .A2(new_n266), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT127), .Z(new_n1013));
  OAI211_X1 g827(.A(new_n872), .B(new_n1013), .C1(new_n877), .C2(new_n878), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n810), .A2(new_n998), .A3(new_n820), .A4(new_n888), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1015), .A2(new_n1010), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n936), .B(new_n1014), .C1(new_n1016), .C2(new_n1011), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n991), .A2(new_n810), .A3(new_n820), .A4(new_n888), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1007), .B1(new_n1018), .B2(new_n1010), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1017), .B1(new_n1021), .B2(new_n1022), .ZN(G57));
endmodule


