

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791;

  XNOR2_X1 U380 ( .A(n525), .B(n524), .ZN(n668) );
  XNOR2_X1 U381 ( .A(n451), .B(G107), .ZN(n769) );
  INV_X1 U382 ( .A(G237), .ZN(n456) );
  NAND2_X2 U383 ( .A1(n562), .A2(n611), .ZN(n393) );
  XNOR2_X1 U384 ( .A(n359), .B(n605), .ZN(n610) );
  NAND2_X1 U385 ( .A1(n604), .A2(n640), .ZN(n359) );
  OR2_X1 U386 ( .A1(n453), .A2(n506), .ZN(n455) );
  XNOR2_X2 U387 ( .A(n653), .B(n655), .ZN(n656) );
  XNOR2_X2 U388 ( .A(n668), .B(KEYINPUT62), .ZN(n669) );
  AND2_X2 U389 ( .A1(n626), .A2(n736), .ZN(n627) );
  INV_X1 U390 ( .A(KEYINPUT68), .ZN(n387) );
  NOR2_X1 U391 ( .A1(G953), .A2(G237), .ZN(n517) );
  INV_X2 U392 ( .A(G953), .ZN(n379) );
  AND2_X2 U393 ( .A1(n426), .A2(n421), .ZN(n366) );
  NAND2_X2 U394 ( .A1(n367), .A2(n435), .ZN(n371) );
  XNOR2_X2 U395 ( .A(n515), .B(KEYINPUT73), .ZN(n452) );
  XNOR2_X2 U396 ( .A(n452), .B(n769), .ZN(n506) );
  NAND2_X2 U397 ( .A1(G234), .A2(G237), .ZN(n461) );
  XNOR2_X1 U398 ( .A(n360), .B(KEYINPUT87), .ZN(n416) );
  NOR2_X1 U399 ( .A1(n789), .A2(n790), .ZN(n413) );
  XNOR2_X1 U400 ( .A(n364), .B(n363), .ZN(n789) );
  NOR2_X1 U401 ( .A1(n595), .A2(n721), .ZN(n607) );
  NOR2_X1 U402 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U403 ( .A(n629), .ZN(n363) );
  XNOR2_X1 U404 ( .A(n418), .B(KEYINPUT93), .ZN(n442) );
  INV_X2 U405 ( .A(KEYINPUT64), .ZN(n445) );
  XNOR2_X2 U406 ( .A(KEYINPUT71), .B(G140), .ZN(n532) );
  XNOR2_X2 U407 ( .A(KEYINPUT8), .B(KEYINPUT69), .ZN(n381) );
  NAND2_X1 U408 ( .A1(n361), .A2(n791), .ZN(n360) );
  XNOR2_X1 U409 ( .A(n362), .B(n392), .ZN(n361) );
  NAND2_X1 U410 ( .A1(n409), .A2(n412), .ZN(n362) );
  NAND2_X1 U411 ( .A1(n646), .A2(n705), .ZN(n364) );
  XNOR2_X2 U412 ( .A(n365), .B(KEYINPUT39), .ZN(n646) );
  NAND2_X1 U413 ( .A1(n627), .A2(n628), .ZN(n365) );
  NAND2_X1 U414 ( .A1(n366), .A2(n419), .ZN(n367) );
  BUF_X1 U415 ( .A(n407), .Z(n368) );
  AND2_X2 U416 ( .A1(n416), .A2(n711), .ZN(n785) );
  BUF_X1 U417 ( .A(n686), .Z(n369) );
  XNOR2_X1 U418 ( .A(n780), .B(n511), .ZN(n686) );
  OR2_X1 U419 ( .A1(n621), .A2(n742), .ZN(n370) );
  OR2_X2 U420 ( .A1(n621), .A2(n742), .ZN(n635) );
  XNOR2_X1 U421 ( .A(n393), .B(n563), .ZN(n372) );
  NAND2_X1 U422 ( .A1(n367), .A2(n435), .ZN(n434) );
  XNOR2_X1 U423 ( .A(n393), .B(n563), .ZN(n674) );
  XNOR2_X2 U424 ( .A(n623), .B(n622), .ZN(n752) );
  AND2_X2 U425 ( .A1(n635), .A2(n395), .ZN(n402) );
  NOR2_X2 U426 ( .A1(n374), .A2(n624), .ZN(n703) );
  NOR2_X1 U427 ( .A1(n403), .A2(n397), .ZN(n396) );
  NAND2_X1 U428 ( .A1(n468), .A2(KEYINPUT0), .ZN(n403) );
  NOR2_X1 U429 ( .A1(n411), .A2(n410), .ZN(n409) );
  XNOR2_X1 U430 ( .A(KEYINPUT4), .B(G137), .ZN(n518) );
  INV_X1 U431 ( .A(KEYINPUT92), .ZN(n436) );
  INV_X1 U432 ( .A(KEYINPUT38), .ZN(n383) );
  AND2_X1 U433 ( .A1(n404), .A2(n469), .ZN(n399) );
  XNOR2_X1 U434 ( .A(KEYINPUT30), .B(KEYINPUT107), .ZN(n605) );
  XNOR2_X1 U435 ( .A(n479), .B(n478), .ZN(n662) );
  XOR2_X1 U436 ( .A(G146), .B(KEYINPUT79), .Z(n504) );
  NAND2_X1 U437 ( .A1(n715), .A2(n428), .ZN(n435) );
  XNOR2_X1 U438 ( .A(n417), .B(n429), .ZN(n428) );
  INV_X1 U439 ( .A(KEYINPUT86), .ZN(n429) );
  NAND2_X1 U440 ( .A1(n433), .A2(n615), .ZN(n410) );
  INV_X1 U441 ( .A(n406), .ZN(n397) );
  INV_X1 U442 ( .A(n649), .ZN(n425) );
  NOR2_X1 U443 ( .A1(n403), .A2(n460), .ZN(n395) );
  NOR2_X1 U444 ( .A1(G953), .A2(n750), .ZN(n466) );
  XNOR2_X1 U445 ( .A(n382), .B(n381), .ZN(n529) );
  AND2_X1 U446 ( .A1(n650), .A2(n716), .ZN(n427) );
  NAND2_X1 U447 ( .A1(n424), .A2(n422), .ZN(n421) );
  NAND2_X1 U448 ( .A1(n649), .A2(n423), .ZN(n422) );
  NAND2_X1 U449 ( .A1(n425), .A2(KEYINPUT66), .ZN(n424) );
  NAND2_X1 U450 ( .A1(KEYINPUT66), .A2(KEYINPUT2), .ZN(n423) );
  XOR2_X1 U451 ( .A(G122), .B(KEYINPUT12), .Z(n471) );
  XNOR2_X1 U452 ( .A(G143), .B(G113), .ZN(n473) );
  XOR2_X1 U453 ( .A(G140), .B(G104), .Z(n474) );
  XNOR2_X1 U454 ( .A(G137), .B(KEYINPUT96), .ZN(n507) );
  INV_X1 U455 ( .A(KEYINPUT48), .ZN(n392) );
  BUF_X1 U456 ( .A(n558), .Z(n565) );
  NOR2_X1 U457 ( .A1(n742), .A2(KEYINPUT19), .ZN(n406) );
  INV_X1 U458 ( .A(G902), .ZN(n526) );
  XNOR2_X1 U459 ( .A(KEYINPUT16), .B(G122), .ZN(n439) );
  XNOR2_X1 U460 ( .A(KEYINPUT97), .B(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U461 ( .A(G137), .B(KEYINPUT78), .ZN(n537) );
  XOR2_X1 U462 ( .A(KEYINPUT9), .B(G122), .Z(n486) );
  XNOR2_X1 U463 ( .A(G116), .B(G107), .ZN(n485) );
  XNOR2_X1 U464 ( .A(n380), .B(n484), .ZN(n488) );
  XOR2_X1 U465 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n484) );
  NAND2_X1 U466 ( .A1(n529), .A2(G217), .ZN(n380) );
  INV_X1 U467 ( .A(KEYINPUT41), .ZN(n622) );
  XNOR2_X1 U468 ( .A(n502), .B(n501), .ZN(n550) );
  XNOR2_X1 U469 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n501) );
  NAND2_X1 U470 ( .A1(n558), .A2(n500), .ZN(n502) );
  AND2_X1 U471 ( .A1(n610), .A2(n609), .ZN(n628) );
  NAND2_X1 U472 ( .A1(n407), .A2(n406), .ZN(n404) );
  NAND2_X1 U473 ( .A1(n370), .A2(KEYINPUT19), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n624) );
  INV_X1 U475 ( .A(KEYINPUT109), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n483), .B(n482), .ZN(n574) );
  AND2_X1 U477 ( .A1(n378), .A2(G953), .ZN(n774) );
  INV_X1 U478 ( .A(G898), .ZN(n378) );
  XNOR2_X1 U479 ( .A(n662), .B(KEYINPUT59), .ZN(n663) );
  INV_X1 U480 ( .A(n435), .ZN(n719) );
  XNOR2_X1 U481 ( .A(n625), .B(KEYINPUT42), .ZN(n790) );
  NOR2_X1 U482 ( .A1(n752), .A2(n624), .ZN(n625) );
  XNOR2_X1 U483 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n629) );
  OR2_X1 U484 ( .A1(n468), .A2(KEYINPUT0), .ZN(n373) );
  AND2_X1 U485 ( .A1(n405), .A2(n404), .ZN(n374) );
  AND2_X1 U486 ( .A1(n736), .A2(n740), .ZN(n375) );
  BUF_X1 U487 ( .A(n727), .Z(n388) );
  AND2_X1 U488 ( .A1(n711), .A2(KEYINPUT2), .ZN(n376) );
  INV_X1 U489 ( .A(KEYINPUT0), .ZN(n469) );
  AND2_X1 U490 ( .A1(n649), .A2(KEYINPUT66), .ZN(n377) );
  NAND2_X1 U491 ( .A1(n379), .A2(G224), .ZN(n440) );
  NAND2_X1 U492 ( .A1(n379), .A2(G234), .ZN(n382) );
  NAND2_X1 U493 ( .A1(n379), .A2(G227), .ZN(n503) );
  NAND2_X1 U494 ( .A1(n786), .A2(n379), .ZN(n787) );
  NAND2_X1 U495 ( .A1(n759), .A2(n379), .ZN(n760) );
  XNOR2_X2 U496 ( .A(n407), .B(n383), .ZN(n736) );
  INV_X2 U497 ( .A(n621), .ZN(n407) );
  BUF_X1 U498 ( .A(n651), .Z(n715) );
  XNOR2_X2 U499 ( .A(n371), .B(KEYINPUT65), .ZN(n384) );
  XNOR2_X1 U500 ( .A(n434), .B(KEYINPUT65), .ZN(n678) );
  BUF_X1 U501 ( .A(n568), .Z(n626) );
  AND2_X1 U502 ( .A1(n640), .A2(n740), .ZN(n385) );
  INV_X2 U503 ( .A(KEYINPUT17), .ZN(n418) );
  INV_X1 U504 ( .A(n368), .ZN(n386) );
  XNOR2_X1 U505 ( .A(n389), .B(KEYINPUT32), .ZN(n553) );
  BUF_X1 U506 ( .A(n550), .Z(n579) );
  BUF_X1 U507 ( .A(n553), .Z(n551) );
  NAND2_X1 U508 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U509 ( .A1(n549), .A2(n638), .ZN(n390) );
  XNOR2_X2 U510 ( .A(n514), .B(n510), .ZN(n780) );
  XNOR2_X2 U511 ( .A(n387), .B(G101), .ZN(n515) );
  NAND2_X1 U512 ( .A1(n550), .A2(n390), .ZN(n389) );
  NAND2_X1 U513 ( .A1(n647), .A2(n427), .ZN(n426) );
  NAND2_X1 U514 ( .A1(n785), .A2(n651), .ZN(n647) );
  XNOR2_X2 U515 ( .A(n458), .B(n457), .ZN(n621) );
  NAND2_X1 U516 ( .A1(n391), .A2(n633), .ZN(n557) );
  XNOR2_X1 U517 ( .A(n566), .B(KEYINPUT104), .ZN(n391) );
  AND2_X2 U518 ( .A1(n555), .A2(n725), .ZN(n566) );
  NAND2_X1 U519 ( .A1(n394), .A2(n373), .ZN(n401) );
  NAND2_X1 U520 ( .A1(n407), .A2(n396), .ZN(n394) );
  NAND2_X1 U521 ( .A1(n400), .A2(n398), .ZN(n558) );
  NAND2_X1 U522 ( .A1(n399), .A2(n405), .ZN(n398) );
  NOR2_X2 U523 ( .A1(n402), .A2(n401), .ZN(n400) );
  OR2_X2 U524 ( .A1(n408), .A2(G902), .ZN(n545) );
  XNOR2_X1 U525 ( .A(n675), .B(n408), .ZN(n677) );
  XNOR2_X1 U526 ( .A(n540), .B(n539), .ZN(n408) );
  NAND2_X1 U527 ( .A1(n620), .A2(n616), .ZN(n411) );
  XNOR2_X1 U528 ( .A(n413), .B(KEYINPUT46), .ZN(n412) );
  NAND2_X1 U529 ( .A1(n598), .A2(n599), .ZN(n415) );
  NAND2_X1 U530 ( .A1(n416), .A2(n376), .ZN(n417) );
  NAND2_X1 U531 ( .A1(n420), .A2(n377), .ZN(n419) );
  XNOR2_X1 U532 ( .A(n589), .B(n588), .ZN(n651) );
  INV_X1 U533 ( .A(n647), .ZN(n420) );
  NAND2_X1 U534 ( .A1(n430), .A2(n572), .ZN(n576) );
  INV_X1 U535 ( .A(n431), .ZN(n430) );
  NAND2_X1 U536 ( .A1(n431), .A2(n705), .ZN(n706) );
  NAND2_X1 U537 ( .A1(n431), .A2(n707), .ZN(n708) );
  XNOR2_X2 U538 ( .A(n567), .B(KEYINPUT31), .ZN(n431) );
  XNOR2_X2 U539 ( .A(n432), .B(G119), .ZN(n438) );
  XNOR2_X2 U540 ( .A(G116), .B(KEYINPUT3), .ZN(n432) );
  INV_X1 U541 ( .A(n709), .ZN(n433) );
  XNOR2_X2 U542 ( .A(G143), .B(G128), .ZN(n446) );
  XNOR2_X2 U543 ( .A(n445), .B(KEYINPUT82), .ZN(n447) );
  XNOR2_X2 U544 ( .A(n447), .B(n446), .ZN(n489) );
  INV_X1 U545 ( .A(KEYINPUT45), .ZN(n588) );
  XNOR2_X1 U546 ( .A(n477), .B(n778), .ZN(n478) );
  XNOR2_X1 U547 ( .A(n481), .B(n480), .ZN(n482) );
  BUF_X1 U548 ( .A(n678), .Z(n682) );
  XNOR2_X1 U549 ( .A(n436), .B(G113), .ZN(n437) );
  XNOR2_X2 U550 ( .A(n438), .B(n437), .ZN(n513) );
  XNOR2_X2 U551 ( .A(n513), .B(n439), .ZN(n770) );
  XNOR2_X2 U552 ( .A(G146), .B(G125), .ZN(n476) );
  XNOR2_X1 U553 ( .A(n476), .B(n440), .ZN(n444) );
  XNOR2_X1 U554 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n441) );
  XNOR2_X1 U555 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U556 ( .A(n443), .B(n444), .ZN(n449) );
  INV_X1 U557 ( .A(n489), .ZN(n448) );
  XNOR2_X1 U558 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U559 ( .A(n770), .B(n450), .ZN(n453) );
  XNOR2_X1 U560 ( .A(G104), .B(G110), .ZN(n451) );
  NAND2_X1 U561 ( .A1(n453), .A2(n506), .ZN(n454) );
  NAND2_X1 U562 ( .A1(n455), .A2(n454), .ZN(n652) );
  XNOR2_X2 U563 ( .A(G902), .B(KEYINPUT15), .ZN(n648) );
  NAND2_X1 U564 ( .A1(n652), .A2(n648), .ZN(n458) );
  NAND2_X1 U565 ( .A1(n526), .A2(n456), .ZN(n459) );
  NAND2_X1 U566 ( .A1(n459), .A2(G210), .ZN(n457) );
  NAND2_X1 U567 ( .A1(n459), .A2(G214), .ZN(n640) );
  INV_X1 U568 ( .A(n640), .ZN(n742) );
  INV_X1 U569 ( .A(KEYINPUT19), .ZN(n460) );
  XNOR2_X1 U570 ( .A(n461), .B(KEYINPUT14), .ZN(n462) );
  XNOR2_X1 U571 ( .A(KEYINPUT76), .B(n462), .ZN(n464) );
  NAND2_X1 U572 ( .A1(n464), .A2(G902), .ZN(n463) );
  XNOR2_X1 U573 ( .A(n463), .B(KEYINPUT95), .ZN(n590) );
  NAND2_X1 U574 ( .A1(n590), .A2(n774), .ZN(n467) );
  NAND2_X1 U575 ( .A1(G952), .A2(n464), .ZN(n750) );
  INV_X1 U576 ( .A(KEYINPUT94), .ZN(n465) );
  XNOR2_X1 U577 ( .A(n466), .B(n465), .ZN(n592) );
  NAND2_X1 U578 ( .A1(n467), .A2(n592), .ZN(n468) );
  NAND2_X1 U579 ( .A1(G214), .A2(n517), .ZN(n470) );
  XNOR2_X1 U580 ( .A(n471), .B(n470), .ZN(n472) );
  XOR2_X1 U581 ( .A(n472), .B(KEYINPUT11), .Z(n479) );
  XNOR2_X1 U582 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X2 U583 ( .A(KEYINPUT70), .B(G131), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n475), .B(n520), .ZN(n477) );
  XNOR2_X1 U585 ( .A(n476), .B(KEYINPUT10), .ZN(n778) );
  NOR2_X1 U586 ( .A1(G902), .A2(n662), .ZN(n483) );
  XNOR2_X1 U587 ( .A(KEYINPUT13), .B(KEYINPUT100), .ZN(n481) );
  INV_X1 U588 ( .A(G475), .ZN(n480) );
  XNOR2_X1 U589 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n488), .B(n487), .ZN(n491) );
  XNOR2_X2 U591 ( .A(n489), .B(G134), .ZN(n514) );
  INV_X1 U592 ( .A(n514), .ZN(n490) );
  XNOR2_X1 U593 ( .A(n491), .B(n490), .ZN(n679) );
  NAND2_X1 U594 ( .A1(n679), .A2(n526), .ZN(n493) );
  XNOR2_X1 U595 ( .A(KEYINPUT102), .B(G478), .ZN(n492) );
  XNOR2_X1 U596 ( .A(n493), .B(n492), .ZN(n573) );
  INV_X1 U597 ( .A(n573), .ZN(n561) );
  NAND2_X1 U598 ( .A1(n574), .A2(n561), .ZN(n494) );
  XNOR2_X2 U599 ( .A(n494), .B(KEYINPUT103), .ZN(n740) );
  XOR2_X1 U600 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n498) );
  NAND2_X1 U601 ( .A1(G234), .A2(n648), .ZN(n495) );
  XNOR2_X1 U602 ( .A(KEYINPUT20), .B(n495), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n541), .A2(G221), .ZN(n496) );
  XNOR2_X1 U604 ( .A(KEYINPUT98), .B(n496), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n498), .B(n497), .ZN(n721) );
  INV_X1 U606 ( .A(n721), .ZN(n499) );
  AND2_X1 U607 ( .A1(n740), .A2(n499), .ZN(n500) );
  XNOR2_X1 U608 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n506), .B(n505), .ZN(n511) );
  XNOR2_X1 U610 ( .A(n520), .B(n532), .ZN(n509) );
  XNOR2_X1 U611 ( .A(n507), .B(KEYINPUT4), .ZN(n508) );
  XNOR2_X1 U612 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U613 ( .A1(n686), .A2(n526), .ZN(n512) );
  XNOR2_X2 U614 ( .A(n512), .B(G469), .ZN(n568) );
  XNOR2_X1 U615 ( .A(n568), .B(KEYINPUT1), .ZN(n555) );
  BUF_X1 U616 ( .A(n555), .Z(n724) );
  XNOR2_X1 U617 ( .A(n513), .B(n514), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n515), .B(G146), .ZN(n516) );
  XNOR2_X1 U619 ( .A(n516), .B(KEYINPUT5), .ZN(n523) );
  NAND2_X1 U620 ( .A1(n517), .A2(G210), .ZN(n519) );
  XNOR2_X1 U621 ( .A(n519), .B(n518), .ZN(n521) );
  XNOR2_X1 U622 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U623 ( .A(n523), .B(n522), .ZN(n524) );
  NAND2_X1 U624 ( .A1(n668), .A2(n526), .ZN(n528) );
  INV_X1 U625 ( .A(G472), .ZN(n527) );
  XNOR2_X2 U626 ( .A(n528), .B(n527), .ZN(n727) );
  NAND2_X1 U627 ( .A1(n529), .A2(G221), .ZN(n535) );
  XNOR2_X1 U628 ( .A(G119), .B(G128), .ZN(n531) );
  XNOR2_X1 U629 ( .A(KEYINPUT24), .B(G110), .ZN(n530) );
  XNOR2_X1 U630 ( .A(n531), .B(n530), .ZN(n533) );
  XNOR2_X1 U631 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U632 ( .A(n535), .B(n534), .ZN(n540) );
  XNOR2_X1 U633 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U634 ( .A(n778), .B(n538), .ZN(n539) );
  AND2_X1 U635 ( .A1(n541), .A2(G217), .ZN(n543) );
  XNOR2_X1 U636 ( .A(KEYINPUT77), .B(KEYINPUT25), .ZN(n542) );
  XNOR2_X1 U637 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X2 U638 ( .A(n545), .B(n544), .ZN(n722) );
  NAND2_X1 U639 ( .A1(n388), .A2(n722), .ZN(n546) );
  NOR2_X1 U640 ( .A1(n724), .A2(n546), .ZN(n547) );
  NAND2_X1 U641 ( .A1(n579), .A2(n547), .ZN(n552) );
  XNOR2_X1 U642 ( .A(n552), .B(G110), .ZN(G12) );
  INV_X1 U643 ( .A(n724), .ZN(n638) );
  XNOR2_X1 U644 ( .A(n727), .B(KEYINPUT6), .ZN(n633) );
  XNOR2_X1 U645 ( .A(n633), .B(KEYINPUT81), .ZN(n548) );
  NAND2_X1 U646 ( .A1(n548), .A2(n722), .ZN(n549) );
  XNOR2_X1 U647 ( .A(n551), .B(G119), .ZN(G21) );
  XNOR2_X1 U648 ( .A(n554), .B(KEYINPUT89), .ZN(n564) );
  NOR2_X1 U649 ( .A1(n722), .A2(n721), .ZN(n725) );
  XNOR2_X1 U650 ( .A(KEYINPUT74), .B(KEYINPUT33), .ZN(n556) );
  XNOR2_X2 U651 ( .A(n557), .B(n556), .ZN(n751) );
  NAND2_X1 U652 ( .A1(n751), .A2(n565), .ZN(n560) );
  XNOR2_X1 U653 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n559) );
  XNOR2_X1 U654 ( .A(n560), .B(n559), .ZN(n562) );
  NOR2_X1 U655 ( .A1(n574), .A2(n561), .ZN(n611) );
  XOR2_X1 U656 ( .A(KEYINPUT80), .B(KEYINPUT35), .Z(n563) );
  NAND2_X1 U657 ( .A1(n564), .A2(n674), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n584), .A2(KEYINPUT44), .ZN(n582) );
  INV_X1 U659 ( .A(n565), .ZN(n571) );
  NAND2_X1 U660 ( .A1(n566), .A2(n604), .ZN(n732) );
  OR2_X2 U661 ( .A1(n571), .A2(n732), .ZN(n567) );
  AND2_X1 U662 ( .A1(n725), .A2(n388), .ZN(n569) );
  NAND2_X1 U663 ( .A1(n626), .A2(n569), .ZN(n570) );
  OR2_X1 U664 ( .A1(n571), .A2(n570), .ZN(n572) );
  INV_X1 U665 ( .A(n572), .ZN(n696) );
  OR2_X1 U666 ( .A1(n574), .A2(n573), .ZN(n631) );
  INV_X1 U667 ( .A(n631), .ZN(n705) );
  AND2_X1 U668 ( .A1(n574), .A2(n573), .ZN(n707) );
  NOR2_X1 U669 ( .A1(n705), .A2(n707), .ZN(n737) );
  XNOR2_X1 U670 ( .A(KEYINPUT83), .B(n737), .ZN(n575) );
  AND2_X1 U671 ( .A1(n576), .A2(n575), .ZN(n580) );
  OR2_X1 U672 ( .A1(n633), .A2(n722), .ZN(n577) );
  NOR2_X1 U673 ( .A1(n724), .A2(n577), .ZN(n578) );
  AND2_X1 U674 ( .A1(n579), .A2(n578), .ZN(n691) );
  NOR2_X2 U675 ( .A1(n580), .A2(n691), .ZN(n581) );
  NAND2_X1 U676 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U677 ( .A(n583), .B(KEYINPUT88), .ZN(n587) );
  BUF_X1 U678 ( .A(n584), .Z(n585) );
  NOR2_X1 U679 ( .A1(n585), .A2(KEYINPUT44), .ZN(n586) );
  NOR2_X2 U680 ( .A1(n587), .A2(n586), .ZN(n589) );
  XNOR2_X1 U681 ( .A(n626), .B(KEYINPUT108), .ZN(n599) );
  NAND2_X1 U682 ( .A1(G953), .A2(n590), .ZN(n591) );
  NOR2_X1 U683 ( .A1(G900), .A2(n591), .ZN(n594) );
  INV_X1 U684 ( .A(n592), .ZN(n593) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT72), .ZN(n596) );
  NAND2_X1 U686 ( .A1(n596), .A2(n722), .ZN(n630) );
  NOR2_X1 U687 ( .A1(n630), .A2(n727), .ZN(n597) );
  XNOR2_X1 U688 ( .A(n597), .B(KEYINPUT28), .ZN(n598) );
  NOR2_X1 U689 ( .A1(KEYINPUT83), .A2(n737), .ZN(n600) );
  NAND2_X1 U690 ( .A1(n703), .A2(n600), .ZN(n601) );
  INV_X1 U691 ( .A(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n601), .A2(n617), .ZN(n603) );
  NAND2_X1 U693 ( .A1(n703), .A2(KEYINPUT47), .ZN(n602) );
  NAND2_X1 U694 ( .A1(n603), .A2(n602), .ZN(n616) );
  INV_X1 U695 ( .A(n727), .ZN(n604) );
  INV_X1 U696 ( .A(n607), .ZN(n608) );
  NOR2_X1 U697 ( .A1(n722), .A2(n608), .ZN(n609) );
  AND2_X1 U698 ( .A1(n628), .A2(n626), .ZN(n614) );
  INV_X1 U699 ( .A(n611), .ZN(n612) );
  NOR2_X1 U700 ( .A1(n612), .A2(n386), .ZN(n613) );
  NAND2_X1 U701 ( .A1(n614), .A2(n613), .ZN(n702) );
  XNOR2_X1 U702 ( .A(KEYINPUT84), .B(n702), .ZN(n615) );
  NAND2_X1 U703 ( .A1(n703), .A2(KEYINPUT83), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U705 ( .A1(n619), .A2(n737), .ZN(n620) );
  NAND2_X1 U706 ( .A1(n385), .A2(n736), .ZN(n623) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U709 ( .A(n634), .B(KEYINPUT105), .ZN(n641) );
  INV_X1 U710 ( .A(n370), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n641), .A2(n636), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n637), .B(KEYINPUT36), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n709) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U715 ( .A1(n642), .A2(n724), .ZN(n643) );
  XOR2_X1 U716 ( .A(KEYINPUT43), .B(n643), .Z(n644) );
  NAND2_X1 U717 ( .A1(n644), .A2(n386), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n645), .B(KEYINPUT106), .ZN(n791) );
  NAND2_X1 U719 ( .A1(n646), .A2(n707), .ZN(n711) );
  INV_X1 U720 ( .A(KEYINPUT2), .ZN(n716) );
  INV_X1 U721 ( .A(n648), .ZN(n649) );
  INV_X1 U722 ( .A(KEYINPUT66), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n384), .A2(G210), .ZN(n657) );
  BUF_X1 U724 ( .A(n652), .Z(n653) );
  XNOR2_X1 U725 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n654) );
  XOR2_X1 U726 ( .A(n654), .B(KEYINPUT90), .Z(n655) );
  XNOR2_X1 U727 ( .A(n657), .B(n656), .ZN(n659) );
  INV_X1 U728 ( .A(G952), .ZN(n658) );
  NAND2_X1 U729 ( .A1(n658), .A2(G953), .ZN(n676) );
  NAND2_X1 U730 ( .A1(n659), .A2(n676), .ZN(n661) );
  XNOR2_X1 U731 ( .A(KEYINPUT119), .B(KEYINPUT56), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n661), .B(n660), .ZN(G51) );
  NAND2_X1 U733 ( .A1(n678), .A2(G475), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n665), .A2(n676), .ZN(n667) );
  INV_X1 U736 ( .A(KEYINPUT60), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n667), .B(n666), .ZN(G60) );
  NAND2_X1 U738 ( .A1(n384), .A2(G472), .ZN(n670) );
  XNOR2_X1 U739 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U740 ( .A1(n671), .A2(n676), .ZN(n673) );
  XOR2_X1 U741 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(G57) );
  XNOR2_X1 U743 ( .A(n372), .B(G122), .ZN(G24) );
  NAND2_X1 U744 ( .A1(n682), .A2(G217), .ZN(n675) );
  INV_X1 U745 ( .A(n676), .ZN(n689) );
  NOR2_X1 U746 ( .A1(n677), .A2(n689), .ZN(G66) );
  NAND2_X1 U747 ( .A1(n384), .A2(G478), .ZN(n680) );
  XOR2_X1 U748 ( .A(n680), .B(n679), .Z(n681) );
  NOR2_X1 U749 ( .A1(n681), .A2(n689), .ZN(G63) );
  NAND2_X1 U750 ( .A1(n682), .A2(G469), .ZN(n688) );
  XOR2_X1 U751 ( .A(KEYINPUT121), .B(KEYINPUT57), .Z(n684) );
  XNOR2_X1 U752 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U754 ( .A(n369), .B(n685), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n690), .A2(n689), .ZN(G54) );
  XOR2_X1 U757 ( .A(G101), .B(n691), .Z(G3) );
  NAND2_X1 U758 ( .A1(n696), .A2(n705), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(G104), .ZN(G6) );
  XOR2_X1 U760 ( .A(KEYINPUT112), .B(KEYINPUT27), .Z(n694) );
  XNOR2_X1 U761 ( .A(G107), .B(KEYINPUT26), .ZN(n693) );
  XNOR2_X1 U762 ( .A(n694), .B(n693), .ZN(n695) );
  XOR2_X1 U763 ( .A(KEYINPUT111), .B(n695), .Z(n698) );
  NAND2_X1 U764 ( .A1(n696), .A2(n707), .ZN(n697) );
  XNOR2_X1 U765 ( .A(n698), .B(n697), .ZN(G9) );
  XOR2_X1 U766 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n700) );
  NAND2_X1 U767 ( .A1(n703), .A2(n707), .ZN(n699) );
  XNOR2_X1 U768 ( .A(n700), .B(n699), .ZN(n701) );
  XOR2_X1 U769 ( .A(G128), .B(n701), .Z(G30) );
  XNOR2_X1 U770 ( .A(G143), .B(n702), .ZN(G45) );
  NAND2_X1 U771 ( .A1(n703), .A2(n705), .ZN(n704) );
  XNOR2_X1 U772 ( .A(n704), .B(G146), .ZN(G48) );
  XNOR2_X1 U773 ( .A(n706), .B(G113), .ZN(G15) );
  XNOR2_X1 U774 ( .A(n708), .B(G116), .ZN(G18) );
  XNOR2_X1 U775 ( .A(n709), .B(G125), .ZN(n710) );
  XNOR2_X1 U776 ( .A(n710), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U777 ( .A(G134), .B(KEYINPUT114), .ZN(n712) );
  XNOR2_X1 U778 ( .A(n712), .B(n711), .ZN(G36) );
  XOR2_X1 U779 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n761) );
  BUF_X1 U780 ( .A(n785), .Z(n713) );
  NOR2_X1 U781 ( .A1(n713), .A2(KEYINPUT2), .ZN(n714) );
  XNOR2_X1 U782 ( .A(n714), .B(KEYINPUT85), .ZN(n718) );
  INV_X1 U783 ( .A(n715), .ZN(n762) );
  NAND2_X1 U784 ( .A1(n762), .A2(n716), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n720) );
  NOR2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n758) );
  XNOR2_X1 U787 ( .A(KEYINPUT51), .B(KEYINPUT115), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U789 ( .A(n723), .B(KEYINPUT49), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U791 ( .A(KEYINPUT50), .B(n726), .Z(n728) );
  NAND2_X1 U792 ( .A1(n728), .A2(n388), .ZN(n729) );
  OR2_X1 U793 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U794 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U795 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U796 ( .A1(n735), .A2(n752), .ZN(n746) );
  INV_X1 U797 ( .A(n736), .ZN(n738) );
  NOR2_X1 U798 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U799 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U800 ( .A1(n742), .A2(n741), .ZN(n743) );
  OR2_X1 U801 ( .A1(n743), .A2(n375), .ZN(n744) );
  AND2_X1 U802 ( .A1(n751), .A2(n744), .ZN(n745) );
  NOR2_X1 U803 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U804 ( .A(n747), .B(KEYINPUT116), .ZN(n748) );
  XNOR2_X1 U805 ( .A(KEYINPUT52), .B(n748), .ZN(n749) );
  NOR2_X1 U806 ( .A1(n750), .A2(n749), .ZN(n755) );
  INV_X1 U807 ( .A(n751), .ZN(n753) );
  NOR2_X1 U808 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U809 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U810 ( .A(n756), .B(KEYINPUT117), .ZN(n757) );
  NOR2_X1 U811 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U812 ( .A(n761), .B(n760), .ZN(G75) );
  NOR2_X1 U813 ( .A1(n762), .A2(G953), .ZN(n763) );
  XNOR2_X1 U814 ( .A(n763), .B(KEYINPUT123), .ZN(n768) );
  NAND2_X1 U815 ( .A1(G953), .A2(G224), .ZN(n764) );
  XNOR2_X1 U816 ( .A(KEYINPUT61), .B(n764), .ZN(n765) );
  NAND2_X1 U817 ( .A1(n765), .A2(G898), .ZN(n766) );
  XNOR2_X1 U818 ( .A(KEYINPUT122), .B(n766), .ZN(n767) );
  NAND2_X1 U819 ( .A1(n768), .A2(n767), .ZN(n776) );
  XOR2_X1 U820 ( .A(n769), .B(KEYINPUT124), .Z(n771) );
  XNOR2_X1 U821 ( .A(n770), .B(n771), .ZN(n772) );
  XNOR2_X1 U822 ( .A(n772), .B(G101), .ZN(n773) );
  NOR2_X1 U823 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U824 ( .A(n776), .B(n775), .ZN(n777) );
  XOR2_X1 U825 ( .A(KEYINPUT125), .B(n777), .Z(G69) );
  XNOR2_X1 U826 ( .A(n778), .B(KEYINPUT126), .ZN(n779) );
  XNOR2_X1 U827 ( .A(n780), .B(n779), .ZN(n784) );
  XNOR2_X1 U828 ( .A(n784), .B(KEYINPUT127), .ZN(n781) );
  XNOR2_X1 U829 ( .A(G227), .B(n781), .ZN(n782) );
  NAND2_X1 U830 ( .A1(G900), .A2(n782), .ZN(n783) );
  NAND2_X1 U831 ( .A1(n783), .A2(G953), .ZN(n788) );
  XNOR2_X1 U832 ( .A(n713), .B(n784), .ZN(n786) );
  NAND2_X1 U833 ( .A1(n788), .A2(n787), .ZN(G72) );
  XOR2_X1 U834 ( .A(n789), .B(G131), .Z(G33) );
  XOR2_X1 U835 ( .A(n790), .B(G137), .Z(G39) );
  XNOR2_X1 U836 ( .A(G140), .B(n791), .ZN(G42) );
endmodule

