//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n461), .B2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(new_n464), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n462), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n467), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n461), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n470), .A2(new_n474), .A3(new_n477), .ZN(G160));
  NAND4_X1  g053(.A1(new_n462), .A2(new_n465), .A3(G2105), .A4(new_n467), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n466), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI22_X1  g057(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n468), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G136), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n465), .A3(new_n467), .A4(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n486), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(G114), .B2(new_n466), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n479), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n491), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  INV_X1    g073(.A(G62), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT67), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT5), .A3(G543), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n499), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT69), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n508), .B(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n506), .B2(new_n505), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n498), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n502), .A2(new_n504), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n512), .A2(new_n519), .ZN(G166));
  INV_X1    g095(.A(new_n515), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(new_n517), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT70), .B(G51), .Z(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g103(.A1(new_n522), .A2(new_n523), .A3(new_n525), .A4(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n498), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n515), .A2(new_n533), .B1(new_n517), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(G171));
  AOI22_X1  g111(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n498), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  INV_X1    g114(.A(G43), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n515), .A2(new_n539), .B1(new_n517), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  XOR2_X1   g122(.A(KEYINPUT71), .B(KEYINPUT9), .Z(new_n548));
  NAND3_X1  g123(.A1(new_n526), .A2(G53), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G53), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT71), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n517), .A2(new_n550), .B1(new_n551), .B2(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n513), .A2(KEYINPUT73), .A3(new_n514), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT73), .B1(new_n513), .B2(new_n514), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G91), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n498), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n549), .A2(KEYINPUT72), .A3(new_n552), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n555), .A2(new_n559), .A3(new_n561), .A4(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  OR2_X1    g139(.A1(new_n512), .A2(new_n519), .ZN(G303));
  OAI21_X1  g140(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT74), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n568), .B(G651), .C1(new_n513), .C2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n515), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n513), .A2(KEYINPUT73), .A3(new_n514), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n572), .A2(G87), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n526), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n558), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(new_n513), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(G48), .B2(new_n526), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(G305));
  XNOR2_X1  g158(.A(KEYINPUT75), .B(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n521), .A2(G85), .B1(new_n526), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n498), .B2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n579), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n517), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n572), .A2(new_n573), .ZN(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n558), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n588), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  INV_X1    g183(.A(new_n600), .ZN(new_n609));
  OAI21_X1  g184(.A(G868), .B1(new_n609), .B2(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n489), .A2(new_n475), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  XOR2_X1   g190(.A(KEYINPUT76), .B(KEYINPUT13), .Z(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n619));
  INV_X1    g194(.A(G123), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n479), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n484), .B2(G135), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(G2096), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n617), .A2(new_n624), .A3(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  INV_X1    g204(.A(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT79), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(new_n635), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n638), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n645), .B1(new_n638), .B2(new_n641), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n628), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n640), .B1(new_n639), .B2(new_n635), .ZN(new_n650));
  AND4_X1   g225(.A1(new_n640), .A2(new_n635), .A3(KEYINPUT14), .A4(new_n636), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n644), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n638), .A2(new_n641), .A3(new_n645), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(new_n627), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n648), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n649), .ZN(new_n657));
  INV_X1    g232(.A(new_n654), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n627), .B1(new_n652), .B2(new_n653), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n657), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n648), .A2(new_n654), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(KEYINPUT80), .A3(new_n657), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n656), .B1(new_n662), .B2(new_n664), .ZN(G401));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  OR3_X1    g244(.A1(new_n668), .A2(KEYINPUT81), .A3(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(KEYINPUT81), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  INV_X1    g246(.A(new_n666), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n667), .B(KEYINPUT17), .Z(new_n673));
  OAI211_X1 g248(.A(new_n670), .B(new_n671), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n669), .A2(new_n666), .A3(new_n667), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT18), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n669), .A3(new_n672), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2096), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT83), .Z(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n683), .A2(new_n684), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(KEYINPUT82), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT20), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n696), .B1(new_n693), .B2(new_n695), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n682), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(new_n682), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(new_n702), .A3(new_n697), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1981), .B(G1986), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n700), .A2(new_n703), .A3(new_n705), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(G229));
  MUX2_X1   g285(.A(G6), .B(G305), .S(G16), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT32), .B(G1981), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G22), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G166), .B2(G16), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(G1971), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(G1971), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n719));
  NAND2_X1  g294(.A1(G288), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT89), .A4(new_n575), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G16), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G16), .B2(G23), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n724), .A2(new_n726), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n718), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT84), .B(G29), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G25), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT85), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n484), .A2(G131), .ZN(new_n735));
  INV_X1    g310(.A(G119), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n466), .A2(G107), .ZN(new_n737));
  OAI21_X1  g312(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n479), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n735), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n734), .B1(new_n740), .B2(new_n732), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT35), .B(G1991), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT86), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n741), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT87), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(KEYINPUT87), .ZN(new_n747));
  INV_X1    g322(.A(G16), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G24), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT88), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G290), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(G1986), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n731), .A2(new_n746), .A3(new_n747), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n729), .A2(new_n730), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(new_n732), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(G35), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G162), .B2(new_n758), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT29), .B(G2090), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n763), .A2(G34), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n763), .A2(G34), .ZN(new_n765));
  NOR3_X1   g340(.A1(new_n758), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G160), .B2(G29), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G2084), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(KEYINPUT96), .ZN(new_n769));
  NOR2_X1   g344(.A1(G171), .A2(new_n748), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G5), .B2(new_n748), .ZN(new_n771));
  INV_X1    g346(.A(G1961), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT31), .B(G11), .Z(new_n774));
  INV_X1    g349(.A(G28), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(KEYINPUT30), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(KEYINPUT30), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n774), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n773), .B(new_n778), .C1(new_n623), .C2(new_n732), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n769), .B(new_n779), .C1(KEYINPUT96), .C2(new_n768), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n748), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT97), .B(G1956), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n732), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT92), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT28), .ZN(new_n788));
  INV_X1    g363(.A(G29), .ZN(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n791));
  INV_X1    g366(.A(G128), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n479), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n484), .B2(G140), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n788), .B1(new_n789), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2067), .ZN(new_n796));
  INV_X1    g371(.A(G139), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n468), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT93), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n489), .A2(G127), .ZN(new_n801));
  INV_X1    g376(.A(G115), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n461), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n804));
  NAND2_X1  g379(.A1(G103), .A2(G2104), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(G2105), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n466), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n803), .A2(G2105), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n809), .A2(new_n789), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n789), .B2(G33), .ZN(new_n811));
  INV_X1    g386(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n796), .B1(G2072), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n767), .A2(G2084), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n771), .B2(new_n772), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n748), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n748), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1966), .ZN(new_n818));
  INV_X1    g393(.A(G2072), .ZN(new_n819));
  AOI211_X1 g394(.A(new_n815), .B(new_n818), .C1(new_n819), .C2(new_n811), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n780), .A2(new_n785), .A3(new_n813), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n789), .A2(G32), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n823));
  AND3_X1   g398(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n824), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n825), .A2(new_n826), .B1(G105), .B2(new_n475), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n484), .A2(G141), .ZN(new_n828));
  INV_X1    g403(.A(G129), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n479), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n822), .B1(new_n831), .B2(new_n789), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT27), .B(G1996), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT95), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(G4), .A2(G16), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(new_n600), .B2(G16), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(G1348), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n760), .A2(new_n761), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n835), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G1348), .B2(new_n837), .ZN(new_n841));
  NOR2_X1   g416(.A1(G16), .A2(G19), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n542), .B2(G16), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT91), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(G1341), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n758), .A2(G27), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G164), .B2(new_n758), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(G2078), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(G1341), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n845), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n821), .A2(new_n841), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n757), .A2(new_n851), .ZN(G150));
  INV_X1    g427(.A(G150), .ZN(G311));
  AOI22_X1  g428(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n854), .A2(new_n498), .ZN(new_n855));
  INV_X1    g430(.A(G93), .ZN(new_n856));
  INV_X1    g431(.A(G55), .ZN(new_n857));
  OAI22_X1  g432(.A1(new_n515), .A2(new_n856), .B1(new_n517), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(G860), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n600), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n542), .A2(new_n859), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n538), .A2(new_n541), .B1(new_n855), .B2(new_n858), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n864), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT98), .Z(new_n871));
  OAI21_X1  g446(.A(new_n860), .B1(new_n869), .B2(KEYINPUT39), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n862), .B1(new_n871), .B2(new_n872), .ZN(G145));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n622), .B(G160), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(G162), .ZN(new_n876));
  INV_X1    g451(.A(new_n496), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n878));
  AOI221_X4 g453(.A(new_n878), .B1(new_n489), .B2(new_n490), .C1(new_n488), .C2(KEYINPUT4), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n489), .A2(new_n490), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT99), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n877), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n809), .A2(KEYINPUT100), .A3(new_n830), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n800), .A2(KEYINPUT100), .A3(new_n808), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n831), .ZN(new_n886));
  INV_X1    g461(.A(new_n794), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n884), .B2(new_n886), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n883), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n884), .A2(new_n886), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n794), .ZN(new_n893));
  INV_X1    g468(.A(new_n883), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n888), .ZN(new_n895));
  INV_X1    g470(.A(new_n740), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n466), .A2(KEYINPUT101), .A3(G118), .ZN(new_n897));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n466), .B2(G118), .ZN(new_n898));
  OR2_X1    g473(.A1(G106), .A2(G2105), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n897), .A2(G2104), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(G142), .ZN(new_n901));
  INV_X1    g476(.A(G130), .ZN(new_n902));
  OAI221_X1 g477(.A(new_n900), .B1(new_n468), .B2(new_n901), .C1(new_n902), .C2(new_n479), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT102), .ZN(new_n904));
  INV_X1    g479(.A(new_n614), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n896), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n910), .A2(new_n740), .A3(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n891), .A2(new_n895), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n891), .B2(new_n895), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n876), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n891), .A2(new_n895), .A3(new_n912), .ZN(new_n916));
  INV_X1    g491(.A(new_n876), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n916), .B(new_n917), .C1(new_n914), .C2(KEYINPUT103), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n914), .A2(KEYINPUT103), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n874), .B(new_n915), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT40), .ZN(G395));
  OR3_X1    g496(.A1(new_n600), .A2(G299), .A3(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n600), .A2(G299), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT105), .B1(new_n600), .B2(G299), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT41), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n600), .B2(G299), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n609), .A2(new_n604), .ZN(new_n928));
  AOI22_X1  g503(.A1(new_n925), .A2(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n867), .B(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n600), .A2(new_n607), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n923), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n933), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  XNOR2_X1  g513(.A(G166), .B(KEYINPUT106), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n939), .A2(new_n722), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n722), .ZN(new_n941));
  XOR2_X1   g516(.A(G305), .B(G290), .Z(new_n942));
  OR3_X1    g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n940), .B2(new_n941), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n937), .A2(new_n938), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n946), .B1(new_n937), .B2(new_n938), .ZN(new_n948));
  OAI21_X1  g523(.A(G868), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(G868), .B2(new_n859), .ZN(G295));
  OAI21_X1  g525(.A(new_n949), .B1(G868), .B2(new_n859), .ZN(G331));
  NAND3_X1  g526(.A1(new_n865), .A2(G301), .A3(new_n866), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(G301), .B1(new_n865), .B2(new_n866), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n953), .A2(new_n954), .A3(G286), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n867), .A2(G171), .ZN(new_n956));
  AOI21_X1  g531(.A(G168), .B1(new_n956), .B2(new_n952), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n934), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(G286), .B1(new_n953), .B2(new_n954), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n956), .A2(G168), .A3(new_n952), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(KEYINPUT107), .A3(new_n934), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n960), .B(new_n964), .C1(new_n929), .C2(new_n963), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n945), .ZN(new_n966));
  OR2_X1    g541(.A1(new_n966), .A2(KEYINPUT108), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n960), .A2(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n925), .A2(new_n926), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n928), .A2(new_n927), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n966), .A2(KEYINPUT108), .B1(new_n946), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT43), .B1(new_n967), .B2(new_n973), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n958), .A2(KEYINPUT110), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n958), .A2(KEYINPUT110), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n934), .A2(new_n926), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n922), .A2(new_n924), .A3(new_n927), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n963), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n975), .B(new_n976), .C1(new_n979), .C2(KEYINPUT109), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(KEYINPUT109), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n945), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n972), .A2(new_n946), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n874), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT44), .B1(new_n974), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n945), .B1(new_n968), .B2(new_n971), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(KEYINPUT108), .A3(new_n874), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n985), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n966), .A2(KEYINPUT108), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT43), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n983), .A2(new_n987), .A3(new_n874), .A4(new_n985), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n989), .B1(new_n997), .B2(KEYINPUT44), .ZN(G397));
  XOR2_X1   g573(.A(KEYINPUT111), .B(G1384), .Z(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT45), .B1(new_n883), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g576(.A(KEYINPUT112), .B(G40), .Z(new_n1002));
  NOR4_X1   g577(.A1(new_n470), .A2(new_n474), .A3(new_n477), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1996), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n830), .B(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n794), .B(G2067), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n740), .B(new_n743), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(G290), .B(G1986), .Z(new_n1012));
  AOI21_X1  g587(.A(new_n1004), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1976), .ZN(new_n1014));
  AND2_X1   g589(.A1(G288), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n1015), .B2(KEYINPUT52), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT113), .B(G8), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n880), .A2(new_n881), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n878), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n491), .A2(KEYINPUT99), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1384), .B1(new_n1021), .B2(new_n877), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1017), .B1(new_n1022), .B2(new_n1003), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n720), .A2(G1976), .A3(new_n721), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT52), .B1(G288), .B2(new_n1014), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT114), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1016), .A2(new_n1023), .A3(new_n1024), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1024), .ZN(new_n1029));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n883), .A2(new_n1030), .A3(new_n1003), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1017), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT52), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n581), .A2(G651), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n526), .A2(G48), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n521), .A2(G86), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(G1981), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n577), .A2(new_n582), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT49), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1041), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(new_n1023), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1028), .A2(new_n1034), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(G166), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n883), .A2(new_n1053), .A3(new_n1030), .ZN(new_n1054));
  INV_X1    g629(.A(G2090), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n474), .A2(new_n477), .ZN(new_n1056));
  INV_X1    g631(.A(new_n470), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1002), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1030), .B1(new_n491), .B2(new_n496), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(KEYINPUT50), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1054), .A2(new_n1055), .A3(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1059), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G1971), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(G8), .B(new_n1052), .C1(new_n1062), .C2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1047), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G288), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1046), .A2(new_n1014), .A3(new_n1069), .ZN(new_n1070));
  XOR2_X1   g645(.A(new_n1041), .B(KEYINPUT115), .Z(new_n1071));
  AOI21_X1  g646(.A(new_n1033), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1067), .A2(new_n1034), .A3(new_n1028), .A4(new_n1046), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1052), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1003), .B1(new_n1060), .B2(KEYINPUT50), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1077), .B(new_n1078), .C1(new_n1022), .C2(new_n1053), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1053), .B1(new_n883), .B2(new_n1030), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT116), .B1(new_n1080), .B2(new_n1076), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1081), .A3(new_n1055), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1066), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1032), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1074), .B1(new_n1075), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1966), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT45), .B1(new_n883), .B2(new_n1030), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1003), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(G2084), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1054), .A2(new_n1091), .A3(new_n1061), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1017), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(G168), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT63), .B1(new_n1086), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1096));
  OAI21_X1  g671(.A(G8), .B1(new_n1062), .B2(new_n1066), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1075), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1074), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1073), .B1(new_n1095), .B2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT56), .B(G2072), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1063), .A2(new_n1065), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n883), .A2(new_n1030), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1076), .B1(new_n1105), .B2(KEYINPUT50), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1106), .B2(G1956), .ZN(new_n1107));
  AND2_X1   g682(.A1(new_n559), .A2(new_n561), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n549), .B2(new_n552), .ZN(new_n1109));
  AOI22_X1  g684(.A1(G299), .A2(KEYINPUT57), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1107), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1114), .A3(new_n1111), .ZN(new_n1115));
  AOI21_X1  g690(.A(G1348), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1031), .A2(G2067), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1113), .B(new_n1115), .C1(new_n609), .C2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1110), .B(new_n1104), .C1(G1956), .C2(new_n1106), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1120), .B(KEYINPUT117), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1112), .B(KEYINPUT121), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT61), .B1(new_n1123), .B2(new_n1121), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1113), .A2(KEYINPUT61), .A3(new_n1115), .A4(new_n1120), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  NOR4_X1   g701(.A1(new_n1116), .A2(new_n1117), .A3(new_n1126), .A4(new_n600), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n609), .B1(new_n1118), .B2(KEYINPUT60), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1131), .B1(new_n1132), .B2(G1996), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1063), .A2(KEYINPUT119), .A3(new_n1065), .A4(new_n1005), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT58), .B(G1341), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1031), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1137), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n542), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n542), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1125), .A2(new_n1130), .A3(new_n1138), .A4(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1122), .B1(new_n1124), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(G286), .A2(new_n1032), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1093), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(G8), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1145), .B1(new_n1149), .B2(new_n1144), .ZN(new_n1150));
  AOI211_X1 g725(.A(G168), .B(new_n1017), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1147), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1132), .B2(G2078), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1054), .A2(new_n1061), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n772), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1001), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1154), .A2(G2078), .ZN(new_n1159));
  AND3_X1   g734(.A1(G160), .A2(G40), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1160), .A3(new_n1063), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1155), .A2(new_n1157), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(G171), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1089), .B1(new_n1105), .B2(new_n1064), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1159), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1155), .A2(new_n1157), .A3(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1163), .B(KEYINPUT54), .C1(G171), .C2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1086), .A2(new_n1153), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(G171), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1155), .A2(new_n1161), .A3(G301), .A4(new_n1157), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT54), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1168), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1102), .B1(new_n1143), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n1177));
  OR2_X1    g752(.A1(new_n1093), .A2(new_n1146), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1050), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1144), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT51), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1178), .B(KEYINPUT62), .C1(new_n1181), .C2(new_n1151), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1086), .A2(new_n1182), .A3(G171), .A4(new_n1166), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1178), .B1(new_n1181), .B2(new_n1151), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1177), .B1(new_n1183), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g763(.A(new_n1169), .B(new_n1074), .C1(new_n1075), .C2(new_n1085), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1189), .A2(KEYINPUT123), .A3(new_n1186), .A4(new_n1182), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1013), .B1(new_n1176), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT46), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1004), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1193), .B1(new_n1194), .B2(new_n1005), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1004), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1196));
  AND2_X1   g771(.A1(new_n1007), .A2(new_n831), .ZN(new_n1197));
  OAI22_X1  g772(.A1(new_n1195), .A2(new_n1196), .B1(new_n1004), .B2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT47), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n896), .A2(new_n743), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1008), .A2(new_n1200), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n887), .A2(G2067), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1004), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OR3_X1    g778(.A1(new_n1004), .A2(G1986), .A3(G290), .ZN(new_n1204));
  INV_X1    g779(.A(new_n1204), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n1205), .A2(KEYINPUT48), .ZN(new_n1206));
  AOI22_X1  g781(.A1(new_n1205), .A2(KEYINPUT48), .B1(new_n1010), .B2(new_n1194), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1203), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1199), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1209), .B1(new_n1199), .B2(new_n1208), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(KEYINPUT125), .B1(new_n1192), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1013), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1073), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1086), .A2(new_n1094), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1216), .B1(new_n1219), .B2(new_n1100), .ZN(new_n1220));
  NAND2_X1  g795(.A1(new_n1123), .A2(new_n1121), .ZN(new_n1221));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AND4_X1   g798(.A1(new_n1125), .A2(new_n1130), .A3(new_n1141), .A4(new_n1138), .ZN(new_n1224));
  AOI22_X1  g799(.A1(new_n1223), .A2(new_n1224), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1225));
  XNOR2_X1  g800(.A(new_n1171), .B(new_n1172), .ZN(new_n1226));
  AND3_X1   g801(.A1(new_n1086), .A2(new_n1153), .A3(new_n1167), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1220), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1215), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1213), .ZN(new_n1233));
  NAND3_X1  g808(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1214), .A2(new_n1234), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n1237));
  NOR2_X1   g811(.A1(G227), .A2(new_n459), .ZN(new_n1238));
  NAND3_X1  g812(.A1(new_n707), .A2(new_n708), .A3(new_n1238), .ZN(new_n1239));
  NOR3_X1   g813(.A1(G401), .A2(KEYINPUT126), .A3(new_n1239), .ZN(new_n1240));
  INV_X1    g814(.A(KEYINPUT126), .ZN(new_n1241));
  AOI21_X1  g815(.A(KEYINPUT80), .B1(new_n663), .B2(new_n657), .ZN(new_n1242));
  AOI211_X1 g816(.A(new_n661), .B(new_n649), .C1(new_n648), .C2(new_n654), .ZN(new_n1243));
  OAI211_X1 g817(.A(G14), .B(new_n655), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  INV_X1    g818(.A(new_n1239), .ZN(new_n1245));
  AOI21_X1  g819(.A(new_n1241), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g820(.A(new_n920), .B1(new_n1240), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g821(.A(new_n1247), .ZN(new_n1248));
  AOI21_X1  g822(.A(new_n1237), .B1(new_n996), .B2(new_n1248), .ZN(new_n1249));
  AOI211_X1 g823(.A(KEYINPUT127), .B(new_n1247), .C1(new_n994), .C2(new_n995), .ZN(new_n1250));
  NOR2_X1   g824(.A1(new_n1249), .A2(new_n1250), .ZN(G308));
  AOI21_X1  g825(.A(new_n987), .B1(new_n967), .B2(new_n973), .ZN(new_n1252));
  INV_X1    g826(.A(new_n995), .ZN(new_n1253));
  OAI21_X1  g827(.A(new_n1248), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g828(.A1(new_n1254), .A2(KEYINPUT127), .ZN(new_n1255));
  NAND3_X1  g829(.A1(new_n996), .A2(new_n1237), .A3(new_n1248), .ZN(new_n1256));
  NAND2_X1  g830(.A1(new_n1255), .A2(new_n1256), .ZN(G225));
endmodule


