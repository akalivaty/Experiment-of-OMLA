//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n563, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n614, new_n616, new_n617, new_n618, new_n619,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT67), .ZN(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n458), .A2(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT69), .B(G2105), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT70), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n470), .A3(new_n467), .ZN(new_n471));
  AND3_X1   g046(.A1(new_n469), .A2(G125), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n473), .B(KEYINPUT71), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n463), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n468), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  XOR2_X1   g056(.A(KEYINPUT69), .B(G2105), .Z(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n482), .C2(G112), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT72), .Z(new_n484));
  NOR2_X1   g059(.A1(new_n476), .A2(new_n482), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n476), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(G124), .A2(new_n485), .B1(new_n486), .B2(G136), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n482), .A2(G138), .A3(new_n468), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n463), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n469), .A3(new_n471), .A4(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G2105), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n498));
  OR2_X1    g073(.A1(new_n498), .A2(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(G114), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n497), .A2(G102), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n468), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n468), .A2(KEYINPUT73), .A3(new_n504), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n496), .A2(new_n509), .ZN(G164));
  OR2_X1    g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n518), .A2(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n516), .A2(new_n526), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n518), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n521), .A2(new_n520), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n517), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n515), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n544), .A2(KEYINPUT76), .A3(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n524), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n522), .A2(new_n523), .ZN(new_n548));
  INV_X1    g123(.A(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(G90), .A2(new_n547), .B1(new_n550), .B2(G52), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n546), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  AND2_X1   g128(.A1(G68), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n513), .B2(G56), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n515), .ZN(new_n556));
  INV_X1    g131(.A(G43), .ZN(new_n557));
  INV_X1    g132(.A(G81), .ZN(new_n558));
  OAI22_X1  g133(.A1(new_n518), .A2(new_n557), .B1(new_n524), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND3_X1  g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G36), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n563), .A2(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(new_n524), .A2(KEYINPUT77), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n513), .A2(new_n517), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(G91), .A3(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n517), .A2(G53), .A3(G543), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n575));
  OAI221_X1 g150(.A(new_n571), .B1(new_n515), .B2(new_n572), .C1(new_n574), .C2(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  AND2_X1   g153(.A1(new_n568), .A2(new_n570), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G87), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n513), .A2(G74), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n550), .B2(G49), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n515), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n550), .A2(G48), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n579), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(G85), .A2(new_n547), .B1(new_n550), .B2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n515), .B2(new_n591), .ZN(G290));
  INV_X1    g167(.A(G868), .ZN(new_n593));
  OR3_X1    g168(.A1(G171), .A2(KEYINPUT78), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT78), .B1(G171), .B2(new_n593), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n511), .B2(new_n512), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n550), .A2(G54), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n568), .A2(G92), .A3(new_n570), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT79), .B(KEYINPUT10), .Z(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n605), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n568), .A2(G92), .A3(new_n570), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n603), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n594), .B(new_n595), .C1(G868), .C2(new_n609), .ZN(G284));
  OAI211_X1 g185(.A(new_n594), .B(new_n595), .C1(G868), .C2(new_n609), .ZN(G321));
  MUX2_X1   g186(.A(G286), .B(G299), .S(new_n593), .Z(G297));
  MUX2_X1   g187(.A(G286), .B(G299), .S(new_n593), .Z(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n609), .B1(new_n614), .B2(G860), .ZN(G148));
  INV_X1    g190(.A(new_n560), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  INV_X1    g192(.A(new_n609), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n618), .A2(G559), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n617), .B1(new_n619), .B2(G868), .ZN(G323));
  XNOR2_X1  g195(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g196(.A1(new_n469), .A2(new_n471), .A3(new_n478), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  AOI22_X1  g202(.A1(G123), .A2(new_n485), .B1(new_n486), .B2(G135), .ZN(new_n628));
  OAI221_X1 g203(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n482), .C2(G111), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n626), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2430), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT82), .Z(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(new_n636), .B2(new_n637), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n641), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2443), .B(G2446), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT83), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n646), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(new_n650), .A3(G14), .ZN(G401));
  XOR2_X1   g226(.A(G2072), .B(G2078), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n660), .B2(new_n654), .ZN(new_n661));
  INV_X1    g236(.A(new_n654), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n662), .B2(new_n659), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n654), .A2(new_n655), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n653), .B1(new_n664), .B2(KEYINPUT17), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n658), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(new_n631), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(new_n625), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n674), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n671), .A2(new_n675), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(KEYINPUT20), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(KEYINPUT20), .ZN(new_n681));
  AOI211_X1 g256(.A(new_n676), .B(new_n678), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n684), .B(new_n687), .ZN(G229));
  NOR2_X1   g263(.A1(G29), .A2(G33), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT89), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT90), .B(KEYINPUT25), .Z(new_n692));
  XOR2_X1   g267(.A(new_n691), .B(new_n692), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n486), .A2(G139), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT91), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n469), .A2(G127), .A3(new_n471), .ZN(new_n696));
  INV_X1    g271(.A(G115), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n465), .ZN(new_n698));
  AOI211_X1 g273(.A(new_n693), .B(new_n695), .C1(new_n463), .C2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n690), .B1(new_n699), .B2(G29), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n700), .A2(G2072), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT92), .ZN(new_n702));
  OR2_X1    g277(.A1(KEYINPUT24), .A2(G34), .ZN(new_n703));
  NAND2_X1  g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n704));
  AOI21_X1  g279(.A(G29), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G160), .B2(G29), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G2084), .ZN(new_n707));
  NOR2_X1   g282(.A1(G29), .A2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n485), .A2(G129), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT93), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n478), .A2(G105), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT26), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n712), .B(new_n714), .C1(new_n486), .C2(G141), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n708), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT94), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT27), .B(G1996), .ZN(new_n720));
  INV_X1    g295(.A(G1348), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n609), .A2(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G4), .B2(G16), .ZN(new_n723));
  OAI22_X1  g298(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n707), .B(new_n724), .C1(new_n721), .C2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(new_n720), .ZN(new_n726));
  NAND2_X1  g301(.A1(G164), .A2(G29), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G27), .B2(G29), .ZN(new_n728));
  INV_X1    g303(.A(G2078), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT86), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(KEYINPUT86), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(G19), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n560), .B2(new_n734), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G1341), .Z(new_n737));
  OR2_X1    g312(.A1(new_n728), .A2(new_n729), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n726), .A2(new_n730), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT31), .B(G11), .Z(new_n740));
  INV_X1    g315(.A(G28), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(KEYINPUT30), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT95), .ZN(new_n743));
  AOI21_X1  g318(.A(G29), .B1(new_n741), .B2(KEYINPUT30), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G29), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n630), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n731), .A2(G21), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G168), .B2(new_n731), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n747), .B1(G1966), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n732), .A2(G20), .A3(new_n733), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT23), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT97), .B(G1956), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n750), .B(new_n755), .C1(G1966), .C2(new_n749), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n700), .A2(G2072), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n753), .B2(new_n754), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n739), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G2090), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n763), .A2(G2090), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n731), .A2(G5), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G171), .B2(new_n731), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1961), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n746), .A2(G26), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT28), .ZN(new_n770));
  AOI22_X1  g345(.A1(G128), .A2(new_n485), .B1(new_n486), .B2(G140), .ZN(new_n771));
  OAI221_X1 g346(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n482), .C2(G116), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AND3_X1   g348(.A1(new_n773), .A2(KEYINPUT88), .A3(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(KEYINPUT88), .B1(new_n773), .B2(G29), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2067), .ZN(new_n777));
  NOR4_X1   g352(.A1(new_n764), .A2(new_n765), .A3(new_n768), .A4(new_n777), .ZN(new_n778));
  AND4_X1   g353(.A1(new_n702), .A2(new_n725), .A3(new_n759), .A4(new_n778), .ZN(new_n779));
  MUX2_X1   g354(.A(G6), .B(G305), .S(G16), .Z(new_n780));
  XOR2_X1   g355(.A(KEYINPUT32), .B(G1981), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n731), .A2(G23), .ZN(new_n783));
  INV_X1    g358(.A(G288), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n731), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT33), .B(G1976), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n734), .A2(G22), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G166), .B2(new_n734), .ZN(new_n789));
  INV_X1    g364(.A(G1971), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n782), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT34), .ZN(new_n794));
  NOR2_X1   g369(.A1(G25), .A2(G29), .ZN(new_n795));
  AOI22_X1  g370(.A1(G119), .A2(new_n485), .B1(new_n486), .B2(G131), .ZN(new_n796));
  OAI221_X1 g371(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n482), .C2(G107), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n795), .B1(new_n799), .B2(G29), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G24), .B(G290), .S(new_n734), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT87), .B(G1986), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n793), .A2(new_n794), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT36), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n779), .A2(new_n807), .ZN(G150));
  INV_X1    g383(.A(G150), .ZN(G311));
  NAND2_X1  g384(.A1(new_n609), .A2(G559), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(KEYINPUT99), .B1(new_n556), .B2(new_n559), .ZN(new_n813));
  INV_X1    g388(.A(G56), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n534), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(G651), .B1(new_n815), .B2(new_n554), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n547), .A2(G81), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n550), .A2(G43), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n517), .A2(G55), .A3(G543), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OAI221_X1 g398(.A(new_n821), .B1(new_n822), .B2(new_n524), .C1(new_n823), .C2(new_n515), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n813), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n823), .A2(new_n515), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n821), .B1(new_n822), .B2(new_n524), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n828), .A2(new_n560), .A3(new_n818), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n812), .B(new_n830), .Z(new_n831));
  OR2_X1    g406(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n832));
  INV_X1    g407(.A(G860), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(KEYINPUT39), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n828), .A2(new_n833), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n699), .B(new_n716), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n491), .A2(new_n495), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT100), .ZN(new_n841));
  INV_X1    g416(.A(new_n509), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n491), .A2(new_n495), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(new_n773), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n839), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n798), .B(new_n623), .ZN(new_n848));
  AOI22_X1  g423(.A1(G130), .A2(new_n485), .B1(new_n486), .B2(G142), .ZN(new_n849));
  OAI221_X1 g424(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n482), .C2(G118), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n848), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT101), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n847), .B(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n480), .B(new_n630), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n488), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n847), .A2(new_n853), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n847), .B2(new_n852), .ZN(new_n859));
  AOI21_X1  g434(.A(G37), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g437(.A1(new_n824), .A2(G868), .ZN(new_n863));
  XNOR2_X1  g438(.A(G305), .B(G303), .ZN(new_n864));
  XNOR2_X1  g439(.A(G288), .B(G290), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n864), .B(new_n865), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT42), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT102), .B1(new_n609), .B2(G299), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n609), .A2(G299), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n609), .A2(G299), .A3(KEYINPUT102), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT41), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OR3_X1    g447(.A1(new_n609), .A2(G299), .A3(KEYINPUT102), .ZN(new_n873));
  XNOR2_X1  g448(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n873), .A2(new_n868), .A3(new_n869), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n619), .B(new_n830), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n868), .A3(new_n869), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n877), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n867), .B(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n863), .B1(new_n881), .B2(G868), .ZN(G295));
  AOI21_X1  g457(.A(new_n863), .B1(new_n881), .B2(G868), .ZN(G331));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n879), .A2(KEYINPUT109), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT109), .B1(new_n879), .B2(new_n885), .ZN(new_n887));
  INV_X1    g462(.A(new_n537), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n550), .A2(G51), .B1(new_n530), .B2(new_n529), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT105), .B1(new_n533), .B2(new_n537), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n546), .A4(new_n551), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n546), .B2(new_n551), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n830), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(G301), .A2(KEYINPUT105), .A3(G286), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n897), .A2(new_n825), .A3(new_n829), .A4(new_n893), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n886), .A2(new_n887), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n879), .ZN(new_n900));
  INV_X1    g475(.A(new_n874), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n898), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n866), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(G37), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n900), .A2(new_n902), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n872), .A2(new_n875), .A3(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT106), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n872), .A2(new_n902), .A3(new_n875), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n907), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n866), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n906), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n884), .B1(new_n918), .B2(KEYINPUT111), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n905), .B1(new_n912), .B2(new_n913), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI211_X1 g497(.A(KEYINPUT107), .B(new_n905), .C1(new_n912), .C2(new_n913), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n914), .ZN(new_n925));
  OAI221_X1 g500(.A(new_n919), .B1(KEYINPUT111), .B2(new_n918), .C1(KEYINPUT43), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n906), .A2(new_n915), .A3(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n917), .B1(new_n924), .B2(new_n914), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(KEYINPUT108), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n915), .B1(new_n922), .B2(new_n923), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n932), .B1(new_n933), .B2(new_n917), .ZN(new_n934));
  AOI211_X1 g509(.A(KEYINPUT110), .B(new_n928), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n925), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n937));
  INV_X1    g512(.A(new_n929), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n939), .B2(new_n927), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n926), .B1(new_n935), .B2(new_n940), .ZN(G397));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n845), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n475), .A2(G40), .A3(new_n479), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n947), .A2(KEYINPUT112), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(KEYINPUT112), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1996), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT46), .Z(new_n953));
  INV_X1    g528(.A(new_n950), .ZN(new_n954));
  INV_X1    g529(.A(G2067), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n773), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n717), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n953), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT47), .ZN(new_n959));
  OR3_X1    g534(.A1(new_n954), .A2(G1986), .A3(G290), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n956), .B1(new_n717), .B2(new_n951), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n962), .B1(new_n951), .B2(new_n717), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n799), .A2(new_n801), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n799), .A2(new_n801), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  OAI22_X1  g542(.A1(new_n960), .A2(new_n961), .B1(new_n954), .B2(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n960), .A2(new_n961), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n773), .A2(G2067), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n965), .B(KEYINPUT127), .Z(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(new_n963), .B2(new_n971), .ZN(new_n972));
  OAI22_X1  g547(.A1(new_n968), .A2(new_n969), .B1(new_n954), .B2(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n959), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n942), .B1(new_n496), .B2(new_n509), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n945), .B1(new_n976), .B2(new_n944), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n845), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n790), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n980), .B(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(KEYINPUT50), .B1(new_n845), .B2(new_n942), .ZN(new_n983));
  OAI211_X1 g558(.A(KEYINPUT50), .B(new_n942), .C1(new_n496), .C2(new_n509), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n946), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(G2090), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n975), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(G166), .A2(new_n975), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n990));
  XNOR2_X1  g565(.A(new_n989), .B(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n976), .A2(new_n944), .ZN(new_n994));
  AOI21_X1  g569(.A(G1966), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G2084), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n997), .B(new_n946), .C1(new_n983), .C2(new_n985), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n992), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n988), .A2(new_n991), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n946), .A2(new_n845), .A3(new_n942), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1005), .A2(new_n975), .ZN(new_n1006));
  OR2_X1    g581(.A1(G305), .A2(G1981), .ZN(new_n1007));
  INV_X1    g582(.A(G86), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n586), .B1(new_n1008), .B2(new_n524), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n585), .B1(new_n1009), .B2(KEYINPUT115), .ZN(new_n1011));
  OAI21_X1  g586(.A(G1981), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1012), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  OAI221_X1 g592(.A(new_n1006), .B1(KEYINPUT49), .B2(new_n1013), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT52), .B1(G288), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1006), .B(new_n1020), .C1(new_n1019), .C2(G288), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1006), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G288), .A2(new_n1019), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT52), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AND3_X1   g599(.A1(new_n1018), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n999), .A2(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1027), .A2(G286), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(KEYINPUT63), .C1(new_n991), .C2(new_n988), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n1003), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT117), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1031), .A3(KEYINPUT63), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1018), .A2(new_n1019), .A3(new_n784), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1022), .B1(new_n1033), .B2(new_n1007), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1003), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(new_n1025), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1026), .A2(new_n1031), .A3(new_n1028), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n729), .A2(KEYINPUT53), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n945), .B(new_n1039), .C1(new_n943), .C2(new_n944), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n994), .ZN(new_n1041));
  INV_X1    g616(.A(G1961), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n986), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n977), .A2(new_n978), .A3(new_n729), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1041), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1047), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G168), .A2(new_n975), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n996), .A2(KEYINPUT123), .A3(new_n998), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT123), .ZN(new_n1052));
  INV_X1    g627(.A(new_n998), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1053), .B2(new_n995), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n1051), .B(new_n1054), .C1(KEYINPUT124), .C2(G168), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1050), .A2(KEYINPUT124), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1027), .A2(new_n1056), .A3(new_n1050), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  OAI221_X1 g637(.A(new_n1048), .B1(new_n1050), .B2(new_n1055), .C1(new_n1060), .C2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1047), .A2(G171), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1064), .A2(KEYINPUT62), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT56), .B(G2072), .Z(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n978), .A2(new_n977), .A3(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(G299), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n1070));
  AND2_X1   g645(.A1(G299), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n845), .A2(KEYINPUT50), .A3(new_n942), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT50), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n976), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n945), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1068), .B(new_n1072), .C1(new_n1076), .C2(G1956), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1068), .B1(new_n1076), .B2(G1956), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1072), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n986), .A2(new_n721), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1005), .A2(new_n955), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n618), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1077), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1078), .B1(new_n1071), .B2(new_n1069), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT61), .B1(new_n1087), .B2(new_n1077), .ZN(new_n1088));
  XNOR2_X1  g663(.A(new_n1088), .B(KEYINPUT122), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT58), .B(G1341), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n979), .A2(G1996), .B1(new_n1005), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n616), .B1(KEYINPUT120), .B2(KEYINPUT59), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT121), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1095), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1097), .A3(new_n1092), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n618), .A2(KEYINPUT60), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1096), .A2(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1083), .A2(new_n618), .A3(new_n1084), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1085), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1077), .A2(KEYINPUT61), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1101), .B(new_n1103), .C1(new_n1082), .C2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1086), .B1(new_n1089), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1043), .A2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1040), .A2(new_n978), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n986), .A2(KEYINPUT125), .A3(new_n1042), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(G301), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT54), .B1(new_n1111), .B2(new_n1064), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT126), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1047), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(G301), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1112), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1065), .B1(new_n1106), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1055), .A2(new_n1050), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1060), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1125), .B2(new_n1061), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1038), .B(new_n1063), .C1(new_n1123), .C2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G2090), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1076), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n980), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n991), .B1(new_n1130), .B2(G8), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1030), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1037), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(G290), .B(G1986), .Z(new_n1134));
  AOI21_X1  g709(.A(new_n954), .B1(new_n967), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n974), .B1(new_n1133), .B2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g711(.A1(new_n668), .A2(G319), .ZN(new_n1138));
  NOR3_X1   g712(.A1(G401), .A2(G229), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n939), .A2(new_n861), .A3(new_n1139), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


