//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT87), .B(G469), .Z(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n189), .A2(G146), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT67), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n193), .A2(new_n200), .A3(new_n195), .A4(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n203));
  OAI21_X1  g017(.A(G128), .B1(new_n194), .B2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G146), .B1(new_n190), .B2(new_n192), .ZN(new_n205));
  INV_X1    g019(.A(G146), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT65), .B1(new_n206), .B2(G143), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(new_n189), .A3(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI211_X1 g024(.A(KEYINPUT68), .B(new_n204), .C1(new_n205), .C2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G143), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n207), .B(new_n209), .C1(new_n213), .C2(G146), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT68), .B1(new_n214), .B2(new_n204), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n202), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n217), .B1(new_n218), .B2(G107), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(G107), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(KEYINPUT84), .A3(G104), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G101), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n218), .B2(G107), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n221), .A3(G104), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n225), .A2(new_n227), .A3(new_n228), .A4(new_n220), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT85), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT85), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n224), .A2(new_n232), .A3(new_n229), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(G128), .B1(new_n205), .B2(new_n203), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n193), .A2(new_n195), .ZN(new_n236));
  AOI22_X1  g050(.A1(new_n199), .A2(new_n201), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI22_X1  g051(.A1(new_n216), .A2(new_n234), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G134), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT11), .B1(new_n239), .B2(G137), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT66), .B1(new_n242), .B2(G134), .ZN(new_n245));
  OR3_X1    g059(.A1(new_n242), .A2(KEYINPUT66), .A3(G134), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n244), .A2(new_n249), .A3(new_n246), .A4(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n238), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n238), .A2(KEYINPUT12), .A3(new_n251), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n216), .A2(KEYINPUT10), .A3(new_n234), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT86), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n204), .B1(new_n205), .B2(new_n210), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n211), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n259), .B1(new_n263), .B2(new_n202), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT86), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(new_n234), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n251), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n259), .B1(new_n237), .B2(new_n230), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n270));
  AND2_X1   g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NOR2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g087(.A1(new_n207), .A2(new_n209), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n191), .A2(G143), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n189), .A2(KEYINPUT64), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n206), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n193), .A2(new_n195), .A3(new_n271), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n270), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n193), .A2(new_n195), .A3(new_n271), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n205), .A2(new_n210), .ZN(new_n282));
  OAI211_X1 g096(.A(KEYINPUT71), .B(new_n281), .C1(new_n282), .C2(new_n273), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n225), .A2(new_n227), .A3(new_n220), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(G101), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(G101), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n280), .A2(new_n283), .A3(new_n286), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n269), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n267), .A2(new_n268), .A3(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n256), .A2(new_n292), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n265), .B1(new_n264), .B2(new_n234), .ZN(new_n299));
  AND4_X1   g113(.A1(new_n265), .A2(new_n216), .A3(KEYINPUT10), .A4(new_n234), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n291), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n251), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n297), .B1(new_n302), .B2(new_n292), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT88), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n268), .B1(new_n267), .B2(new_n291), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n251), .B(new_n290), .C1(new_n258), .C2(new_n266), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n296), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(KEYINPUT88), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n187), .B(new_n188), .C1(new_n305), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT89), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(KEYINPUT88), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n303), .A2(new_n304), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n298), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n315), .A2(KEYINPUT89), .A3(new_n187), .A4(new_n188), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G469), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n307), .A2(new_n296), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n302), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n256), .A2(new_n292), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n296), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n318), .B1(new_n323), .B2(new_n187), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n317), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G221), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT9), .B(G234), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(new_n187), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G237), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n294), .A3(G214), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n190), .A3(new_n192), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n332), .A2(new_n294), .A3(G143), .A4(G214), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G131), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT93), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT93), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n339), .A3(G131), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT95), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT17), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n334), .A2(new_n249), .A3(new_n335), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT16), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n348), .A2(G140), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(KEYINPUT16), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n206), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n347), .B(G146), .C1(KEYINPUT16), .C2(new_n349), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n339), .B1(new_n336), .B2(G131), .ZN(new_n354));
  AOI211_X1 g168(.A(KEYINPUT93), .B(new_n249), .C1(new_n334), .C2(new_n335), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n353), .B1(KEYINPUT17), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n344), .B(new_n343), .C1(new_n354), .C2(new_n355), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT95), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n345), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n346), .B(new_n206), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT18), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n249), .ZN(new_n363));
  OAI221_X1 g177(.A(new_n361), .B1(new_n336), .B2(new_n363), .C1(new_n337), .C2(new_n362), .ZN(new_n364));
  XNOR2_X1  g178(.A(G113), .B(G122), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(G104), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(KEYINPUT94), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n341), .A2(new_n344), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n346), .B(KEYINPUT19), .Z(new_n370));
  OAI21_X1  g184(.A(new_n352), .B1(new_n370), .B2(G146), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n364), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n366), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(G475), .A2(G902), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT92), .B(KEYINPUT20), .Z(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n374), .A2(new_n380), .A3(new_n375), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n368), .ZN(new_n383));
  INV_X1    g197(.A(new_n366), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n360), .B2(new_n364), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n187), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT96), .B(G475), .Z(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n213), .A2(G128), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n196), .A2(G143), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n239), .A3(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G116), .B(G122), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n393), .B(new_n221), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n390), .A2(KEYINPUT13), .A3(new_n391), .ZN(new_n395));
  OAI21_X1  g209(.A(G134), .B1(new_n390), .B2(KEYINPUT13), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n392), .B(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G116), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n221), .B1(new_n399), .B2(KEYINPUT14), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n393), .ZN(new_n401));
  INV_X1    g215(.A(new_n392), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n239), .B1(new_n390), .B2(new_n391), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n397), .A2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n329), .A2(G217), .A3(new_n294), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n397), .A2(new_n404), .A3(new_n406), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n187), .ZN(new_n411));
  INV_X1    g225(.A(G478), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(KEYINPUT15), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n397), .A2(new_n404), .A3(new_n406), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n406), .B1(new_n397), .B2(new_n404), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n187), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(KEYINPUT97), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT97), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n415), .B1(new_n410), .B2(new_n187), .ZN(new_n421));
  INV_X1    g235(.A(new_n418), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G952), .ZN(new_n425));
  AOI211_X1 g239(.A(G953), .B(new_n425), .C1(G234), .C2(G237), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(G898), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT98), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n187), .B(new_n294), .C1(G234), .C2(G237), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n426), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(new_n431), .B(KEYINPUT99), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n389), .A2(new_n424), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G214), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G110), .B(G122), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT2), .ZN(new_n440));
  INV_X1    g254(.A(G113), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT70), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT70), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(KEYINPUT2), .B2(G113), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(KEYINPUT2), .A2(G113), .ZN(new_n446));
  XNOR2_X1  g260(.A(G116), .B(G119), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n441), .B1(new_n447), .B2(KEYINPUT5), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT5), .ZN(new_n451));
  INV_X1    g265(.A(G119), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n452), .A3(G116), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT90), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n449), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n234), .A2(new_n439), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n445), .A2(new_n446), .ZN(new_n457));
  INV_X1    g271(.A(new_n447), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n448), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n286), .A3(new_n288), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n439), .B1(new_n234), .B2(new_n455), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n438), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n463), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n465), .A2(new_n437), .A3(new_n461), .A4(new_n456), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT6), .ZN(new_n467));
  INV_X1    g281(.A(G224), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n262), .A2(new_n211), .B1(new_n201), .B2(new_n199), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n278), .A2(new_n279), .A3(new_n348), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n216), .B2(new_n348), .ZN(new_n474));
  INV_X1    g288(.A(new_n469), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(new_n438), .C1(new_n462), .C2(new_n463), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n467), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n473), .B(new_n476), .C1(KEYINPUT7), .C2(new_n469), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n437), .B(KEYINPUT8), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n234), .A2(new_n455), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n455), .B1(new_n229), .B2(new_n224), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n474), .A2(new_n487), .A3(new_n475), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n481), .A2(new_n466), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n187), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G210), .B1(G237), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n480), .A2(new_n489), .A3(new_n187), .A4(new_n491), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n436), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n434), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n326), .A2(new_n331), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT100), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n324), .B1(new_n312), .B2(new_n316), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n499), .A2(new_n330), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT100), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n496), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G472), .A2(G902), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n239), .A2(G137), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n242), .A2(G134), .ZN(new_n506));
  OAI21_X1  g320(.A(G131), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n250), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT69), .B1(new_n470), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT69), .ZN(new_n510));
  INV_X1    g324(.A(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n216), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n278), .A2(new_n279), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n251), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n509), .A2(new_n512), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT73), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n508), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n250), .A2(KEYINPUT73), .A3(new_n507), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n263), .A2(new_n202), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n280), .A2(new_n251), .A3(new_n283), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n280), .A2(KEYINPUT72), .A3(new_n251), .A4(new_n283), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n516), .B1(new_n525), .B2(new_n515), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n460), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT31), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n447), .B1(new_n445), .B2(new_n446), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n449), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT74), .B1(new_n459), .B2(new_n448), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n525), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT75), .B(KEYINPUT27), .Z(new_n535));
  NAND3_X1  g349(.A1(new_n332), .A2(new_n294), .A3(G210), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT26), .B(G101), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n527), .A2(new_n528), .A3(new_n534), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT76), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n531), .A2(new_n532), .ZN(new_n542));
  AOI211_X1 g356(.A(new_n542), .B(new_n520), .C1(new_n523), .C2(new_n524), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n526), .B2(new_n460), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT76), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n528), .A4(new_n539), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n539), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT28), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n509), .A2(new_n512), .A3(new_n514), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n460), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n534), .B2(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n250), .A2(KEYINPUT73), .A3(new_n507), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT73), .B1(new_n250), .B2(new_n507), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n533), .B(new_n521), .C1(new_n470), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n549), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT77), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n559), .A3(new_n549), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n548), .B1(new_n552), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT78), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n527), .A2(new_n534), .A3(new_n539), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT31), .ZN(new_n566));
  OAI211_X1 g380(.A(KEYINPUT78), .B(new_n548), .C1(new_n552), .C2(new_n561), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n504), .B1(new_n547), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT32), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n504), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n547), .B2(new_n568), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT80), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n523), .A2(new_n524), .ZN(new_n577));
  INV_X1    g391(.A(new_n520), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n533), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT28), .B1(new_n543), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n556), .A2(new_n559), .A3(new_n549), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n559), .B1(new_n556), .B2(new_n549), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n558), .A2(KEYINPUT79), .A3(new_n560), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n548), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n580), .A2(new_n584), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n544), .A2(new_n548), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n539), .B1(new_n552), .B2(new_n561), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(new_n187), .B(new_n588), .C1(new_n591), .C2(KEYINPUT29), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  OAI211_X1 g407(.A(KEYINPUT80), .B(new_n573), .C1(new_n547), .C2(new_n568), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n571), .A2(new_n576), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G234), .ZN(new_n596));
  OAI21_X1  g410(.A(G217), .B1(new_n596), .B2(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n452), .A2(G128), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n452), .A2(G128), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(KEYINPUT23), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT24), .B(G110), .Z(new_n602));
  XNOR2_X1  g416(.A(G119), .B(G128), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n601), .A2(G110), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n353), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT81), .B(G110), .Z(new_n606));
  OAI22_X1  g420(.A1(new_n601), .A2(new_n606), .B1(new_n602), .B2(new_n603), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n346), .A2(new_n206), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n352), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT22), .B(G137), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n327), .A2(new_n596), .A3(G953), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n611), .B(new_n612), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n610), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT82), .B1(new_n615), .B2(G902), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT25), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n597), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n617), .B2(new_n616), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n597), .A2(new_n187), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT83), .Z(new_n621));
  NAND2_X1  g435(.A1(new_n614), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n595), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n503), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT101), .B(G101), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G3));
  OAI21_X1  g442(.A(new_n187), .B1(new_n547), .B2(new_n568), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(G472), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n569), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n623), .ZN(new_n632));
  INV_X1    g446(.A(new_n389), .ZN(new_n633));
  NAND2_X1  g447(.A1(KEYINPUT102), .A2(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n410), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(KEYINPUT102), .A2(KEYINPUT33), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n637), .A2(G478), .A3(new_n187), .ZN(new_n638));
  AOI21_X1  g452(.A(G478), .B1(new_n410), .B2(new_n187), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n495), .A2(new_n432), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n632), .A2(new_n500), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n218), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT103), .B(KEYINPUT34), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n374), .A2(new_n377), .A3(new_n375), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n377), .B1(new_n374), .B2(new_n375), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n388), .B(new_n424), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n649), .B1(new_n653), .B2(new_n433), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n379), .A2(new_n650), .B1(new_n386), .B2(new_n387), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n655), .A2(KEYINPUT104), .A3(new_n424), .A4(new_n432), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n654), .A2(new_n656), .A3(new_n495), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT105), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n654), .A2(new_n656), .A3(new_n495), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n632), .A2(new_n500), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  INV_X1    g478(.A(new_n613), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n610), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n621), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n619), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n631), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n503), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  INV_X1    g488(.A(new_n495), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n576), .A2(new_n594), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n541), .A2(new_n546), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n572), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n593), .B1(new_n680), .B2(KEYINPUT32), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n676), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n430), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n426), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n653), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n326), .A2(new_n331), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n682), .B2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n688), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n499), .A2(new_n330), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n692), .A2(new_n595), .A3(new_n693), .A4(new_n676), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NAND2_X1  g510(.A1(new_n493), .A2(new_n494), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(KEYINPUT38), .Z(new_n698));
  AOI22_X1  g512(.A1(new_n382), .A2(new_n388), .B1(new_n419), .B2(new_n423), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n698), .A2(new_n436), .A3(new_n700), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n543), .A2(new_n579), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n187), .B1(new_n702), .B2(new_n539), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n544), .A2(new_n548), .ZN(new_n704));
  OAI21_X1  g518(.A(G472), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n571), .A2(new_n576), .A3(new_n594), .A4(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n701), .A2(new_n670), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT107), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n686), .B(KEYINPUT39), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n500), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT40), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(new_n712), .B(new_n213), .Z(G45));
  NOR3_X1   g527(.A1(new_n499), .A2(new_n330), .A3(new_n687), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n595), .A3(new_n641), .A4(new_n676), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  AOI21_X1  g530(.A(new_n318), .B1(new_n315), .B2(new_n187), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n330), .B(new_n717), .C1(new_n312), .C2(new_n316), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n595), .A2(new_n718), .A3(new_n624), .A4(new_n644), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND4_X1  g535(.A1(new_n595), .A2(new_n661), .A3(new_n718), .A4(new_n624), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NAND4_X1  g537(.A1(new_n595), .A2(new_n718), .A3(new_n434), .A4(new_n676), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND3_X1  g539(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n548), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT108), .A3(new_n566), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n679), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT108), .B1(new_n727), .B2(new_n566), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n504), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT109), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(new_n504), .C1(new_n729), .C2(new_n730), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n732), .A2(new_n624), .A3(new_n630), .A4(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n717), .B1(new_n312), .B2(new_n316), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n643), .A2(new_n700), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(new_n331), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n398), .ZN(G24));
  NAND4_X1  g554(.A1(new_n732), .A2(new_n630), .A3(new_n669), .A4(new_n734), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT110), .ZN(new_n742));
  AOI22_X1  g556(.A1(new_n731), .A2(KEYINPUT109), .B1(G472), .B2(new_n629), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n669), .A4(new_n734), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n718), .A2(new_n495), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n642), .A2(new_n687), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  NAND3_X1  g566(.A1(new_n493), .A2(new_n435), .A3(new_n494), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n499), .A2(new_n330), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n595), .A3(new_n624), .A4(new_n748), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n569), .A2(new_n570), .B1(G472), .B2(new_n592), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n623), .B1(new_n758), .B2(new_n574), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n759), .A2(new_n754), .A3(KEYINPUT42), .A4(new_n748), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  AND4_X1   g576(.A1(new_n595), .A2(new_n754), .A3(new_n624), .A4(new_n688), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n239), .ZN(G36));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n323), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n320), .A2(KEYINPUT45), .A3(new_n322), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(G469), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n769), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n770), .A2(KEYINPUT111), .A3(new_n771), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n774), .A2(new_n317), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n331), .A3(new_n709), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n753), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n680), .B1(G472), .B2(new_n629), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n783), .B2(new_n670), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n631), .A2(KEYINPUT115), .A3(new_n669), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  XOR2_X1   g601(.A(new_n640), .B(KEYINPUT113), .Z(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n389), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n640), .A2(new_n389), .A3(new_n787), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT114), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n786), .A2(KEYINPUT44), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n792), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n780), .A2(new_n781), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NAND2_X1  g612(.A1(new_n777), .A2(new_n331), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n595), .A2(new_n749), .A3(new_n624), .A4(new_n753), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  XOR2_X1   g618(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n675), .A2(new_n700), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n714), .A2(new_n706), .A3(new_n670), .A4(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n715), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n751), .A2(new_n809), .A3(new_n695), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n751), .A2(new_n809), .A3(new_n695), .A4(KEYINPUT52), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n763), .B1(new_n757), .B2(new_n760), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n722), .B1(new_n735), .B2(new_n738), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n414), .A2(new_n418), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(KEYINPUT116), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n389), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n641), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n643), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n500), .A2(new_n821), .A3(new_n624), .A4(new_n783), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n719), .A2(new_n724), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n816), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n502), .B(new_n498), .C1(new_n625), .C2(new_n671), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n655), .A2(new_n669), .A3(new_n686), .A4(new_n818), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n754), .A2(new_n595), .A3(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n754), .A2(new_n748), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n746), .B2(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n815), .A2(new_n824), .A3(new_n825), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n814), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n806), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n824), .A2(new_n815), .A3(new_n825), .A4(new_n829), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n832), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n751), .A2(new_n836), .A3(new_n695), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n751), .B2(new_n695), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n500), .A2(new_n686), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n641), .B(new_n676), .C1(new_n677), .C2(new_n681), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n705), .B1(new_n680), .B2(KEYINPUT32), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n670), .B(new_n807), .C1(new_n677), .C2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n694), .B2(new_n690), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT52), .B1(new_n846), .B2(new_n751), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n835), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT52), .A2(new_n751), .A3(new_n809), .A4(new_n695), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n851), .A2(new_n832), .A3(new_n834), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n830), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n834), .A2(KEYINPUT117), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n854), .B(new_n855), .C1(new_n840), .C2(new_n847), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n852), .B1(new_n856), .B2(new_n832), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n736), .ZN(new_n860));
  NOR4_X1   g674(.A1(new_n860), .A2(new_n330), .A3(new_n685), .A4(new_n753), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n706), .A2(new_n623), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n389), .A2(new_n639), .A3(new_n638), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n746), .A2(new_n792), .A3(new_n861), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n792), .A2(new_n426), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n870), .A2(new_n735), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n718), .A2(new_n436), .A3(new_n698), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT50), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n753), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n860), .A2(new_n331), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n875), .B1(new_n801), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n869), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n869), .A2(KEYINPUT51), .A3(new_n874), .A4(new_n877), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n861), .A2(new_n792), .A3(new_n759), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT48), .Z(new_n883));
  NOR2_X1   g697(.A1(new_n871), .A2(new_n747), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n863), .A2(new_n641), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(G952), .A3(new_n294), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n883), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n880), .A2(new_n881), .A3(new_n887), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n859), .A2(new_n888), .B1(G952), .B2(G953), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n640), .A2(new_n330), .A3(new_n436), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n698), .A2(new_n633), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n860), .B2(KEYINPUT49), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n892), .B(new_n862), .C1(KEYINPUT49), .C2(new_n860), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n889), .A2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n294), .A2(G952), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n895), .B(KEYINPUT121), .Z(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n467), .A2(new_n479), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n477), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT55), .Z(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n832), .B1(new_n851), .B2(new_n834), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n848), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(G210), .A3(G902), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n901), .B1(new_n905), .B2(KEYINPUT56), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n904), .A2(new_n907), .A3(new_n900), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n897), .B1(new_n906), .B2(new_n908), .ZN(G51));
  XOR2_X1   g723(.A(new_n769), .B(KEYINPUT57), .Z(new_n910));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n902), .A2(new_n848), .A3(new_n911), .A4(new_n805), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n719), .A2(new_n724), .A3(new_n822), .ZN(new_n913));
  AND4_X1   g727(.A1(new_n595), .A2(new_n661), .A3(new_n718), .A4(new_n624), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n739), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n913), .A2(new_n915), .A3(new_n825), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(KEYINPUT53), .A3(new_n815), .A4(new_n829), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n751), .A2(new_n695), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT118), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n751), .A2(new_n695), .A3(new_n836), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(KEYINPUT52), .A3(new_n920), .A4(new_n809), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n917), .B1(new_n921), .B2(new_n812), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT53), .B1(new_n814), .B2(new_n830), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n806), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n912), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n911), .B1(new_n833), .B2(new_n848), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n910), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n315), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n922), .A2(new_n923), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n929), .A2(new_n187), .A3(new_n768), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n895), .B1(new_n928), .B2(new_n930), .ZN(G54));
  AND2_X1   g745(.A1(KEYINPUT58), .A2(G475), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n903), .A2(G902), .A3(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n374), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n933), .A2(KEYINPUT123), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT123), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n933), .A2(new_n934), .ZN(new_n937));
  NOR4_X1   g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n895), .ZN(G60));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT59), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n637), .B(new_n940), .C1(new_n925), .C2(new_n926), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n896), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n637), .B1(new_n859), .B2(new_n940), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n615), .B1(new_n929), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n903), .A2(new_n667), .A3(new_n946), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(new_n896), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n429), .B2(new_n468), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n916), .B2(G953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n898), .B1(G898), .B2(new_n294), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  NAND3_X1  g770(.A1(new_n780), .A2(new_n759), .A3(new_n807), .ZN(new_n957));
  AND4_X1   g771(.A1(new_n797), .A2(new_n957), .A3(new_n803), .A4(new_n815), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n837), .A2(new_n838), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n715), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n958), .A2(new_n294), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n683), .A2(new_n294), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(G227), .A2(G900), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n526), .B(new_n370), .Z(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(G953), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n961), .B2(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(G953), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n797), .A2(new_n803), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n820), .A2(new_n753), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n625), .A2(new_n710), .A3(new_n970), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT125), .Z(new_n972));
  NAND3_X1  g786(.A1(new_n959), .A2(new_n712), .A3(new_n715), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n969), .B(new_n972), .C1(new_n973), .C2(KEYINPUT62), .ZN(new_n974));
  INV_X1    g788(.A(new_n973), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT124), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n973), .A2(new_n978), .A3(KEYINPUT62), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n974), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n965), .A2(G953), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n967), .B(new_n968), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n966), .A2(new_n982), .ZN(G72));
  INV_X1    g797(.A(new_n704), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n977), .A2(new_n979), .ZN(new_n985));
  INV_X1    g799(.A(new_n974), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n916), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  AOI21_X1  g803(.A(new_n984), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n958), .A2(new_n916), .A3(new_n960), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n989), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n589), .B(KEYINPUT126), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n895), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n984), .A2(new_n589), .A3(new_n989), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT127), .Z(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n857), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n990), .A2(new_n997), .ZN(G57));
endmodule


