//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1343, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n203), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n204), .A2(new_n205), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n209), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT0), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n219), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G68), .Z(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G1), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G274), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT66), .B(G41), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n249), .B1(new_n250), .B2(G45), .ZN(new_n251));
  INV_X1    g0051(.A(G226), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n247), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n251), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1698), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G222), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G77), .ZN(new_n267));
  INV_X1    g0067(.A(G223), .ZN(new_n268));
  XNOR2_X1  g0068(.A(KEYINPUT3), .B(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G1698), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n263), .B(new_n267), .C1(new_n268), .C2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n257), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G179), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n223), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n224), .B1(new_n220), .B2(new_n221), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n224), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G150), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  OAI22_X1  g0083(.A1(new_n279), .A2(new_n280), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n277), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n286), .A2(new_n224), .A3(G1), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n277), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n221), .B1(new_n247), .B2(G20), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(new_n289), .B1(new_n221), .B2(new_n287), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n275), .B(new_n291), .C1(G169), .C2(new_n273), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g0093(.A(new_n291), .ZN(new_n294));
  INV_X1    g0094(.A(new_n273), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT67), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(new_n298), .A3(new_n275), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n293), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n277), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n279), .A2(new_n283), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(G20), .B2(G77), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT15), .B(G87), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(new_n280), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n247), .A2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n288), .A2(G77), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n286), .A2(G1), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(G77), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G244), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n251), .B1(new_n313), .B2(new_n256), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n262), .A2(G232), .ZN(new_n315));
  INV_X1    g0115(.A(G107), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n315), .B1(new_n316), .B2(new_n269), .C1(new_n211), .C2(new_n270), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n314), .B1(new_n317), .B2(new_n272), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n312), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(G190), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n312), .B(KEYINPUT68), .C1(new_n319), .C2(new_n318), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n317), .A2(new_n272), .ZN(new_n326));
  INV_X1    g0126(.A(new_n314), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n296), .ZN(new_n329));
  INV_X1    g0129(.A(new_n312), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n318), .A2(new_n274), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n300), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT9), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n291), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n335), .B(KEYINPUT69), .Z(new_n336));
  INV_X1    g0136(.A(KEYINPUT10), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT70), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n295), .B2(G200), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n294), .A2(KEYINPUT9), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n273), .A2(G190), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n336), .A2(new_n337), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n341), .A3(new_n340), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n335), .B(KEYINPUT69), .ZN(new_n345));
  OAI21_X1  g0145(.A(KEYINPUT10), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n269), .B2(G20), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n266), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n203), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G58), .A2(G68), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n204), .A2(new_n205), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n282), .A2(G159), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n348), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT7), .B1(new_n266), .B2(new_n224), .ZN(new_n359));
  NOR4_X1   g0159(.A1(new_n264), .A2(new_n265), .A3(new_n349), .A4(G20), .ZN(new_n360));
  OAI21_X1  g0160(.A(G68), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n354), .A2(G20), .B1(G159), .B2(new_n282), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(KEYINPUT16), .A3(new_n362), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n358), .A2(new_n363), .A3(new_n277), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n279), .B1(new_n247), .B2(G20), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n365), .A2(new_n288), .B1(new_n287), .B2(new_n279), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT18), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n251), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G33), .A2(G87), .ZN(new_n372));
  INV_X1    g0172(.A(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n268), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n252), .A2(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n372), .B1(new_n376), .B2(new_n266), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n272), .ZN(new_n378));
  AOI21_X1  g0178(.A(G169), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT66), .A2(G41), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT66), .A2(G41), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G45), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n248), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT77), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n251), .A2(new_n387), .A3(new_n369), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n269), .A2(new_n374), .A3(new_n375), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n254), .B1(new_n390), .B2(new_n372), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n391), .A2(G179), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n379), .B1(new_n389), .B2(new_n392), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n367), .A2(new_n368), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n368), .B1(new_n367), .B2(new_n393), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n386), .A2(new_n397), .A3(new_n378), .A4(new_n388), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n319), .B1(new_n391), .B2(new_n370), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n364), .A2(new_n400), .A3(new_n366), .ZN(new_n401));
  XNOR2_X1  g0201(.A(new_n401), .B(KEYINPUT17), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n333), .A2(new_n347), .A3(new_n396), .A4(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT75), .B1(new_n310), .B2(G68), .ZN(new_n404));
  XOR2_X1   g0204(.A(new_n404), .B(KEYINPUT12), .Z(new_n405));
  NAND3_X1  g0205(.A1(new_n288), .A2(G68), .A3(new_n307), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT11), .ZN(new_n407));
  INV_X1    g0207(.A(G77), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n280), .A2(new_n408), .B1(new_n224), .B2(G68), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n409), .A2(KEYINPUT74), .B1(new_n221), .B2(new_n283), .ZN(new_n410));
  AND2_X1   g0210(.A1(new_n409), .A2(KEYINPUT74), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n277), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OAI211_X1 g0212(.A(new_n405), .B(new_n406), .C1(new_n407), .C2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n407), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  OAI211_X1 g0216(.A(G232), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT71), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n269), .A2(KEYINPUT71), .A3(G232), .A4(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G97), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n269), .A2(G226), .A3(new_n373), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n272), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n254), .A2(G238), .A3(new_n255), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n251), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n416), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  AOI211_X1 g0228(.A(KEYINPUT13), .B(new_n426), .C1(new_n423), .C2(new_n272), .ZN(new_n429));
  OAI21_X1  g0229(.A(G169), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT14), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT14), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(G169), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT73), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n426), .B1(new_n423), .B2(new_n272), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT72), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT13), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI211_X1 g0238(.A(KEYINPUT72), .B(new_n426), .C1(new_n423), .C2(new_n272), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n424), .A2(new_n427), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT72), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n436), .A2(new_n437), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n442), .A2(KEYINPUT73), .A3(KEYINPUT13), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n429), .A2(new_n274), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT76), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n434), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n446), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n440), .B2(new_n444), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n431), .A2(new_n433), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT76), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n415), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n429), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G190), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n440), .B2(new_n444), .ZN(new_n457));
  OAI21_X1  g0257(.A(G200), .B1(new_n428), .B2(new_n429), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n415), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n403), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n247), .B(G45), .C1(new_n462), .C2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n380), .B2(new_n381), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n272), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n250), .B2(new_n462), .ZN(new_n467));
  INV_X1    g0267(.A(G274), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n272), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n466), .A2(G270), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g0270(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n471));
  OAI211_X1 g0271(.A(G257), .B(new_n373), .C1(new_n264), .C2(new_n265), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n260), .A2(G303), .A3(new_n261), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n272), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT88), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(KEYINPUT88), .A3(new_n475), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n310), .A2(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n247), .A2(G33), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(KEYINPUT79), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n247), .B2(G33), .ZN(new_n485));
  NOR4_X1   g0285(.A1(new_n483), .A2(new_n287), .A3(new_n485), .A4(new_n277), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n481), .B1(new_n486), .B2(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n224), .C1(G33), .C2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n490), .B(new_n277), .C1(new_n224), .C2(G116), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT20), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n491), .B(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n296), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT21), .B1(new_n480), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(KEYINPUT88), .B1(new_n470), .B2(new_n475), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n466), .A2(G270), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n467), .A2(new_n469), .ZN(new_n498));
  AND4_X1   g0298(.A1(KEYINPUT88), .A2(new_n475), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n494), .B(KEYINPUT21), .C1(new_n496), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n493), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n274), .B1(new_n474), .B2(new_n272), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n470), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT89), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n500), .A2(KEYINPUT89), .A3(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n501), .B1(new_n480), .B2(G200), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n397), .B2(new_n480), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n283), .A2(new_n408), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n316), .A2(KEYINPUT6), .A3(G97), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  XNOR2_X1  g0315(.A(G97), .B(G107), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(KEYINPUT78), .B(new_n512), .C1(new_n517), .C2(new_n224), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT78), .ZN(new_n519));
  AND2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n224), .B1(new_n522), .B2(new_n513), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n519), .B1(new_n523), .B2(new_n511), .ZN(new_n524));
  OAI21_X1  g0324(.A(G107), .B1(new_n359), .B2(new_n360), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n518), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n277), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n310), .A2(G97), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n486), .B2(G97), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G250), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n531));
  OAI211_X1 g0331(.A(G244), .B(new_n373), .C1(new_n264), .C2(new_n265), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT4), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n488), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT4), .B1(new_n262), .B2(G244), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n272), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n466), .A2(G257), .B1(new_n467), .B2(new_n469), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n538), .A2(new_n397), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n530), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n537), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(KEYINPUT80), .B(new_n272), .C1(new_n534), .C2(new_n535), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n541), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT81), .ZN(new_n546));
  OAI21_X1  g0346(.A(G200), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n532), .A2(new_n533), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n269), .A2(KEYINPUT4), .A3(G244), .A4(new_n373), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(new_n488), .A4(new_n531), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT80), .B1(new_n551), .B2(new_n272), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n537), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n540), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n527), .A2(new_n529), .B1(new_n296), .B2(new_n538), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n274), .B(new_n537), .C1(new_n548), .C2(new_n552), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT83), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT83), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n269), .A2(new_n562), .A3(G244), .A4(G1698), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g0364(.A(G238), .B(new_n373), .C1(new_n264), .C2(new_n265), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G33), .A2(G116), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n254), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  OAI22_X1  g0369(.A1(KEYINPUT82), .A2(new_n213), .B1(new_n383), .B2(G1), .ZN(new_n570));
  NAND2_X1  g0370(.A1(KEYINPUT82), .A2(G250), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n571), .A2(new_n247), .A3(G45), .A4(new_n468), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n572), .A3(new_n254), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n569), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT84), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT84), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT19), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n421), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n576), .B1(new_n581), .B2(G20), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n521), .A2(new_n212), .ZN(new_n583));
  XNOR2_X1  g0383(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n584));
  OAI211_X1 g0384(.A(KEYINPUT85), .B(new_n224), .C1(new_n584), .C2(new_n421), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n224), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT86), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT86), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n269), .A2(new_n589), .A3(new_n224), .A4(G68), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n224), .A2(G33), .A3(G97), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(new_n578), .A3(new_n580), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n584), .A2(KEYINPUT87), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n277), .B1(new_n586), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n304), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(new_n310), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n486), .A2(G87), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n575), .A2(new_n599), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n567), .B1(new_n563), .B2(new_n561), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n573), .B1(new_n605), .B2(new_n254), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(new_n397), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n482), .B(new_n484), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n288), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n304), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n611), .A2(new_n597), .A3(new_n591), .ZN(new_n612));
  AOI211_X1 g0412(.A(new_n601), .B(new_n610), .C1(new_n612), .C2(new_n277), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n274), .B(new_n573), .C1(new_n605), .C2(new_n254), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n564), .A2(new_n568), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n574), .B1(new_n615), .B2(new_n272), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(G169), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n604), .A2(new_n607), .B1(new_n613), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n269), .A2(G257), .A3(G1698), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n269), .A2(G250), .A3(new_n373), .ZN(new_n620));
  INV_X1    g0420(.A(G294), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n619), .B(new_n620), .C1(new_n259), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n272), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n466), .A2(G264), .B1(new_n467), .B2(new_n469), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n296), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n262), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n254), .B1(new_n627), .B2(new_n619), .ZN(new_n628));
  OR2_X1    g0428(.A1(KEYINPUT66), .A2(G41), .ZN(new_n629));
  NAND2_X1  g0429(.A1(KEYINPUT66), .A2(G41), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT5), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(G264), .B(new_n254), .C1(new_n631), .C2(new_n463), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n498), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n628), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n274), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n626), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n224), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT90), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(KEYINPUT22), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n269), .A2(new_n224), .A3(G87), .A4(new_n639), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(KEYINPUT22), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n224), .A2(G107), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT23), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT23), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n224), .B2(G107), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT91), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n566), .B2(G20), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n224), .A2(KEYINPUT91), .A3(G33), .A4(G116), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n646), .A2(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n644), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT24), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n301), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n644), .A2(new_n652), .A3(KEYINPUT24), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n309), .A2(new_n645), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT92), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT25), .ZN(new_n660));
  OR2_X1    g0460(.A1(new_n659), .A2(KEYINPUT25), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(KEYINPUT25), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n661), .A2(new_n309), .A3(new_n645), .A4(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n660), .B(new_n663), .C1(new_n609), .C2(new_n316), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n636), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n664), .B1(new_n655), .B2(new_n656), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n319), .B1(new_n628), .B2(new_n633), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n625), .B2(G190), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n559), .A2(new_n618), .A3(new_n672), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n461), .A2(new_n510), .A3(new_n673), .ZN(G372));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n618), .A2(new_n558), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n604), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n607), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n601), .B1(new_n612), .B2(new_n277), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(KEYINPUT93), .A3(new_n575), .A4(new_n603), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n558), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n613), .A2(new_n617), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n676), .B1(new_n675), .B2(new_n686), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n556), .A2(new_n557), .B1(new_n668), .B2(new_n670), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n555), .A2(new_n682), .A3(new_n685), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n626), .A2(new_n635), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n668), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n504), .A2(new_n691), .A3(new_n495), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n685), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n461), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n402), .ZN(new_n695));
  INV_X1    g0495(.A(new_n415), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n448), .B1(new_n434), .B2(new_n447), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n451), .A2(new_n452), .A3(KEYINPUT76), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n460), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n695), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n396), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n347), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n694), .A2(new_n705), .A3(new_n300), .ZN(G369));
  NAND2_X1  g0506(.A1(new_n309), .A2(new_n224), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G213), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G343), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n667), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n666), .A2(new_n712), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n667), .A2(new_n714), .A3(new_n671), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n691), .A2(new_n712), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT95), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(KEYINPUT95), .A3(new_n716), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n712), .B1(new_n506), .B2(new_n507), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n713), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n501), .A2(new_n712), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT94), .Z(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n504), .B2(new_n495), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n506), .A2(new_n726), .A3(new_n507), .A4(new_n509), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n721), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n723), .A2(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n227), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n250), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n583), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n222), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n738), .B2(new_n735), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  INV_X1    g0540(.A(new_n712), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n693), .B2(new_n687), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT29), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n504), .A2(new_n505), .ZN(new_n745));
  INV_X1    g0545(.A(new_n495), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n507), .A3(new_n746), .A4(new_n667), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n607), .B1(new_n604), .B2(new_n677), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n684), .B1(new_n748), .B2(new_n681), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n558), .A2(new_n671), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n527), .B(new_n529), .C1(new_n397), .C2(new_n538), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n319), .B1(new_n553), .B2(KEYINPUT81), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n545), .A2(new_n546), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n747), .A2(new_n749), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n618), .A2(new_n558), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n684), .B1(new_n758), .B2(new_n675), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n760), .A2(KEYINPUT29), .A3(new_n741), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n744), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n673), .A2(new_n510), .A3(new_n741), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT30), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n616), .A2(new_n537), .A3(new_n536), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n502), .A2(new_n497), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n634), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n606), .A2(new_n538), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n769), .A2(KEYINPUT30), .A3(new_n634), .A4(new_n766), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(G179), .B1(new_n623), .B2(new_n624), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n606), .B(new_n772), .C1(new_n499), .C2(new_n496), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n545), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT31), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n741), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT96), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n773), .B2(new_n545), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n616), .A2(new_n634), .A3(G179), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n780), .A2(new_n480), .A3(KEYINPUT96), .A4(new_n553), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n771), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT97), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n771), .A3(KEYINPUT97), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n741), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n763), .B(new_n777), .C1(new_n787), .C2(KEYINPUT31), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G330), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n762), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n740), .B1(new_n791), .B2(G1), .ZN(G364));
  NOR2_X1   g0592(.A1(new_n286), .A2(G20), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n247), .B1(new_n793), .B2(G45), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n734), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n223), .B1(G20), .B2(new_n296), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n224), .A2(new_n319), .A3(G179), .A4(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n316), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n224), .A2(new_n274), .A3(new_n397), .A4(G200), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n266), .B(new_n802), .C1(G58), .C2(new_n803), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n224), .A2(new_n397), .A3(new_n319), .A4(G179), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G179), .A2(G200), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(G20), .A3(new_n397), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G159), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n212), .A2(new_n806), .B1(new_n810), .B2(KEYINPUT32), .ZN(new_n811));
  NAND3_X1  g0611(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G190), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n224), .B1(new_n807), .B2(G190), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n814), .A2(new_n203), .B1(new_n815), .B2(new_n489), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n224), .A2(new_n274), .A3(G190), .A4(G200), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT98), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G77), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n812), .A2(new_n397), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n810), .A2(KEYINPUT32), .B1(G50), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n804), .A2(new_n817), .A3(new_n824), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(G311), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n809), .A2(G329), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n269), .B(new_n829), .C1(G322), .C2(new_n803), .ZN(new_n830));
  INV_X1    g0630(.A(G283), .ZN(new_n831));
  INV_X1    g0631(.A(G326), .ZN(new_n832));
  INV_X1    g0632(.A(new_n825), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n801), .A2(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT33), .B(G317), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n813), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n815), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n805), .A2(G303), .B1(new_n837), .B2(G294), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n828), .A2(new_n830), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n799), .B1(new_n827), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(G13), .A2(G33), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(G20), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n798), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n733), .A2(new_n266), .ZN(new_n845));
  INV_X1    g0645(.A(G116), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n845), .A2(G355), .B1(new_n846), .B2(new_n733), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n245), .A2(new_n383), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n733), .A2(new_n269), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n738), .B2(G45), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI211_X1 g0651(.A(new_n797), .B(new_n840), .C1(new_n844), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n728), .A2(new_n729), .ZN(new_n853));
  INV_X1    g0653(.A(new_n843), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n730), .A2(new_n796), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(G330), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(G396));
  NAND2_X1  g0658(.A1(new_n701), .A2(KEYINPUT99), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT99), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n332), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n325), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n330), .A2(new_n712), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n701), .A2(new_n712), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n742), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n862), .A2(new_n863), .A3(new_n712), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n693), .B2(new_n687), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n872), .A2(new_n789), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n796), .B1(new_n872), .B2(new_n789), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n868), .A2(new_n841), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n814), .A2(new_n281), .ZN(new_n877));
  INV_X1    g0677(.A(new_n803), .ZN(new_n878));
  INV_X1    g0678(.A(G143), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n878), .A2(new_n879), .B1(new_n880), .B2(new_n833), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n877), .B(new_n881), .C1(G159), .C2(new_n823), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(KEYINPUT34), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(KEYINPUT34), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n801), .A2(new_n203), .ZN(new_n885));
  INV_X1    g0685(.A(G132), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n269), .B1(new_n808), .B2(new_n886), .C1(new_n202), .C2(new_n815), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n885), .B(new_n887), .C1(G50), .C2(new_n805), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n883), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n823), .A2(G116), .ZN(new_n890));
  OAI22_X1  g0690(.A1(new_n806), .A2(new_n316), .B1(new_n831), .B2(new_n814), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(G303), .B2(new_n825), .ZN(new_n892));
  INV_X1    g0692(.A(G311), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n266), .B1(new_n808), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(G294), .B2(new_n803), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n801), .A2(new_n212), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(G97), .B2(new_n837), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n890), .A2(new_n892), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n799), .B1(new_n889), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n798), .A2(new_n841), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n797), .B(new_n899), .C1(new_n408), .C2(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n874), .A2(new_n875), .B1(new_n876), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(G384));
  INV_X1    g0703(.A(new_n517), .ZN(new_n904));
  OR2_X1    g0704(.A1(new_n904), .A2(KEYINPUT35), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(KEYINPUT35), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n905), .A2(G116), .A3(new_n225), .A4(new_n906), .ZN(new_n907));
  XOR2_X1   g0707(.A(new_n907), .B(KEYINPUT36), .Z(new_n908));
  NAND3_X1  g0708(.A1(new_n222), .A2(G77), .A3(new_n353), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n910), .A2(KEYINPUT100), .B1(new_n221), .B2(G68), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(KEYINPUT100), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n247), .A2(G13), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n782), .A2(new_n771), .A3(KEYINPUT97), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT97), .B1(new_n782), .B2(new_n771), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n776), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n763), .B(new_n917), .C1(new_n787), .C2(KEYINPUT31), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n866), .A2(new_n867), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n415), .A2(new_n741), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n699), .B2(new_n700), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n454), .A2(new_n460), .A3(new_n921), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT107), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n699), .A2(new_n700), .A3(new_n922), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n921), .B1(new_n454), .B2(new_n460), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT107), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n929), .A2(new_n918), .A3(new_n930), .A4(new_n919), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  INV_X1    g0732(.A(new_n710), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n367), .B1(new_n393), .B2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n401), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n364), .A2(new_n400), .A3(KEYINPUT104), .A4(new_n366), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT37), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT105), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT37), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n941), .A3(new_n401), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT105), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n938), .A2(new_n943), .A3(KEYINPUT37), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n367), .B(new_n933), .C1(new_n704), .C2(new_n695), .ZN(new_n946));
  AOI21_X1  g0746(.A(KEYINPUT38), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT16), .B1(new_n361), .B2(new_n362), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT102), .B1(new_n949), .B2(new_n301), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT102), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n358), .A2(new_n951), .A3(new_n277), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n363), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n366), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT103), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(new_n955), .A3(new_n933), .ZN(new_n956));
  INV_X1    g0756(.A(new_n366), .ZN(new_n957));
  INV_X1    g0757(.A(new_n363), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n358), .A2(new_n277), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(KEYINPUT102), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n957), .B1(new_n960), .B2(new_n952), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT103), .B1(new_n961), .B2(new_n710), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n956), .A2(new_n962), .B1(new_n396), .B2(new_n402), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n955), .B1(new_n954), .B2(new_n933), .ZN(new_n965));
  AOI211_X1 g0765(.A(KEYINPUT103), .B(new_n710), .C1(new_n953), .C2(new_n366), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n401), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n954), .B2(new_n393), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n941), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n942), .ZN(new_n971));
  OAI211_X1 g0771(.A(KEYINPUT38), .B(new_n964), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n932), .B1(new_n948), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n926), .A2(new_n931), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT38), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n962), .A2(new_n969), .A3(new_n956), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n971), .B1(new_n976), .B2(KEYINPUT37), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n975), .B1(new_n977), .B2(new_n963), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n972), .A2(new_n978), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n979), .A2(new_n929), .A3(new_n919), .A4(new_n918), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n932), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n918), .A2(new_n461), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(G330), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n982), .B2(new_n983), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n704), .A2(new_n710), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT101), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n862), .A2(new_n741), .ZN(new_n989));
  AND3_X1   g0789(.A1(new_n871), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n871), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n929), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n979), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n454), .A2(new_n741), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n972), .B(new_n978), .C1(new_n947), .C2(KEYINPUT106), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n977), .A2(new_n975), .A3(new_n963), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n996), .A2(new_n947), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT106), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(KEYINPUT39), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n995), .A2(KEYINPUT39), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n987), .B1(new_n992), .B2(new_n993), .C1(new_n994), .C2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n744), .A2(new_n461), .A3(new_n761), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n1002), .A2(new_n300), .A3(new_n705), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1001), .B(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n986), .A2(new_n1005), .B1(new_n247), .B2(new_n793), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n986), .A2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n914), .B1(new_n1006), .B2(new_n1007), .ZN(G367));
  NAND2_X1  g0808(.A1(new_n680), .A2(new_n603), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n712), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n685), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(new_n749), .B2(new_n1010), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n843), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n823), .A2(G50), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n806), .A2(new_n202), .B1(new_n879), .B2(new_n833), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G68), .B2(new_n837), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(KEYINPUT113), .B(G137), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1017), .A2(new_n808), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n266), .B(new_n1018), .C1(G150), .C2(new_n803), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n800), .A2(G77), .B1(G159), .B2(new_n813), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n823), .A2(G283), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n801), .A2(new_n489), .B1(new_n621), .B2(new_n814), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n833), .A2(new_n893), .B1(new_n815), .B2(new_n316), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT112), .B(G317), .Z(new_n1026));
  OAI21_X1  g0826(.A(new_n266), .B1(new_n1026), .B2(new_n808), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G303), .B2(new_n803), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n805), .A2(G116), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT46), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1022), .A2(new_n1025), .A3(new_n1028), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1021), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n798), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n849), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n844), .B1(new_n227), .B2(new_n304), .C1(new_n238), .C2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1013), .A2(new_n796), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n731), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT111), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n558), .A2(new_n741), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT109), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n530), .A2(new_n712), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n555), .A2(new_n558), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1039), .B1(new_n723), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n720), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT95), .B1(new_n715), .B2(new_n716), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n722), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n713), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(KEYINPUT111), .A3(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n1053));
  AND3_X1   g0853(.A1(new_n1045), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1053), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1039), .B(new_n1055), .C1(new_n723), .C2(new_n1044), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT45), .B1(new_n723), .B2(new_n1044), .ZN(new_n1057));
  AND4_X1   g0857(.A1(KEYINPUT45), .A2(new_n1048), .A3(new_n1044), .A4(new_n1049), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1038), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n722), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1061), .A2(new_n719), .A3(new_n720), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n1062), .A2(new_n730), .A3(new_n1048), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n730), .B1(new_n1062), .B2(new_n1048), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1066), .A2(new_n790), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1045), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT45), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n1044), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1072), .A3(new_n731), .A4(new_n1056), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1060), .A2(new_n1067), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n791), .ZN(new_n1075));
  XOR2_X1   g0875(.A(new_n734), .B(KEYINPUT41), .Z(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n795), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n558), .B1(new_n1051), .B2(new_n667), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n741), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1044), .A2(new_n721), .A3(new_n722), .ZN(new_n1081));
  OR2_X1    g0881(.A1(new_n1081), .A2(KEYINPUT42), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(KEYINPUT42), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT43), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1012), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1012), .A2(new_n1085), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT108), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1084), .A2(new_n1089), .A3(new_n1086), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n731), .A2(new_n1051), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1091), .A2(new_n1094), .A3(new_n1092), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1037), .B1(new_n1078), .B2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT114), .Z(G387));
  INV_X1    g0900(.A(new_n736), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1101), .A2(new_n845), .B1(new_n316), .B2(new_n733), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n235), .A2(new_n383), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n279), .A2(G50), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT50), .Z(new_n1105));
  OAI211_X1 g0905(.A(new_n736), .B(new_n383), .C1(new_n203), .C2(new_n408), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n849), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1102), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n797), .B1(new_n1108), .B2(new_n844), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n822), .A2(new_n203), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n805), .A2(G77), .B1(new_n837), .B2(new_n600), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n279), .B2(new_n814), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n269), .B1(new_n808), .B2(new_n281), .C1(new_n878), .C2(new_n221), .ZN(new_n1113));
  INV_X1    g0913(.A(G159), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n801), .A2(new_n489), .B1(new_n1114), .B2(new_n833), .ZN(new_n1115));
  NOR4_X1   g0915(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n266), .B1(new_n808), .B2(new_n832), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n878), .A2(new_n1026), .B1(new_n893), .B2(new_n814), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(G322), .B2(new_n825), .ZN(new_n1119));
  INV_X1    g0919(.A(G303), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n822), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT48), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n805), .A2(G294), .B1(new_n837), .B2(G283), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT49), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1117), .B(new_n1128), .C1(G116), .C2(new_n800), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1116), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1109), .B1(new_n721), .B2(new_n854), .C1(new_n1131), .C2(new_n799), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1067), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n734), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n791), .A2(new_n1065), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1132), .B1(new_n794), .B2(new_n1066), .C1(new_n1134), .C2(new_n1135), .ZN(G393));
  NAND3_X1  g0936(.A1(new_n1060), .A2(new_n795), .A3(new_n1073), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n844), .B1(new_n489), .B2(new_n227), .C1(new_n242), .C2(new_n1035), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n796), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n822), .A2(new_n279), .B1(new_n221), .B2(new_n814), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT115), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n266), .B(new_n896), .C1(G143), .C2(new_n809), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n878), .A2(new_n1114), .B1(new_n281), .B2(new_n833), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT51), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n805), .A2(G68), .B1(new_n837), .B2(G77), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1142), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n814), .A2(new_n1120), .B1(new_n815), .B2(new_n846), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G283), .B2(new_n805), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n269), .B(new_n802), .C1(G322), .C2(new_n809), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(new_n621), .C2(new_n822), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n803), .A2(G311), .B1(G317), .B2(new_n825), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT52), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1141), .A2(new_n1148), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1139), .B1(new_n1155), .B2(new_n798), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1044), .B2(new_n854), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1137), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1074), .A2(new_n734), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1060), .A2(new_n1073), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1133), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1158), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G390));
  NAND2_X1  g0963(.A1(new_n871), .A2(new_n989), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT101), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n871), .A2(new_n988), .A3(new_n989), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n925), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n994), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1000), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n760), .A2(new_n741), .A3(new_n864), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1170), .A2(new_n989), .B1(new_n927), .B2(new_n928), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n994), .B1(new_n996), .B2(new_n947), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1169), .A2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n929), .A2(new_n918), .A3(G330), .A4(new_n919), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n918), .A2(G330), .A3(new_n461), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT116), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n918), .A2(new_n461), .A3(KEYINPUT116), .A4(G330), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1002), .A2(new_n300), .A3(new_n705), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n788), .A2(G330), .A3(new_n919), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n925), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n1176), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1170), .A2(new_n989), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n918), .A2(G330), .A3(new_n919), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n1192), .B2(new_n925), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n929), .A2(G330), .A3(new_n788), .A4(new_n919), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1185), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1169), .A2(new_n1194), .A3(new_n1174), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1178), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1003), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1187), .A2(new_n1176), .B1(new_n1166), .B2(new_n1165), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1194), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n992), .A2(new_n994), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1173), .C1(new_n1204), .C2(new_n1000), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1176), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1202), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1198), .A2(new_n1207), .A3(new_n734), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1173), .B1(new_n1204), .B2(new_n1000), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1197), .B(new_n795), .C1(new_n1176), .C2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT120), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1000), .A2(new_n841), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n797), .B1(new_n279), .B2(new_n900), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT117), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n266), .B1(new_n621), .B2(new_n808), .C1(new_n806), .C2(new_n212), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n885), .B1(G107), .B2(new_n813), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n831), .B2(new_n833), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G97), .C2(new_n823), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n803), .A2(G116), .B1(new_n837), .B2(G77), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT119), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT54), .B(G143), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n822), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(G125), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n269), .B1(new_n808), .B2(new_n1223), .C1(new_n878), .C2(new_n886), .ZN(new_n1224));
  INV_X1    g1024(.A(G128), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n833), .A2(new_n1225), .B1(new_n815), .B2(new_n1114), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n801), .A2(new_n221), .B1(new_n814), .B2(new_n1017), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1222), .A2(new_n1224), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n805), .A2(G150), .ZN(new_n1229));
  XOR2_X1   g1029(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1230));
  XNOR2_X1  g1030(.A(new_n1229), .B(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1218), .A2(new_n1220), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1212), .B(new_n1214), .C1(new_n799), .C2(new_n1232), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1210), .A2(new_n1211), .A3(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1211), .B1(new_n1210), .B2(new_n1233), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1208), .B1(new_n1234), .B2(new_n1235), .ZN(G378));
  AOI21_X1  g1036(.A(new_n724), .B1(new_n980), .B2(new_n932), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n347), .A2(new_n292), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n291), .A2(new_n933), .ZN(new_n1239));
  XOR2_X1   g1039(.A(new_n1239), .B(KEYINPUT55), .Z(new_n1240));
  NAND2_X1  g1040(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(KEYINPUT123), .B(KEYINPUT56), .Z(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1238), .A2(new_n1240), .ZN(new_n1245));
  OR3_X1    g1045(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1242), .B2(new_n1245), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n974), .A2(new_n1237), .A3(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n974), .B2(new_n1237), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1001), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n931), .A2(new_n973), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n712), .B1(new_n915), .B2(new_n916), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n785), .A2(new_n786), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1253), .A2(new_n775), .B1(new_n1254), .B2(new_n776), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n868), .B1(new_n1255), .B2(new_n763), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n930), .B1(new_n1256), .B2(new_n929), .ZN(new_n1257));
  OAI211_X1 g1057(.A(G330), .B(new_n981), .C1(new_n1252), .C2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1248), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1000), .A2(new_n994), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n974), .A2(new_n1237), .A3(new_n1248), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1260), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1251), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1259), .A2(new_n841), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n269), .A2(new_n250), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n878), .A2(new_n316), .B1(new_n831), .B2(new_n808), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1271), .B1(G68), .B2(new_n837), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n801), .A2(new_n202), .B1(new_n489), .B2(new_n814), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G116), .B2(new_n825), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1272), .B(new_n1274), .C1(new_n304), .C2(new_n822), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1268), .B1(new_n806), .B2(new_n408), .ZN(new_n1276));
  XOR2_X1   g1076(.A(new_n1276), .B(KEYINPUT121), .Z(new_n1277));
  NOR2_X1   g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1270), .B1(new_n1278), .B2(KEYINPUT58), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n803), .A2(G128), .B1(G132), .B2(new_n813), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n806), .B2(new_n1221), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n837), .A2(G150), .B1(G125), .B2(new_n825), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(KEYINPUT122), .ZN(new_n1283));
  AOI211_X1 g1083(.A(new_n1281), .B(new_n1283), .C1(G137), .C2(new_n823), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT59), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n800), .A2(G159), .ZN(new_n1287));
  AOI211_X1 g1087(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1285), .A2(KEYINPUT59), .ZN(new_n1290));
  OAI221_X1 g1090(.A(new_n1279), .B1(KEYINPUT58), .B2(new_n1278), .C1(new_n1289), .C2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1291), .A2(new_n798), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n797), .B(new_n1292), .C1(new_n221), .C2(new_n900), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1266), .A2(new_n795), .B1(new_n1267), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1197), .B1(new_n1176), .B2(new_n1209), .ZN(new_n1295));
  AOI22_X1  g1095(.A1(new_n1188), .A2(new_n1189), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1199), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1266), .A3(KEYINPUT57), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n734), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT57), .B1(new_n1297), .B2(new_n1266), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1294), .B1(new_n1299), .B2(new_n1300), .ZN(G375));
  INV_X1    g1101(.A(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n925), .A2(new_n841), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n823), .A2(G107), .ZN(new_n1304));
  OAI22_X1  g1104(.A1(new_n806), .A2(new_n489), .B1(new_n621), .B2(new_n833), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1305), .B1(G116), .B2(new_n813), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n266), .B1(new_n808), .B2(new_n1120), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(G283), .B2(new_n803), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n837), .A2(new_n600), .B1(new_n800), .B2(G77), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1304), .A2(new_n1306), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n823), .A2(G150), .ZN(new_n1311));
  OAI22_X1  g1111(.A1(new_n806), .A2(new_n1114), .B1(new_n886), .B2(new_n833), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(G50), .B2(new_n837), .ZN(new_n1313));
  OAI221_X1 g1113(.A(new_n269), .B1(new_n808), .B2(new_n1225), .C1(new_n878), .C2(new_n1017), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1221), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n813), .A2(new_n1316), .B1(new_n800), .B2(G58), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1311), .A2(new_n1313), .A3(new_n1315), .A4(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n799), .B1(new_n1310), .B2(new_n1318), .ZN(new_n1319));
  AOI211_X1 g1119(.A(new_n797), .B(new_n1319), .C1(new_n203), .C2(new_n900), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1302), .A2(new_n795), .B1(new_n1303), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1296), .A2(new_n1185), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1322), .A2(new_n1202), .A3(new_n1077), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1321), .A2(new_n1323), .ZN(G381));
  INV_X1    g1124(.A(G387), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1249), .A2(new_n1250), .A3(new_n1001), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1263), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n795), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1267), .A2(new_n1293), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1297), .A2(new_n1266), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT57), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1332), .B1(new_n1251), .B2(new_n1265), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n735), .B1(new_n1334), .B2(new_n1297), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1330), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1210), .A2(new_n1233), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1208), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  OR2_X1    g1139(.A1(G393), .A2(G396), .ZN(new_n1340));
  NOR4_X1   g1140(.A1(new_n1340), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1325), .A2(new_n1336), .A3(new_n1339), .A4(new_n1341), .ZN(G407));
  NAND3_X1  g1142(.A1(new_n1336), .A2(new_n711), .A3(new_n1339), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(G407), .A2(G213), .A3(new_n1343), .ZN(G409));
  XOR2_X1   g1144(.A(G393), .B(G396), .Z(new_n1345));
  NAND3_X1  g1145(.A1(new_n1099), .A2(KEYINPUT125), .A3(new_n1162), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1076), .B1(new_n1074), .B2(new_n791), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1097), .B(new_n1096), .C1(new_n1347), .C2(new_n795), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(G390), .A2(new_n1348), .A3(new_n1037), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1346), .A2(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(KEYINPUT125), .B1(new_n1099), .B2(new_n1162), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1345), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(KEYINPUT126), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT126), .ZN(new_n1354));
  OAI211_X1 g1154(.A(new_n1354), .B(new_n1345), .C1(new_n1350), .C2(new_n1351), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(G387), .A2(new_n1162), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1349), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1357), .A2(new_n1345), .ZN(new_n1358));
  AOI22_X1  g1158(.A1(new_n1353), .A2(new_n1355), .B1(new_n1356), .B2(new_n1358), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1296), .A2(KEYINPUT60), .A3(new_n1185), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(KEYINPUT124), .ZN(new_n1361));
  INV_X1    g1161(.A(KEYINPUT124), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1296), .A2(new_n1362), .A3(KEYINPUT60), .A4(new_n1185), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1361), .A2(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(KEYINPUT60), .B1(new_n1296), .B2(new_n1185), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1365), .A2(new_n1196), .A3(new_n735), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1364), .A2(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1367), .A2(new_n1321), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1368), .A2(new_n902), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1367), .A2(G384), .A3(new_n1321), .ZN(new_n1370));
  INV_X1    g1170(.A(G213), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1371), .A2(G343), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1372), .A2(G2897), .ZN(new_n1373));
  NAND3_X1  g1173(.A1(new_n1369), .A2(new_n1370), .A3(new_n1373), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1373), .ZN(new_n1375));
  AND3_X1   g1175(.A1(new_n1367), .A2(G384), .A3(new_n1321), .ZN(new_n1376));
  AOI21_X1  g1176(.A(G384), .B1(new_n1367), .B2(new_n1321), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1375), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1297), .A2(new_n1266), .A3(new_n1077), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1338), .B1(new_n1294), .B2(new_n1379), .ZN(new_n1380));
  AOI21_X1  g1180(.A(new_n1380), .B1(new_n1336), .B2(G378), .ZN(new_n1381));
  OAI211_X1 g1181(.A(new_n1374), .B(new_n1378), .C1(new_n1381), .C2(new_n1372), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT61), .ZN(new_n1383));
  OAI211_X1 g1183(.A(G378), .B(new_n1294), .C1(new_n1299), .C2(new_n1300), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1294), .A2(new_n1379), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1385), .A2(new_n1339), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1384), .A2(new_n1386), .ZN(new_n1387));
  INV_X1    g1187(.A(KEYINPUT62), .ZN(new_n1388));
  INV_X1    g1188(.A(new_n1372), .ZN(new_n1389));
  NOR2_X1   g1189(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1390));
  NAND4_X1  g1190(.A1(new_n1387), .A2(new_n1388), .A3(new_n1389), .A4(new_n1390), .ZN(new_n1391));
  NAND3_X1  g1191(.A1(new_n1382), .A2(new_n1383), .A3(new_n1391), .ZN(new_n1392));
  XNOR2_X1  g1192(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1393));
  AOI21_X1  g1193(.A(new_n1372), .B1(new_n1384), .B2(new_n1386), .ZN(new_n1394));
  AOI21_X1  g1194(.A(new_n1393), .B1(new_n1394), .B2(new_n1390), .ZN(new_n1395));
  OAI21_X1  g1195(.A(new_n1359), .B1(new_n1392), .B2(new_n1395), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1356), .A2(new_n1358), .ZN(new_n1397));
  INV_X1    g1197(.A(new_n1355), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1099), .A2(new_n1162), .ZN(new_n1399));
  INV_X1    g1199(.A(KEYINPUT125), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1399), .A2(new_n1400), .ZN(new_n1401));
  NAND3_X1  g1201(.A1(new_n1401), .A2(new_n1346), .A3(new_n1349), .ZN(new_n1402));
  AOI21_X1  g1202(.A(new_n1354), .B1(new_n1402), .B2(new_n1345), .ZN(new_n1403));
  OAI21_X1  g1203(.A(new_n1397), .B1(new_n1398), .B2(new_n1403), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1387), .A2(new_n1389), .ZN(new_n1405));
  AND2_X1   g1205(.A1(new_n1378), .A2(new_n1374), .ZN(new_n1406));
  AOI21_X1  g1206(.A(KEYINPUT61), .B1(new_n1405), .B2(new_n1406), .ZN(new_n1407));
  NAND2_X1  g1207(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1408));
  NOR4_X1   g1208(.A1(new_n1381), .A2(KEYINPUT63), .A3(new_n1372), .A4(new_n1408), .ZN(new_n1409));
  INV_X1    g1209(.A(KEYINPUT63), .ZN(new_n1410));
  AOI21_X1  g1210(.A(new_n1410), .B1(new_n1394), .B2(new_n1390), .ZN(new_n1411));
  OAI211_X1 g1211(.A(new_n1404), .B(new_n1407), .C1(new_n1409), .C2(new_n1411), .ZN(new_n1412));
  NAND2_X1  g1212(.A1(new_n1396), .A2(new_n1412), .ZN(G405));
  NAND2_X1  g1213(.A1(G375), .A2(new_n1339), .ZN(new_n1414));
  NAND2_X1  g1214(.A1(new_n1414), .A2(new_n1384), .ZN(new_n1415));
  NAND2_X1  g1215(.A1(new_n1415), .A2(new_n1390), .ZN(new_n1416));
  NAND3_X1  g1216(.A1(new_n1414), .A2(new_n1384), .A3(new_n1408), .ZN(new_n1417));
  NAND2_X1  g1217(.A1(new_n1416), .A2(new_n1417), .ZN(new_n1418));
  XNOR2_X1  g1218(.A(new_n1418), .B(new_n1359), .ZN(G402));
endmodule


