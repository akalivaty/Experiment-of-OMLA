//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT76), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G113), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n193), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(new_n191), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT30), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G134), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G137), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(KEYINPUT67), .A3(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n199), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n203), .B2(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT11), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(G134), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(G137), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n212), .A2(new_n216), .A3(new_n200), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n218), .A2(KEYINPUT68), .A3(G131), .A4(new_n206), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n208), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n208), .A2(new_n217), .A3(new_n219), .A4(KEYINPUT70), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  AOI21_X1  g041(.A(G128), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(KEYINPUT1), .A3(G146), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n232));
  XNOR2_X1  g046(.A(G143), .B(G146), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n232), .B(new_n229), .C1(new_n233), .C2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n225), .A2(new_n227), .A3(new_n236), .A4(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n222), .A2(new_n223), .A3(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT65), .B1(new_n201), .B2(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n216), .B1(new_n240), .B2(new_n213), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n210), .A2(KEYINPUT11), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT66), .A3(new_n217), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n233), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n225), .A2(new_n227), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n249), .A2(new_n245), .A3(new_n246), .A4(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n255), .B(G131), .C1(new_n241), .C2(new_n242), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n244), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n198), .B1(new_n239), .B2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n208), .A2(new_n217), .A3(new_n219), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n238), .A2(new_n259), .ZN(new_n260));
  AND3_X1   g074(.A1(new_n260), .A2(new_n257), .A3(new_n198), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n197), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n197), .B(KEYINPUT71), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n239), .A2(new_n257), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT72), .B(KEYINPUT27), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(G237), .A2(G953), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G210), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n267), .B(KEYINPUT73), .ZN(new_n273));
  INV_X1    g087(.A(new_n271), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n266), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n269), .A2(new_n271), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n265), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g094(.A1(new_n264), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n262), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n262), .A2(new_n281), .A3(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n280), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT28), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n264), .A2(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(KEYINPUT75), .B(KEYINPUT28), .Z(new_n291));
  NAND2_X1  g105(.A1(new_n260), .A2(new_n257), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n197), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n293), .B2(new_n264), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n288), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n190), .B1(new_n286), .B2(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n262), .A2(new_n281), .A3(KEYINPUT31), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT31), .B1(new_n262), .B2(new_n281), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n190), .B(new_n295), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n189), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(KEYINPUT32), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT32), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n295), .B1(new_n297), .B2(new_n298), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT76), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n188), .B1(new_n306), .B2(new_n299), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n304), .B1(new_n307), .B2(KEYINPUT78), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT80), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n264), .A2(new_n289), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(KEYINPUT29), .A3(new_n280), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n239), .A2(new_n257), .ZN(new_n315));
  INV_X1    g129(.A(new_n263), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n264), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n314), .B1(new_n318), .B2(KEYINPUT28), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n239), .A2(new_n257), .A3(new_n263), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n263), .B1(new_n239), .B2(new_n257), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n314), .B(KEYINPUT28), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n310), .B(new_n313), .C1(new_n319), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G902), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT28), .B1(new_n320), .B2(new_n321), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n312), .B1(new_n328), .B2(new_n322), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(new_n310), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT81), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G902), .B1(new_n329), .B2(new_n310), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n313), .B1(new_n319), .B2(new_n323), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT80), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n262), .A2(new_n264), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(new_n280), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT29), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n288), .A2(new_n290), .A3(new_n294), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n331), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G472), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n309), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G119), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT83), .B1(new_n345), .B2(G128), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n346), .A2(KEYINPUT23), .B1(new_n345), .B2(G128), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(KEYINPUT23), .B2(new_n346), .ZN(new_n348));
  XNOR2_X1  g162(.A(G119), .B(G128), .ZN(new_n349));
  XOR2_X1   g163(.A(KEYINPUT24), .B(G110), .Z(new_n350));
  OAI22_X1  g164(.A1(new_n348), .A2(G110), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G125), .ZN(new_n353));
  INV_X1    g167(.A(G125), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G140), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT16), .ZN(new_n356));
  OR3_X1    g170(.A1(new_n354), .A2(KEYINPUT16), .A3(G140), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(G146), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n355), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G146), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n351), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n348), .A2(G110), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n357), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n224), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n358), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT82), .B1(new_n350), .B2(new_n349), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n350), .A2(KEYINPUT82), .A3(new_n349), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n363), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G137), .ZN(new_n371));
  INV_X1    g185(.A(G953), .ZN(new_n372));
  AND3_X1   g186(.A1(new_n372), .A2(G221), .A3(G234), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n371), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n374), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n362), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n375), .A2(new_n325), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT25), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G217), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(G234), .B2(new_n325), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(G902), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n375), .A2(new_n377), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n385), .A2(KEYINPUT84), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(KEYINPUT84), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n384), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n244), .A2(new_n256), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n237), .B(new_n229), .C1(G128), .C2(new_n233), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT85), .B(G101), .ZN(new_n394));
  INV_X1    g208(.A(G104), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n395), .B2(G107), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n397));
  INV_X1    g211(.A(G107), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(G104), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(G107), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n394), .A2(new_n396), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT86), .B1(new_n395), .B2(G107), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n400), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n395), .A2(KEYINPUT86), .A3(G107), .ZN(new_n404));
  OAI21_X1  g218(.A(G101), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n393), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n237), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n407), .B1(new_n231), .B2(new_n234), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(KEYINPUT10), .A3(new_n401), .ZN(new_n409));
  OAI22_X1  g223(.A1(new_n406), .A2(KEYINPUT10), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n396), .A2(new_n399), .A3(new_n400), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G101), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT4), .A3(new_n401), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n414), .A3(G101), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n254), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n392), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n409), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n238), .A2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n393), .A2(new_n401), .A3(new_n405), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n420), .A2(new_n391), .A3(new_n416), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(KEYINPUT88), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(new_n392), .C1(new_n410), .C2(new_n417), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G140), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n372), .A2(G227), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n405), .A2(new_n401), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n408), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n421), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n392), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n430), .ZN(new_n438));
  NOR2_X1   g252(.A1(KEYINPUT87), .A2(KEYINPUT12), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n392), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n437), .A2(new_n424), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n431), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n325), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n425), .A2(new_n427), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n438), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n437), .A2(new_n424), .A3(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n430), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(G469), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n443), .A2(new_n325), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G221), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n453), .B1(new_n455), .B2(new_n325), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G214), .B1(G237), .B2(G902), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT94), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n354), .B1(new_n252), .B2(new_n253), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n465), .B1(G125), .B2(new_n408), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n372), .A2(G224), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT91), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n464), .B1(new_n238), .B2(new_n354), .ZN(new_n470));
  INV_X1    g284(.A(new_n468), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n413), .A2(new_n197), .A3(new_n415), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n193), .A2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g290(.A(G116), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n477), .A2(KEYINPUT5), .A3(G119), .ZN(new_n478));
  INV_X1    g292(.A(G113), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI22_X1  g294(.A1(new_n476), .A2(new_n480), .B1(new_n192), .B2(new_n193), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n401), .A3(new_n405), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n474), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT6), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT6), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n475), .A2(new_n474), .A3(new_n482), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT89), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n475), .A2(new_n482), .A3(new_n490), .A4(new_n474), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n475), .A2(new_n482), .ZN(new_n492));
  INV_X1    g306(.A(new_n474), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n473), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(new_n491), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n500));
  OAI22_X1  g314(.A1(new_n470), .A2(new_n499), .B1(new_n500), .B2(new_n471), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n471), .A2(new_n500), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n466), .A2(new_n502), .A3(new_n498), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n482), .A2(KEYINPUT92), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n481), .A2(new_n505), .A3(new_n401), .A4(new_n405), .ZN(new_n506));
  INV_X1    g320(.A(new_n481), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n432), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n504), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n474), .B(KEYINPUT8), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n497), .A2(new_n501), .A3(new_n503), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n325), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n463), .B1(new_n496), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n494), .B2(KEYINPUT90), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n483), .A2(new_n484), .A3(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n495), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n469), .A2(new_n472), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(new_n325), .A3(new_n462), .A4(new_n512), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT101), .ZN(new_n523));
  INV_X1    g337(.A(G478), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(KEYINPUT15), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n477), .A2(G122), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n477), .A2(G122), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT98), .B(G107), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR3_X1    g345(.A1(new_n226), .A2(KEYINPUT100), .A3(G128), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT100), .B1(new_n226), .B2(G128), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n226), .A2(G128), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n203), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n530), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT13), .B1(new_n226), .B2(G128), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(KEYINPUT99), .ZN(new_n540));
  INV_X1    g354(.A(new_n535), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n532), .A2(new_n533), .B1(new_n541), .B2(KEYINPUT13), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n203), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n527), .A2(KEYINPUT14), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n529), .A3(G107), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n527), .B(new_n528), .C1(KEYINPUT14), .C2(new_n398), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n535), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G134), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n550), .B2(new_n536), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n454), .A2(new_n381), .A3(G953), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n544), .B2(new_n551), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n526), .B1(new_n557), .B2(new_n325), .ZN(new_n558));
  AOI211_X1 g372(.A(G902), .B(new_n525), .C1(new_n554), .C2(new_n556), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G475), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n359), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n353), .A2(new_n355), .A3(KEYINPUT96), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(G146), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n270), .A2(G214), .ZN(new_n566));
  NOR2_X1   g380(.A1(KEYINPUT95), .A2(G143), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OR2_X1    g382(.A1(KEYINPUT95), .A2(G143), .ZN(new_n569));
  NAND2_X1  g383(.A1(KEYINPUT95), .A2(G143), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n569), .A2(new_n570), .B1(new_n270), .B2(G214), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(KEYINPUT18), .A2(G131), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n565), .A2(new_n361), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT18), .B(G131), .C1(new_n568), .C2(new_n571), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n570), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n566), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n578), .B(new_n215), .C1(new_n566), .C2(new_n567), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n580));
  OAI21_X1  g394(.A(G131), .B1(new_n568), .B2(new_n571), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n365), .B(new_n358), .C1(new_n581), .C2(new_n580), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n576), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G113), .B(G122), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(new_n395), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n576), .B(new_n586), .C1(new_n582), .C2(new_n583), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n561), .B1(new_n590), .B2(new_n325), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n563), .A2(KEYINPUT19), .A3(new_n564), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n359), .A2(KEYINPUT19), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n224), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n358), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n579), .B2(new_n581), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n595), .A2(new_n597), .B1(new_n574), .B2(new_n575), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT97), .B1(new_n598), .B2(new_n586), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n595), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n576), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n587), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n603), .A3(new_n589), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT20), .ZN(new_n605));
  NOR2_X1   g419(.A1(G475), .A2(G902), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n605), .B1(new_n604), .B2(new_n606), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n560), .B(new_n592), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(G952), .ZN(new_n611));
  AOI211_X1 g425(.A(G953), .B(new_n611), .C1(G234), .C2(G237), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n325), .B(new_n372), .C1(G234), .C2(G237), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT21), .B(G898), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n523), .B1(new_n610), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n604), .A2(new_n606), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT20), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n591), .B1(new_n618), .B2(new_n607), .ZN(new_n619));
  INV_X1    g433(.A(new_n615), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(KEYINPUT101), .A3(new_n620), .A4(new_n560), .ZN(new_n621));
  AOI211_X1 g435(.A(new_n461), .B(new_n522), .C1(new_n616), .C2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n344), .A2(new_n390), .A3(new_n459), .A4(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(new_n394), .Z(G3));
  NAND2_X1  g438(.A1(new_n306), .A2(new_n299), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n325), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n307), .B1(new_n626), .B2(G472), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n458), .A2(new_n389), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n462), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n496), .B2(new_n513), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n461), .B1(new_n631), .B2(new_n521), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(KEYINPUT102), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n634), .B(new_n461), .C1(new_n631), .C2(new_n521), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT33), .B1(new_n553), .B2(KEYINPUT103), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n557), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n557), .A2(new_n637), .ZN(new_n639));
  OAI21_X1  g453(.A(G478), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI211_X1 g454(.A(G478), .B(G902), .C1(new_n554), .C2(new_n556), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n524), .A2(new_n325), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n619), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n636), .A2(new_n620), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n629), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  NAND2_X1  g463(.A1(new_n636), .A2(new_n620), .ZN(new_n650));
  INV_X1    g464(.A(new_n560), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n619), .A2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n629), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT35), .B(G107), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  OR3_X1    g469(.A1(new_n370), .A2(KEYINPUT36), .A3(new_n374), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n370), .B1(KEYINPUT36), .B2(new_n374), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n384), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n658), .A2(KEYINPUT104), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n383), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n661), .A2(new_n452), .A3(new_n457), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n622), .A2(new_n627), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT105), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n663), .B(new_n665), .ZN(G12));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n308), .A2(new_n303), .B1(new_n342), .B2(G472), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n613), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n612), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n652), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n636), .A2(new_n662), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n667), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n632), .A2(KEYINPUT102), .ZN(new_n677));
  INV_X1    g491(.A(new_n635), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n677), .A2(new_n662), .A3(new_n678), .A4(new_n674), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n301), .A2(new_n302), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n304), .B1(new_n625), .B2(new_n189), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n680), .A2(new_n304), .B1(new_n681), .B2(new_n302), .ZN(new_n682));
  INV_X1    g496(.A(G472), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n332), .A2(new_n335), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n684), .A2(KEYINPUT81), .B1(new_n340), .B2(new_n339), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n683), .B1(new_n685), .B2(new_n336), .ZN(new_n686));
  OAI211_X1 g500(.A(KEYINPUT106), .B(new_n679), .C1(new_n682), .C2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n676), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XNOR2_X1  g503(.A(new_n522), .B(KEYINPUT38), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n592), .B1(new_n608), .B2(new_n609), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n651), .ZN(new_n692));
  NOR4_X1   g506(.A1(new_n690), .A2(new_n461), .A3(new_n661), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n282), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n288), .B2(new_n318), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n695), .B2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n309), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n672), .B(KEYINPUT39), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n459), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n700));
  OR2_X1    g514(.A1(new_n699), .A2(KEYINPUT40), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n697), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  INV_X1    g517(.A(new_n644), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n691), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n673), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n636), .A2(new_n662), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n668), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT107), .B(G146), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G48));
  NAND2_X1  g524(.A1(new_n442), .A2(new_n325), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(G469), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n457), .A3(new_n444), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n390), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n646), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n344), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  INV_X1    g533(.A(new_n652), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n714), .A2(new_n390), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n650), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n344), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND3_X1  g538(.A1(new_n677), .A2(new_n678), .A3(new_n714), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n616), .A2(new_n621), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n661), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n344), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NOR2_X1   g544(.A1(new_n713), .A2(new_n692), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n677), .A3(new_n678), .A4(new_n620), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n311), .B1(new_n319), .B2(new_n323), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n288), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n188), .B1(new_n734), .B2(new_n286), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(G902), .B1(new_n306), .B2(new_n299), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n736), .B(new_n390), .C1(new_n683), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(G122), .Z(G24));
  AOI21_X1  g554(.A(new_n735), .B1(new_n626), .B2(G472), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n633), .A2(new_n635), .A3(new_n713), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n661), .A4(new_n706), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  NAND2_X1  g558(.A1(new_n446), .A2(new_n448), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT108), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n448), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(G469), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n444), .A3(new_n451), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n456), .A2(new_n461), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n522), .A2(new_n751), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n706), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n307), .B(KEYINPUT32), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n390), .B(new_n753), .C1(new_n686), .C2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT42), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT42), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n344), .A2(new_n757), .A3(new_n390), .A4(new_n753), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G131), .ZN(G33));
  AND2_X1   g574(.A1(new_n752), .A2(new_n750), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n344), .A2(new_n390), .A3(new_n674), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  NAND2_X1  g577(.A1(new_n522), .A2(new_n460), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n691), .B(KEYINPUT109), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(KEYINPUT43), .A3(new_n704), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT43), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n691), .B2(new_n644), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n661), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT110), .B1(new_n766), .B2(new_n768), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n770), .A2(new_n627), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n764), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n746), .A2(KEYINPUT45), .A3(new_n748), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT45), .B1(new_n446), .B2(new_n448), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n775), .A2(new_n443), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n450), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n444), .B1(new_n778), .B2(KEYINPUT46), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n457), .B(new_n698), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n774), .B(new_n782), .C1(new_n773), .C2(new_n772), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT111), .B(G137), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G39));
  OAI21_X1  g599(.A(new_n457), .B1(new_n779), .B2(new_n780), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT47), .B(new_n457), .C1(new_n779), .C2(new_n780), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n764), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n668), .A2(new_n389), .A3(new_n706), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT112), .B1(new_n790), .B2(new_n792), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n352), .ZN(G42));
  AND2_X1   g612(.A1(new_n712), .A2(new_n444), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT49), .Z(new_n800));
  INV_X1    g614(.A(new_n690), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n765), .A2(new_n390), .A3(new_n704), .A4(new_n751), .ZN(new_n802));
  OR4_X1    g616(.A1(new_n697), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n671), .B1(new_n766), .B2(new_n768), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n764), .A2(new_n713), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n754), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n389), .B1(new_n807), .B2(new_n343), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT48), .ZN(new_n810));
  INV_X1    g624(.A(new_n738), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n804), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n725), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT118), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n805), .A2(new_n390), .A3(new_n612), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n697), .A2(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n611), .B(G953), .C1(new_n816), .C2(new_n645), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n810), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n619), .A3(new_n644), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n736), .B(new_n661), .C1(new_n683), .C2(new_n737), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n806), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT117), .Z(new_n824));
  NOR2_X1   g638(.A1(new_n812), .A2(new_n764), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n799), .A2(new_n456), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n790), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n714), .A2(new_n461), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT114), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n690), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n828), .B1(new_n831), .B2(new_n812), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT50), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(KEYINPUT51), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n827), .A2(new_n833), .A3(new_n822), .A4(new_n819), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n835), .A2(KEYINPUT116), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT116), .B1(new_n835), .B2(new_n836), .ZN(new_n838));
  OAI221_X1 g652(.A(new_n818), .B1(new_n824), .B2(new_n834), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n743), .B1(new_n668), .B2(new_n707), .ZN(new_n841));
  INV_X1    g655(.A(new_n692), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n661), .A2(new_n456), .A3(new_n673), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n636), .A2(new_n842), .A3(new_n750), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n309), .B2(new_n696), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n846), .A2(new_n688), .A3(KEYINPUT52), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(new_n846), .B2(new_n688), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n344), .B1(new_n722), .B2(new_n728), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n301), .B1(new_n737), .B2(new_n683), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n459), .A2(new_n390), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n461), .B1(new_n514), .B2(new_n521), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n645), .A2(new_n620), .A3(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n851), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n739), .A2(new_n855), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n623), .A2(new_n850), .A3(new_n856), .A4(new_n717), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n853), .A2(new_n620), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n627), .A2(new_n628), .A3(new_n720), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n663), .A3(KEYINPUT113), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT113), .B1(new_n859), .B2(new_n663), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n661), .A2(new_n672), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n764), .A2(new_n864), .A3(new_n458), .A4(new_n610), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n344), .A2(new_n865), .B1(new_n821), .B2(new_n753), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n866), .A2(new_n762), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n857), .A2(new_n759), .A3(new_n863), .A4(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n840), .B1(new_n849), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n846), .A2(new_n688), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n846), .A2(new_n688), .A3(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n756), .A2(new_n866), .A3(new_n758), .A4(new_n762), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n623), .A2(new_n850), .A3(new_n856), .A4(new_n717), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n859), .A2(new_n663), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n860), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n875), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n874), .A2(KEYINPUT53), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n869), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n869), .A2(KEYINPUT54), .A3(new_n882), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n839), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n803), .B1(new_n887), .B2(new_n888), .ZN(G75));
  AOI21_X1  g703(.A(KEYINPUT120), .B1(new_n883), .B2(G902), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n891));
  AOI211_X1 g705(.A(new_n891), .B(new_n325), .C1(new_n869), .C2(new_n882), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n463), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n518), .B(new_n519), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n325), .B1(new_n869), .B2(new_n882), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G210), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n901), .A2(KEYINPUT119), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n901), .B2(KEYINPUT119), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n896), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n372), .A2(G952), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n899), .A2(new_n905), .A3(new_n907), .ZN(G51));
  NOR3_X1   g722(.A1(new_n849), .A2(new_n868), .A3(new_n840), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT53), .B1(new_n874), .B2(new_n881), .ZN(new_n910));
  OAI21_X1  g724(.A(G902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n891), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n900), .A2(KEYINPUT120), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n777), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT122), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n450), .B(KEYINPUT57), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n885), .A2(new_n886), .A3(new_n916), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n914), .A2(KEYINPUT122), .B1(new_n917), .B2(new_n442), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n906), .B1(new_n915), .B2(new_n918), .ZN(G54));
  AND2_X1   g733(.A1(KEYINPUT58), .A2(G475), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n604), .B1(new_n893), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n604), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n912), .A2(new_n913), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n907), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT123), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n912), .A2(new_n913), .A3(new_n920), .ZN(new_n926));
  INV_X1    g740(.A(new_n604), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n928), .A2(new_n929), .A3(new_n907), .A4(new_n923), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n930), .ZN(G60));
  XOR2_X1   g745(.A(new_n642), .B(KEYINPUT59), .Z(new_n932));
  NAND3_X1  g746(.A1(new_n885), .A2(new_n886), .A3(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n638), .A2(new_n639), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n907), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n934), .B2(new_n933), .ZN(G63));
  XNOR2_X1  g750(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n381), .A2(new_n325), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n883), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n386), .A2(new_n387), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n906), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n656), .A2(new_n657), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G66));
  INV_X1    g760(.A(G224), .ZN(new_n947));
  OAI21_X1  g761(.A(G953), .B1(new_n614), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n876), .A2(new_n880), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(G953), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n487), .B(new_n495), .C1(G898), .C2(new_n372), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  AOI21_X1  g766(.A(new_n372), .B1(G227), .B2(G900), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n795), .A2(new_n796), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n782), .A2(new_n636), .A3(new_n842), .A4(new_n808), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n759), .A2(new_n783), .A3(new_n762), .A4(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n841), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n688), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT125), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n955), .A2(new_n957), .A3(new_n372), .A4(new_n960), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n258), .A2(new_n261), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n593), .A2(new_n594), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(G900), .B2(G953), .ZN(new_n965));
  AOI21_X1  g779(.A(KEYINPUT126), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n791), .B1(new_n645), .B2(new_n720), .ZN(new_n967));
  OR4_X1    g781(.A1(new_n668), .A2(new_n389), .A3(new_n699), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n783), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n797), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n960), .A2(new_n702), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n974), .A2(new_n372), .ZN(new_n975));
  INV_X1    g789(.A(new_n964), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n954), .B(new_n966), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n961), .A2(new_n965), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n976), .B1(new_n974), .B2(new_n372), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n953), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n977), .A2(new_n982), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  NAND3_X1  g799(.A1(new_n955), .A2(new_n957), .A3(new_n960), .ZN(new_n986));
  INV_X1    g800(.A(new_n949), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n280), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n989), .A3(new_n337), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n985), .B1(new_n338), .B2(new_n694), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT127), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n906), .B1(new_n883), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n970), .A2(new_n949), .A3(new_n972), .A4(new_n973), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n989), .B(new_n337), .C1(new_n995), .C2(new_n985), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n994), .A2(new_n996), .ZN(G57));
endmodule


