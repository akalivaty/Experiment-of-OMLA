//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT16), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  OR3_X1    g005(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(G146), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(G146), .B1(new_n190), .B2(new_n192), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G237), .ZN(new_n197));
  INV_X1    g011(.A(G953), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G214), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT89), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n200), .B(new_n201), .C1(new_n202), .C2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G143), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n199), .B1(new_n205), .B2(KEYINPUT89), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT17), .A4(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n206), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n206), .A3(G131), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n196), .B(new_n207), .C1(new_n212), .C2(KEYINPUT17), .ZN(new_n213));
  XNOR2_X1  g027(.A(G113), .B(G122), .ZN(new_n214));
  INV_X1    g028(.A(G104), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT18), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n208), .B1(new_n217), .B2(new_n209), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n189), .B(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n218), .B(new_n220), .C1(new_n217), .C2(new_n211), .ZN(new_n221));
  AND3_X1   g035(.A1(new_n213), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  XOR2_X1   g036(.A(new_n189), .B(KEYINPUT19), .Z(new_n223));
  OR2_X1    g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n193), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n190), .A2(KEYINPUT71), .A3(G146), .A4(new_n192), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n224), .A2(new_n212), .A3(new_n226), .A4(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n216), .B1(new_n228), .B2(new_n221), .ZN(new_n229));
  OR2_X1    g043(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G475), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n230), .A2(KEYINPUT20), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n216), .B1(new_n213), .B2(new_n221), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n222), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G475), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n231), .B(new_n232), .C1(new_n222), .C2(new_n229), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT20), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n233), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G952), .ZN(new_n241));
  AOI211_X1 g055(.A(G953), .B(new_n241), .C1(G234), .C2(G237), .ZN(new_n242));
  XOR2_X1   g056(.A(KEYINPUT21), .B(G898), .Z(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT92), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n232), .B(new_n198), .C1(G234), .C2(G237), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n201), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n202), .A2(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n249), .B1(new_n252), .B2(G128), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(KEYINPUT13), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  OR3_X1    g071(.A1(new_n205), .A2(KEYINPUT13), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(G134), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n255), .B1(new_n259), .B2(KEYINPUT91), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT91), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n256), .A2(new_n261), .A3(G134), .A4(new_n258), .ZN(new_n262));
  XNOR2_X1  g076(.A(G116), .B(G122), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G107), .ZN(new_n265));
  INV_X1    g079(.A(G107), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n265), .A2(KEYINPUT90), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(KEYINPUT90), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n260), .A2(new_n262), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(G116), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT14), .A3(G122), .ZN(new_n273));
  OAI211_X1 g087(.A(G107), .B(new_n273), .C1(new_n264), .C2(KEYINPUT14), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n253), .A2(new_n254), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n274), .B(new_n267), .C1(new_n255), .C2(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(KEYINPUT9), .B(G234), .Z(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(G217), .A3(new_n198), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n271), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n271), .B2(new_n276), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n232), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G478), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(KEYINPUT15), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI221_X1 g099(.A(new_n232), .B1(KEYINPUT15), .B2(new_n283), .C1(new_n280), .C2(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n240), .A2(new_n248), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n272), .A2(G119), .ZN(new_n290));
  AND2_X1   g104(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n291));
  NOR2_X1   g105(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT83), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT83), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n290), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n295), .ZN(new_n299));
  INV_X1    g113(.A(new_n290), .ZN(new_n300));
  INV_X1    g114(.A(G119), .ZN(new_n301));
  NOR3_X1   g115(.A1(new_n301), .A2(KEYINPUT67), .A3(G116), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n303), .B1(new_n272), .B2(G119), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n299), .B(new_n300), .C1(new_n302), .C2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n298), .A2(KEYINPUT84), .A3(G113), .A4(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n294), .A2(G113), .A3(new_n297), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n300), .B1(new_n304), .B2(new_n302), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n309), .A2(new_n295), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n309), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT2), .B(G113), .Z(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n215), .A2(G107), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n215), .A2(G107), .ZN(new_n317));
  OAI21_X1  g131(.A(G101), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n215), .B2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n266), .A3(G104), .ZN(new_n321));
  INV_X1    g135(.A(G101), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .A4(new_n315), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n306), .A2(new_n311), .A3(new_n314), .A4(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n309), .B(new_n313), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n319), .A2(new_n321), .A3(new_n315), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G101), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g148(.A(G110), .B(G122), .Z(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT85), .ZN(new_n336));
  OR2_X1    g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n250), .A2(new_n251), .A3(new_n219), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n201), .A2(G146), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT66), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n250), .A2(new_n251), .A3(new_n341), .A4(new_n219), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n201), .A2(G146), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n345));
  OAI21_X1  g159(.A(G128), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n344), .B1(new_n252), .B2(G146), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n345), .A3(G128), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT64), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT0), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(new_n257), .ZN(new_n353));
  NAND3_X1  g167(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n353), .A2(new_n354), .B1(new_n352), .B2(new_n257), .ZN(new_n355));
  AOI211_X1 g169(.A(new_n257), .B(new_n344), .C1(new_n252), .C2(G146), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n343), .A2(new_n355), .B1(new_n356), .B2(KEYINPUT0), .ZN(new_n357));
  MUX2_X1   g171(.A(new_n350), .B(new_n357), .S(G125), .Z(new_n358));
  INV_X1    g172(.A(G224), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G953), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT7), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n336), .B(KEYINPUT8), .Z(new_n364));
  AOI21_X1  g178(.A(new_n308), .B1(new_n312), .B2(KEYINPUT5), .ZN(new_n365));
  INV_X1    g179(.A(new_n314), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n325), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n306), .A2(new_n314), .A3(new_n311), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n364), .B(new_n367), .C1(new_n368), .C2(new_n325), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n358), .A2(new_n362), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n337), .A2(new_n363), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n334), .A2(new_n336), .ZN(new_n372));
  NAND2_X1  g186(.A1(KEYINPUT86), .A2(KEYINPUT6), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n334), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n336), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n337), .A3(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(new_n358), .B(new_n360), .Z(new_n377));
  AND3_X1   g191(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT87), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT87), .B1(new_n376), .B2(new_n377), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n232), .B(new_n371), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G210), .B1(G237), .B2(G902), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT88), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n376), .A2(new_n377), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT87), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n232), .A3(new_n381), .A4(new_n371), .ZN(new_n390));
  AOI211_X1 g204(.A(new_n188), .B(new_n289), .C1(new_n384), .C2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n343), .A2(new_n355), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT11), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(new_n254), .B2(G137), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n254), .A2(G137), .ZN(new_n396));
  INV_X1    g210(.A(G137), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(KEYINPUT11), .A3(G134), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(G131), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(G131), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n356), .A2(KEYINPUT0), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n393), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT30), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n343), .A2(new_n346), .B1(new_n356), .B2(new_n345), .ZN(new_n406));
  INV_X1    g220(.A(new_n396), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n254), .A2(G137), .ZN(new_n408));
  OAI21_X1  g222(.A(G131), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n400), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n404), .B(new_n405), .C1(new_n406), .C2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n410), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n350), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n405), .B1(new_n414), .B2(new_n404), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n328), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT31), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n393), .A2(new_n402), .A3(new_n403), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n410), .B1(new_n347), .B2(new_n349), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(new_n328), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n197), .A2(new_n198), .A3(G210), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(G101), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n416), .A2(new_n417), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT30), .B1(new_n418), .B2(new_n419), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n327), .B1(new_n428), .B2(new_n411), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n414), .A2(new_n327), .A3(new_n404), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n424), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT31), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n328), .B1(new_n418), .B2(new_n419), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n430), .A3(KEYINPUT28), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT68), .B1(new_n418), .B2(new_n419), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT68), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n414), .A2(new_n436), .A3(new_n404), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n328), .A2(KEYINPUT28), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n434), .A2(new_n439), .A3(new_n425), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(new_n432), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(G472), .A2(G902), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n441), .A2(KEYINPUT69), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT69), .B1(new_n441), .B2(new_n442), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n392), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT70), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n434), .A2(new_n439), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n424), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n429), .A2(new_n420), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n448), .B(new_n449), .C1(new_n424), .C2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n451), .B(new_n232), .C1(new_n449), .C2(new_n448), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n441), .A2(new_n442), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n452), .A2(G472), .B1(KEYINPUT32), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT70), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n455), .B(new_n392), .C1(new_n443), .C2(new_n444), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n446), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT22), .B(G137), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n198), .A2(G221), .A3(G234), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n301), .A2(G128), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT23), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n301), .B2(G128), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n463), .B(new_n465), .C1(G119), .C2(new_n257), .ZN(new_n466));
  XNOR2_X1  g280(.A(G119), .B(G128), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT24), .B(G110), .Z(new_n468));
  OAI22_X1  g282(.A1(new_n466), .A2(G110), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n189), .A2(new_n219), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n469), .A2(new_n226), .A3(new_n470), .A4(new_n227), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(G110), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n467), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n473), .B(new_n474), .C1(new_n194), .C2(new_n195), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n471), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n471), .B2(new_n475), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n461), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n475), .A3(new_n460), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n232), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT25), .ZN(new_n481));
  INV_X1    g295(.A(G217), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(G234), .B2(new_n232), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n478), .A2(new_n484), .A3(new_n232), .A4(new_n479), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT73), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n483), .A2(G902), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT74), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n478), .A2(new_n479), .A3(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n491), .B(KEYINPUT75), .Z(new_n492));
  NAND4_X1  g306(.A1(new_n481), .A2(KEYINPUT73), .A3(new_n483), .A4(new_n485), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n488), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G140), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n198), .A2(G227), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n495), .B(new_n496), .Z(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n324), .B1(new_n347), .B2(new_n349), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n499), .A2(KEYINPUT10), .B1(new_n332), .B2(new_n357), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n257), .B1(new_n338), .B2(KEYINPUT1), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT77), .B1(new_n501), .B2(new_n348), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT77), .ZN(new_n503));
  INV_X1    g317(.A(new_n344), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n205), .B2(new_n219), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n345), .B1(new_n205), .B2(new_n219), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n503), .B(new_n505), .C1(new_n506), .C2(new_n257), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n507), .A3(new_n349), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n325), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT10), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n402), .B(KEYINPUT78), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n500), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n402), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n500), .B2(new_n511), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n498), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT81), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(KEYINPUT81), .B(new_n498), .C1(new_n513), .C2(new_n515), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n500), .A2(new_n511), .A3(new_n512), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n347), .A2(new_n324), .A3(new_n349), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT79), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT79), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n406), .A2(new_n523), .A3(new_n324), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n522), .A2(new_n524), .A3(new_n509), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT80), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT12), .B1(new_n402), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n525), .A2(new_n402), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n525), .B2(new_n402), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n520), .B(new_n497), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n518), .A2(new_n519), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G469), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n533), .A3(new_n232), .ZN(new_n534));
  INV_X1    g348(.A(new_n515), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n520), .A3(new_n497), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n402), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n527), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n525), .A2(new_n402), .A3(new_n528), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n513), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n536), .B(G469), .C1(new_n540), .C2(new_n497), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n533), .A2(new_n232), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n534), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G221), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n545), .B1(new_n277), .B2(new_n232), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT76), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n391), .A2(new_n457), .A3(new_n494), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(G101), .ZN(G3));
  INV_X1    g364(.A(new_n381), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n380), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n188), .B1(new_n552), .B2(new_n390), .ZN(new_n553));
  INV_X1    g367(.A(new_n281), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n271), .A2(new_n276), .A3(new_n279), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  NAND2_X1  g373(.A1(KEYINPUT93), .A2(KEYINPUT33), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n559), .B(new_n560), .C1(new_n280), .C2(new_n281), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(G478), .A3(new_n232), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n282), .A2(new_n283), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n233), .A2(new_n236), .A3(new_n239), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n553), .A2(new_n248), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n443), .A2(new_n444), .ZN(new_n571));
  INV_X1    g385(.A(G472), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n441), .B2(new_n232), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  AND4_X1   g388(.A1(new_n494), .A2(new_n574), .A3(new_n544), .A4(new_n547), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT34), .B(G104), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G6));
  NAND4_X1  g392(.A1(new_n287), .A2(new_n236), .A3(new_n233), .A4(new_n239), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n553), .A2(new_n248), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n575), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G107), .Z(new_n584));
  XNOR2_X1  g398(.A(new_n583), .B(new_n584), .ZN(G9));
  OR2_X1    g399(.A1(new_n476), .A2(new_n477), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n461), .A2(KEYINPUT36), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT94), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n586), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n490), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n488), .A2(new_n493), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n544), .A2(new_n547), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n391), .A2(new_n574), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(G110), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT95), .B(KEYINPUT37), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G12));
  INV_X1    g410(.A(new_n246), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n598));
  OR3_X1    g412(.A1(new_n597), .A2(new_n598), .A3(G900), .ZN(new_n599));
  INV_X1    g413(.A(new_n242), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n597), .B2(G900), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n240), .A2(KEYINPUT97), .A3(new_n287), .A4(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n604));
  INV_X1    g418(.A(new_n602), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n579), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n457), .A2(new_n592), .A3(new_n553), .A4(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G128), .ZN(G30));
  NOR2_X1   g425(.A1(new_n240), .A2(new_n288), .ZN(new_n612));
  INV_X1    g426(.A(new_n384), .ZN(new_n613));
  INV_X1    g427(.A(new_n390), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT38), .ZN(new_n616));
  NOR3_X1   g430(.A1(new_n616), .A2(new_n188), .A3(new_n591), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n602), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n548), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n450), .A2(new_n425), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n433), .A2(new_n430), .A3(new_n425), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n232), .ZN(new_n626));
  OAI21_X1  g440(.A(G472), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n446), .A2(new_n623), .A3(new_n456), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n612), .A2(new_n617), .A3(new_n622), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n252), .ZN(G45));
  NAND3_X1  g448(.A1(new_n565), .A2(new_n566), .A3(new_n602), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n457), .A2(new_n592), .A3(new_n553), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G146), .ZN(G48));
  INV_X1    g452(.A(new_n534), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n533), .B1(new_n532), .B2(new_n232), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n639), .A2(new_n640), .A3(new_n546), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n457), .A2(new_n494), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n570), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT41), .B(G113), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G15));
  NAND2_X1  g460(.A1(new_n643), .A2(new_n582), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G116), .ZN(G18));
  INV_X1    g462(.A(new_n289), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n457), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n553), .A2(new_n641), .A3(new_n591), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n301), .ZN(G21));
  NOR2_X1   g467(.A1(new_n453), .A2(new_n573), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n494), .A2(new_n248), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n553), .A2(new_n655), .A3(new_n612), .A4(new_n641), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G122), .ZN(G24));
  NAND2_X1  g471(.A1(new_n654), .A2(new_n591), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n635), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n553), .A3(new_n641), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G125), .ZN(G27));
  NAND2_X1  g475(.A1(new_n541), .A2(KEYINPUT102), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n520), .B1(new_n529), .B2(new_n530), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n498), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n664), .A2(new_n665), .A3(G469), .A4(new_n536), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n534), .A2(new_n662), .A3(new_n543), .A4(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n669), .A2(new_n670), .A3(new_n546), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n454), .B1(KEYINPUT32), .B2(new_n453), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n672), .A2(new_n494), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n384), .A2(new_n390), .A3(new_n187), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n635), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n671), .A2(new_n673), .A3(KEYINPUT42), .A4(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n674), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n457), .A3(new_n494), .ZN(new_n678));
  INV_X1    g492(.A(new_n670), .ZN(new_n679));
  INV_X1    g493(.A(new_n546), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n667), .A2(new_n668), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n678), .A2(new_n682), .A3(new_n635), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n676), .B1(new_n683), .B2(KEYINPUT42), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G131), .ZN(G33));
  AND2_X1   g499(.A1(new_n457), .A2(new_n494), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n671), .A3(new_n607), .A4(new_n677), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n678), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(KEYINPUT104), .A3(new_n607), .A4(new_n671), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G134), .ZN(G36));
  NAND2_X1  g507(.A1(new_n664), .A2(new_n536), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n695), .A2(KEYINPUT105), .A3(G469), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n543), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(KEYINPUT46), .A3(new_n543), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n534), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n680), .A3(new_n619), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n591), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n574), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT106), .ZN(new_n710));
  INV_X1    g524(.A(new_n565), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n566), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT43), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT107), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT44), .B1(new_n710), .B2(new_n713), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n674), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n707), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT108), .B(G137), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G39));
  INV_X1    g534(.A(new_n457), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n674), .A2(new_n494), .A3(new_n635), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n705), .A2(KEYINPUT47), .A3(new_n680), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT47), .B1(new_n705), .B2(new_n680), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n721), .B(new_n722), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G140), .ZN(G42));
  NAND3_X1  g541(.A1(new_n494), .A2(new_n187), .A3(new_n547), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n632), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n639), .A2(new_n640), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT49), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n729), .A2(new_n616), .A3(new_n712), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n600), .B1(new_n630), .B2(new_n631), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n677), .A2(new_n641), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n734), .A2(new_n494), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n568), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n713), .A2(new_n242), .A3(new_n494), .A4(new_n654), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n553), .A3(new_n641), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n739), .A3(G952), .A4(new_n198), .ZN(new_n740));
  INV_X1    g554(.A(new_n725), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n723), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n639), .A2(new_n547), .A3(new_n640), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n677), .B(new_n738), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n734), .A2(new_n242), .A3(new_n713), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n658), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n240), .A2(new_n733), .A3(new_n711), .A4(new_n735), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n748), .A2(KEYINPUT111), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n187), .B1(KEYINPUT111), .B2(new_n748), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n616), .A2(new_n738), .A3(new_n641), .A4(new_n750), .ZN(new_n751));
  AOI211_X1 g565(.A(new_n746), .B(new_n747), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n749), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n744), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n740), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n734), .A2(new_n673), .A3(new_n242), .A4(new_n713), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT112), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT48), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n744), .A2(new_n752), .A3(KEYINPUT51), .A4(new_n753), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n671), .A2(new_n659), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n566), .A2(new_n287), .A3(new_n605), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n457), .A2(new_n592), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n677), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n692), .A2(new_n684), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n637), .A2(new_n660), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n553), .A2(new_n602), .A3(new_n612), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n671), .A2(new_n770), .A3(new_n708), .A4(new_n628), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n608), .A2(new_n609), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n608), .A2(new_n609), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n769), .B(new_n771), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n610), .A2(KEYINPUT52), .A3(new_n769), .A4(new_n771), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI221_X4 g592(.A(new_n188), .B1(new_n567), .B2(new_n579), .C1(new_n384), .C2(new_n390), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n575), .A3(new_n248), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n549), .A3(new_n593), .ZN(new_n781));
  OAI22_X1  g595(.A1(new_n642), .A2(new_n581), .B1(new_n650), .B2(new_n651), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n656), .B1(new_n642), .B2(new_n569), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n768), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT54), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n782), .A2(new_n783), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n786), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n781), .B1(new_n790), .B2(new_n791), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n768), .A3(new_n778), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n785), .A2(new_n796), .A3(new_n786), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n796), .B1(new_n785), .B2(new_n786), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n789), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n788), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n756), .A2(KEYINPUT113), .A3(new_n759), .A4(new_n760), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n763), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n241), .A2(new_n198), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT114), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n732), .B1(new_n802), .B2(new_n804), .ZN(G75));
  OAI21_X1  g619(.A(new_n795), .B1(new_n797), .B2(new_n798), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(G902), .A3(new_n383), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n376), .B(new_n377), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n807), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n198), .A2(G952), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n776), .A2(new_n777), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n784), .A2(new_n692), .A3(new_n684), .A4(new_n767), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n786), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n785), .A2(new_n796), .A3(new_n786), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n232), .B1(new_n820), .B2(new_n795), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT56), .B1(new_n821), .B2(G210), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n814), .B1(new_n822), .B2(new_n811), .ZN(new_n823));
  INV_X1    g637(.A(new_n811), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n806), .A2(G210), .A3(G902), .ZN(new_n825));
  OAI211_X1 g639(.A(KEYINPUT116), .B(new_n824), .C1(new_n825), .C2(KEYINPUT56), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n812), .B(new_n813), .C1(new_n823), .C2(new_n826), .ZN(G51));
  XNOR2_X1  g641(.A(new_n542), .B(KEYINPUT57), .ZN(new_n828));
  INV_X1    g642(.A(new_n799), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n789), .B1(new_n820), .B2(new_n795), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n532), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n821), .A2(new_n698), .A3(new_n699), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n813), .B1(new_n832), .B2(new_n833), .ZN(G54));
  NAND3_X1  g648(.A1(new_n821), .A2(KEYINPUT58), .A3(G475), .ZN(new_n835));
  INV_X1    g649(.A(new_n230), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n836), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n837), .A2(new_n838), .A3(new_n813), .ZN(G60));
  INV_X1    g653(.A(new_n813), .ZN(new_n840));
  NAND2_X1  g654(.A1(G478), .A2(G902), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT59), .Z(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n788), .B2(new_n799), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n840), .B1(new_n843), .B2(new_n562), .ZN(new_n844));
  INV_X1    g658(.A(new_n562), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n806), .A2(KEYINPUT54), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n845), .B(new_n842), .C1(new_n846), .C2(new_n799), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT117), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n845), .B1(new_n800), .B2(new_n842), .ZN(new_n849));
  INV_X1    g663(.A(new_n842), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n562), .B(new_n850), .C1(new_n829), .C2(new_n830), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(new_n851), .A3(new_n852), .A4(new_n840), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n848), .A2(new_n853), .ZN(G63));
  NAND2_X1  g668(.A1(G217), .A2(G902), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT60), .Z(new_n856));
  XOR2_X1   g670(.A(new_n589), .B(KEYINPUT118), .Z(new_n857));
  NAND3_X1  g671(.A1(new_n806), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n806), .A2(new_n856), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n478), .A2(new_n479), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n840), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT61), .B1(new_n858), .B2(KEYINPUT119), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(G66));
  NOR2_X1   g677(.A1(new_n784), .A2(G953), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(G953), .B1(new_n245), .B2(new_n359), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n865), .A2(KEYINPUT120), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(KEYINPUT120), .B2(new_n865), .ZN(new_n868));
  INV_X1    g682(.A(G898), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n376), .B1(new_n869), .B2(G953), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n868), .B(new_n870), .ZN(G69));
  AOI21_X1  g685(.A(new_n198), .B1(G227), .B2(G900), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT125), .ZN(new_n873));
  XOR2_X1   g687(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n610), .A2(new_n769), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n874), .B1(new_n633), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n620), .B1(new_n567), .B2(new_n579), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n690), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n726), .A2(new_n876), .A3(new_n718), .A4(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n880));
  AOI211_X1 g694(.A(new_n875), .B(new_n633), .C1(new_n880), .C2(KEYINPUT62), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n198), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n428), .A2(new_n411), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT121), .Z(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n223), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(G900), .A2(G953), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n553), .A2(new_n612), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n707), .A2(new_n673), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT123), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n707), .A2(new_n891), .A3(new_n673), .A4(new_n888), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n875), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n692), .A2(new_n684), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT124), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n718), .A3(new_n726), .A4(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n887), .B1(new_n896), .B2(G953), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n873), .B(new_n886), .C1(new_n897), .C2(new_n885), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n872), .A2(KEYINPUT125), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(G72));
  NOR3_X1   g714(.A1(new_n429), .A2(new_n424), .A3(new_n420), .ZN(new_n901));
  NAND2_X1  g715(.A1(G472), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT63), .Z(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n787), .B(new_n905), .C1(new_n425), .C2(new_n450), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT127), .Z(new_n907));
  INV_X1    g721(.A(new_n784), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n879), .A2(new_n881), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n624), .B1(new_n909), .B2(new_n904), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT126), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n912), .B(new_n624), .C1(new_n909), .C2(new_n904), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n813), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n903), .B1(new_n896), .B2(new_n908), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n901), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n907), .A2(new_n914), .A3(new_n916), .ZN(G57));
endmodule


